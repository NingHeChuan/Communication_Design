`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R7Su66EFP3j7HdSRwT0ufavHZ21RJuR7GdMa5N1qrx05vZRLzNZT/TrlIe3c6DsFCenpiZCD2noZ
QAoR4Rt+mA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CMEJWch+GbdZ7DIDA14J94rfET0XyGxfytAfvkgCwK+buy8C6yPuTyczckBiUAmLYwq3N0YLZZjn
gsyXn6e48OgTdLuKlj0b1I+R+nOfWP/cHyUHpk91Upohu0q4i+T1Z7YlZ2KevK2O/yOn6S3pNXlM
CA1hIxQSQLLJQcJjXBI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IDWChuOHJQwebqfYcE88tSCCIBnxLv1aLHU6OnUVlxJuAYH1Wr0uPmJkkVb7CXm2iZXQx/jo6XaT
TumCKxTZIL3ET0tLNKmedouL0GaXfUzXVCSzEoTXiWf2gNPQB6+v0sryyUdggn9CbJglWE9UkluW
rCPI7feYIVKqODl/+/XlmC+0ONTNrMlZjktMivGmmfgFiOaVxlj7ZiVhYDRk2pmK7N0SbS8Yhqtp
tu4XIZyivSAfozOEYzRk3aC5YLPqYEODky8fadXC0TifmV1/9ihpE9MdNVbsAfiU6jAuYaPtixy1
eWfPyz8p770Y8aO4Ymmlv6Cov/zwD1Zr7rP3ng==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D4tWnXwgYbtbYBATOz3rKT5u236p/210UA0/0NawJUvRuLLRIOY863EXCqmoNKd3cdAJGfRGO/fA
mX3MQnn8fORd5NV0Drcjtq7LVURk4LrUaNUiho8FoaaKgENLoHWz5zN6jL9cfE19cPf5q6X+HSoS
vhMpVULwvEeloyESsidHnjc6Leo2s08QmBHWIJ4gX6Y353OK7qNS3bZaZnw5UMLbMBvsopLT0HMU
QgsF83OsAoA/LETx2kFpFT62GHW7Xr0WQupO68ddkWdncI1pQ1ry5DiS4IAcjHmDYTyo542wmUO5
kUoT65xdo6CgR0mBfndpvcIfOPFrzBLsA3X/8A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TYxxwxeYhuHcZvmvIoDp6PM6jwmqvK/EOpQJuzYEJwksrBgERfR0MxeEKttmbgtW3IAljWYtUY74
488K1yihiHHoprJ33R35ZxUze+TipXVo/GLAiCGp6aVvDPTACRhogMPXLJypmeRU1yO394pPbgS6
wC0P27Oimz3cJkJrwIhG7UV3FbbvFXVTh6Lp9wme459SE3zFnKsJYjUpffIirIVsuN+DETk1csWY
DA9UX9JySwER9tWjcgC7RtzEV1hjIG9WuwYm3zkOqr4FZ/dkK9PLm51AgWpaMXgB/7ws+/P8fkKm
QNdT6izgEuqxwJScjWNpExqD7cRIM9y2FibGuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y058Y7qqyKaMCwzJEnFzRJA1mSsdLWRJPV8jeagM24nQRyHL6Of41SQjwa7S6UfHPjaxh3kStD/R
iqFSj7BMeRnjDwKkql9QbQCQ1AEtG8kKMw6X1Sw8vQdkSSWaY8A0qHxlAj9yFFRWps0IUCT20y4r
a1FWV0KSxSpJrwls87U=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BkCcTwW7IOFCvnzvt27BUy3KHmy1QJwSQsGYOAQoWdJnp7bpQCB3MV/YrDTHZ6GeuEjTv+Y4jK1+
AUi7wPge8Y2zeEpQSTFjwsHrg0a6KicpWuoUxj9ZsRjp7lihT95V1Q0eAIg8YhlL39mGtTcQ5Vdp
7z8wKvjx++phq/T2pWg3qojhz3yoqaCG4uvKWuNn2R3f0YfPc7K1qQ8cRTBYuIfje99ZizVelHfv
/gPaALzJb7mtbJVe83NohlYy8IyL0cxXXClT+sW1XPYiN9k5NbywIoRmRDobstBVd3O4Ukd5mT3V
p/qjzuZHyCC/I/jJRQFyZvHI5rcbT8On+yp5MA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558368)
`protect data_block
inIHoKuztb9az5nMezpT+npf5U6KYQsfYW5Q5+6khYjIfg3alrIpTgmkKi/UvjzZogbrKLLT6ysx
56fYYqs9ckk2mE3P5H9LwfMFas1SEgH82G9Y6+5Br1Xbzh4Ng3/nORjYFCnh5bvNHjdnuwzzdW7z
xpqgLhGPbBblkNWOhsEfSA9+3JWF1F6pHy0xTb5GfqEHq6joix6PGPNgLTbbEzwQ5kB+cP4tDbIw
Y4ErMPeilEIdK9i3U5Ry5KBMx2xMOWIpGYjJpJgx/tgYXc+d3BaeVmLbF4dpGmN++MKR7XU0G1GO
uZyUNMdrpEFeIIt0gQzKvb0/nbioD1gnpCYLe129lcU1JLT4mwSUeclmpcXUj9ORP5BkRGv9Qxah
AKVepMghDBz5fgRHUUli7MJVt9p1aoadXkuQPudfmBf42GfpXKMi4lMjGwkKR4QHCTnl7tmntMKi
vEXewm6PKaDxFCtwNlerSY7IulTRduZhZ1bQ7xqf+8+HyAI3yYmp2dUqnlmiSB3SQ1bzfwwNsQvG
45TBj54x7ZOd5nOUBPLzAmF41n7Jehg7gpfeXdROONpH4us0xdSKCDarMx9E4CUnWbHj+2bQmW1N
h+G0u5u8jdX1FDeYseLW3+7P51D7FSmLDLwJCJPdambVs9fEvFe0UrNbloAK3G3W6xT6rveYIiDM
Vn2D8Cgs0smEcl2LR6rIEwONArRGPWoXEiby1NKvPGAWoDzpnt4skh7vtDtDkh6yO6yeBjIjEU1w
7DKF6aT87TIf552hKA8TDmjHeZGEv7CfnhQ2lF/pUx9J9AWcLu62VxdIYciD27ak3hhKB9j7ahHh
u0YVM2DC30Oqnic2rTxOCUle9Sv0rbM5Sn7psRYjCrhl/w413My89ndrfNZzO3WrzWv6njd4ydQk
SGWoVqhrn92SACa868cLACBVltd3e4y1ItK7tir4SLmFMy4S5hjMzgVFYo2imAF9p1AH/4SsScl4
m3fRsqjKlnqwKM4gwJdORlLUi6qYUMfIb4wZOZzh4BN31rSjwKBcyC9HXDYNoGZW3GGsYL2ME3wc
hGQfAAa3Q7EQOF4M5tNlzoKUE/fRCkqlncp14WKMTaPUCKKHBfPSCMAKMvWVCFguVPF2NU09O4xD
yhmt+RblkenHVOh2m24oRrUOL0Tw89QgZubkPIvnXp5s/K6FtavWVbF82l/4MH+vmfXQAyjgWw3C
LMII7iXsGgkVTrxBeiDpmE3GJHUJt02va7OmwqrxAaGblXSXnuOG0RP35gaXNYY3Lt4v7gcOnpP8
zVDlZksqpIePm/o6d9MPM99rRIiFu6X7OVWltC6ms1eVZw4TsJOqA1kBVIdH39sMa7J6sXkAgq9g
XQXwf3AeEt4+Gf5QW/ZGItHeCg07GZJTU81Xq065ZCOa8M4kXe11h3QUFBB9YbD1K8ea/F8hUpgN
kEC4ij9eV2R1pLNQcKNsbK6cay9nIv8KAbICZbkqi/Yhg4tG5LKWl0Mo3UmEmc4gR7VEyVlg2wgF
/JdyZrBOIMFy00fCW3LZVgsKOELrQI8gLSOqK/Aif6U0TD062YjlRjXL9EmbyhTTWTZmYxzDqpHe
dyPiEVybaKjvHhQEp4xOMb09c39PHK16a+L5NVVYpTux8Pvxs6uEQv1hzinfgj4LvMIO32S4lYyI
RZKYl15ZPReWlfyMTqaXio5I1UqliQhjjpNTsrhbV41W72rTagrSpRZ833twLXobwW1L1ifTzNdY
h8x73IK/OdShaQ1CPX8QI9S+ipB4cX/MGf2wNPLBqCPB3W7T3n4WPZJNfU4wXf1mTaUdE+MtxFi2
RLQ47prF8rx0rr+PUowBx9m40w4SYAsx9+lrrBwkvwONP/FLKSFVP8G3+EwktZHcobge+zVfkRnt
MX+MPzzhUg53HAdcdAF/+rc/4tcLZpc4OVmBO7Kt4DsmTMQWN3WVBKsaxdHARFH7Z+hJ2Wyr87EA
p9Y87VO3U6WMUa/JZhNda+qxVZd4TCRUm7qbmGz/BoDq3DyecZjRJ368AZxNCS4TqLxHKVwSoOaJ
dELJvZj2ph2FFYeXBeKJMzPabxfhCUUUUBHSyFLIa26LG3etITSXgimENnmi2lBzoy0062rw8s40
gl7NNncGr+Yj2O4IbSEJAI41juUyVo4G0s0BEhR/s8AQ+rpP4lPhH5drhkyJVGgd4+v1A+JFTcRt
847Tu30c1OTQtI3dAB1l6a7RSH1CMVNlhpmOHnDcvLlFm4YhopyuI2jM62cpoYNRD0iPqT5ELzFr
A6ZK6XIzcHF0zB+NGnfAz+0jxv/I+v5ybqo3GD+y3Ji5bB7+Q4UNdepSso6037NWOuY9RcmNGjwS
z0b2OOrLZIw1sSKwtVE/nviLaL4XujmzmnBUo0xy5bKYut6FNDIgBpee1Iamx7kO4+Qe0gffHdHT
8ZxL3gVfY+YUfm3G16InZ5ycGSgB3JifzIRoNa+6ubB0Zrf/y5GDt1oRWFTNLRmNR02mmRPkXjEF
Ru9g6ryPNnIy2ecuGPRiK6O6xgNWSer0m3i9YyC1btkhHG9C9w1tRj6CmwAudQY98KVL+FLd1khM
CGJdGNakZ++OU03F5nrJ4gK+Aqzk37Z3ZroGfCXjuxEz56y02wFFQl7AzJ50Ug5ZdBmtEuNIdpYH
53I2oFGQclPNQ27ya32BeKw/cZ7Zc5fLDgxtjqbD+k6VuzKDclJxVae+NZsc9ZM/Ydjf4F1aircP
2wa4piQiMqdfpWcqFGGDunN/O4C7FW7/vOj4Y2qIjteCuYdTMXUEuq2kVAVZUfL7qO+0GpR79zW1
P1QbO9KpNdaAbrYi3Hr8fyo7sffGhspaNqzpZ9MOU0AM8uJPecg7nk82EpqFSxW+PLFYfEbJm+zr
so+KXL/4VxxsVKUNR/tWNHJcos9DsJkspOLqKY4W00PIKu6Lxm0trMTXp5lLgJ8vgVervcyanmGK
xYPx2aVy4EzwgBnzR2OeQpIel/Bq0Cp3beQZAwQb3v/9YXZGnT8L2H+LX7aruRu2NSp4jCJmes1P
KZkGkmzWl7DunhjOecAEo5BNI5mdrY4FgY0pseikfv5fOWATgEUHgW3daLHZ7AU6AZeejzphSl7c
IPpnmn+nDhOVAWen2PBQNLH1xWRY5cP7hwuJXX5GE5o0Y3AFiY4hqg0NlEOq8IFoHGsS8IuNH3n+
JqUSkWcitVKbDx4vj0TEQ+beLxTYcHiCc2OnP57EavJ6+p7WQimAxOqza/Rct5eXs7mF+N4Y6J9V
Ra3X9sDO8wDgIwkkQnNR6HMlbgcumIK2UuM4aCd3mVQ5tDNA0T9XcPf3OBmwwMhvkQ1QWRQVw4Ma
lpjhNndw7DYFnNbwTu/WAN920Lpk8nzilb7cF4uaSloX6aMoKdZlPJ8vG4Ler59nmRQh4PcTdMce
uASNQJ7EBrGzC5oXTwU7jz0DhVAG15xeoH+aNcqaf9tyG3a4FxTXfW6YzkuT5wqg6oldiMe1cWQE
5ApxZWaBBcDoVHTJLL8f+ybvQqv/+XPnUZ/eCGvrwhrt1/60wqFYhEETqUPq1ov+ImDyFKd5QMve
a8yF3f4VfABvsLXgnx2R/Nqot0toaD3ZtJB28ywu7uYNrsnZPdm3AxD3JzoNrVfFoLyfjPXA6nnM
8fYi8f26PpVgpdFvhfxxWzJcVqorvB194a3FWoi6NntUkQbYioWL1wLEUKBrlsJy3KJiZjoNNejM
kXRcDUJE0LCatJXN2iBT0RbaAfQSFpUBfLnvZ8QGOsfmXFkLDPU6w8y569OAoJUm4/BoTsy6wW4r
e4eNA5EfPZ5uFCM9WyrxiJhz8PVw3jMo6WgUjx2y6IvWM37geF3YhE+WOTR8jXwySq1BwgKE/apy
+Pye+PkT/JOt6nMvMlc2KQ1HvVuEPr+q6BwVpBNFL7agL8NlSwImy/3LJ/r1xNXen/x2lWSCmbQ+
CYdRHrKoT3lfG1AsVM+IOg5mCEPRpuOOQ3ZHnvKulCcf3zEK6YAS4U0/+6SjXh/gP1Rx4LcOPa7a
Zp1+uL0uC68XgE3FUaFMbfKYuX5dk5jGzMPPfwPMMvwAQDdVjqXv4CABarzCugFJRLJv2ZCCQ2wm
iY74D2QBYfvZ4ZFwrcdlAUpqbIBl8imXdSNGHlR8cnSIK9B6ldphVIOIg/WoFJsoWTcBeTf+9zS3
sX9aW+XmM+vGvUqjV4DY8aNHUUXfLLt7V21z6JsCIGL6ad2w6e559D8fJfyHBr/FcOimPtm7rl2D
Ph9PMSIODi/kp9YsSudBRG4GRMuuPfPWcyJC/zp+DYNMgrw9bM3SE8aLBcqU3+XfSpXYioTHXsrc
vzwIa4jBkMM3PHAaxXHzbNtME9LRWtgyGbFH8i9U2KgETbZJnSz3I05o9xDyNcwAkPqQo+wMfZ2H
mU/LGi9LxlbQjp7VGQWcZOjzws6idhEw6hCqRnaElT9bcz5oAdS/P0inpwPJNTECnasSYJz+ywxm
EGN1h2XwbAORId9OTMAdYqa0ism/DerDiSN++wVZ0cGShcBgc0djdAPiD9YiexxXhfbUEiQzrf0w
ASpY8C6su04TCaLJ0p0Z2FM8ugOmBVMPN4u6WgHmHtrQ+NYNHpp0k8b6wiapbXhEvSuTmPa3ny1u
BO1BIL+YRDtjtNNOXqB1TkR8R5a6upFHg+bmO95q04hI4mMAlIQM7cmVNq1jBh1P9z8m8ak1RtZh
g6f6LLTUjTwrUiaRMVOUFo3JsjcyQM/Y6s77XTgUD+WQYS54h/Wv1GhTbS1IQE1yd1f38Bj8sjeB
lGlwmcwRZ5U1j0MaZ+UJIHFdiiM8anSUMuEITr3vdzcrZ/wJj+lmLdARs2hIuFUthPFPyAnxJIKO
DGLFaiuYtSWp3Sc8M4sz/u43r+G68Elu3i9PTyvOwhkzpTY8pik81x5tZvENmsaX2HLxrGbkIIgB
39py+K+5d51Y+yB4Yu6hlBz9PxS7QVB0GvgEr/+EBqV/BOgzUqJOgSgngRvMb49ptkrGDul9Dv4c
hQA/+37rtOsq0+lzH0kcMVreFoP3ErDw+2/snpl8kW26/YFKfeKm1Di1kX3xoSG56JkBvE1XeRM3
KVeTnXZMkzblaobRrA10w8LmpCgWo6lQa7Wh6Cyi5sGZfe5cX24BHkPu1SP9SgzX70utQJGamShF
auDhKvPBc8JaYH7IWcesIeWlJ15iKPVw2pG3HrRx4BvBbuPj7n++XbhD5qx2XAfkmrfXmJ4LmV46
KqrZgAZI2OPwgJsv4m70CrFZakNgIFAlLaTrrVKJ+QLMXJen2X3Hrfho0icQicAq3aJVpAOf8ObB
LizW4vgsO9/HwwSvkL0pCMsLGeIzY5YdnHBgLAdqLdvEln3qtKTqbqNJcALFsMP/aWcSM6+r39AY
rUGdOVBnpKBEIh77ovoPf4raPgqow96DX6DiRlj+mlNcPEz1W0OkH99AnHIMDU27chNhWzFJ8x7b
uib7yTsuhD2r8SaCR49c4QASFMmL2dHdOEqtuKJI6OKQXmOerMi2/YlQ2yF8RFkcXMsIAVIy2kAe
pWBEKqJNPo0qZZKFv99UPK2RHrofcND2rkAIRnTfLMyvm9ZqkHWT7k6WqL4UYhSnOWUcLmSJMIX1
NKG/nLK4ytj/7nTTI0OVWN0oxK/IuXTO1HF1A+wJ+odtsciZ13EgCp51hodtbyAgKZN1LUmOGUGu
zmvOVGWnqaquTwUCzQXj67u2sIDQjmtlX7/cTidj9fNLX7EkjNKI2f9FnXCtSm9xezbEZPkx01jH
VSuJ2bVM84rCsSwGCsMZMX3Ia9tBePuvyekpsXcGBtPS1m4V39kW65lOlNWMsy24+yjYQ0zLCnCg
a0mDFRsG8AaJRuwLGz5QRMHZf6Ue4u1ey1lOpTeohq5l4S8+ZHks6sKnELfW4FzeUWrMgW7lqDWL
gcV5zw5XiA4fwXGU2RQU9fNVgSNWwEFUNKRS7lwQdcM2svBlIO2SJ5x9qRT7sjdj+9dbcoYslTjm
swrRqSK2BT4jP8IH7hmIlpo9WrIpzRMhvMvzuGzxQ/BAjZwrCdcjpfvql5rfEY7qzAYB61wFNYTb
eZCMTNkbJqYg33Ld4T5WHn033E29dU7pncQbB5cxipvx7fqJFchTSh8jAelfntfRF38IRHSnc5lx
i1RuqKmRAe1jiNiahM9a7P3OsUwCKJf6PcztyiiQAPaCzFqSDRMxnTW787nFX4QVwd7gKIcfZL10
7lfi3QW/LdtctA/5Snv0ZnwIVSJ7mlLDJ0SutyxTvra/7E9emIyRlWnyA75dn91vPz+FDpCuUnAv
RimGnqanKe9d62LatHFkDih5EDkCqRtTQ50W6ox6Ts8quMEAraQK84IjzG41RIxqnroYxYD47R66
nzUa+wFYnrNtSVZfqc0pTKgsAqc9ktYo3TuwPi+H9jvN+NW2Tljtu8GN9RECXdhRaVxwMaduIH99
12qLZd/ALJpxY+9mPV6opwzQDsdWJFqN+Y6ml1a+DE9USwb4OxKlZnA6NmG3TpyGqFxMhL6Ppxlj
geq9NV7khYJuN30WsOSX36pixdiAd+2Ct9Gt4DTK7DgXh1sPglsrj5UqkGYZx4YaYGu7ppsN5uYK
Mds6iBAE6gpWOoV5gx2jxlf4Fbdg+jwlLVHB+J0PFu+i8s582AdlE5mTEFy13I2eZ/x9aJPa9pWW
EHCqGJjlDe+1gyN11rroBI+zu2EUZr0RTJI6h0uQBm9vbFzvLfpjS0GZ4vyfEbU5y/U9oSquEfuN
habgb4T0u6WpePlb4ktgBsrp0U+O0FQtxK0Udf4DcV790fJg4385cKBVCJxXQ9J6TsgmtCgK3uY5
xXHsYmRkXGSihufAb6gDwlKZ2GBRwVEW4RhptTV413FJnkHd2GfAzGYW1cWlpg0fjfBrxYEtv54a
+AA0ucDnrNBLH/FskrBGfiP5a1rLM25Scf0EGKp0J84gEzYuI7bXXRgVaW7dv5m6n8FAICQyBCFI
6hUNoSw9NVP5PonRj3I+4P/BTfL1gWtUo4hGdDAfYP1b1Li5IbUSlY4EEoiNlG5IWyLt05TrZ+lv
FXP0O+MN8kdw8S3G0Dz/Cao25rtp+k7OFxX5qOX0E7ZeKOOHc5/OrPqIAyS5YB8yBsBCZ7s15CKI
8Lo5m56rUFLh4LTOr9VTYZcNCrnQBv8aF7BPSXYVJPMzN8XYpX67vYpLep0RalO4Sw7Sfx86luWA
V0NacT1Yc8PD8pq5XWhwXVvWrWMXKHO5SeJfbAegWI9PmY34XluS0Xvx5U6RRv+OkFxpipUDnhBv
/+sCbrZQ1Sp3+Knbd1MQn6RdLUFaKElpd4VFHwchMnZi7D+9tTZensbMOME3BCSS+E532mTmWNd3
IvLWx7nGPDpcX+YYeE8d2H49gpaFlntDKpwewwXRilEhagI2IJ7INX4VsR8zUPj11wt3o2RS3kTV
fVlcjdQFFlY9x1kbQ383B4o10rEAe5JNDQUA55W8X5xlz2ZHtqSKCWT0f7ETbx5lTHu8wXqP2hd/
LbdV7QT8Xmh8TTbRqWqi+DKTWXK9hWXZm2b0ufDk7mWbmz9fVEjR56PsaMo/Cu0QI9Mx7XWfGk0Z
dAV5looSpOfswRX+ZTBSG7iyoMbJ18UngXiq9tX9yXv4INAEWQ4NlpImuFAz02eAYc2SNXonIHEw
VgAajg7FEpxU/zbLUmGozX6scEROh2v/m3cBglKLPw9QK6DlQNWRhGNJKpR6s8B4p0UJGb7VRNlm
r17T9OsbGCa2M00t2znnhP8BlHy8v1xbXa1dWiaDMDfspfatNXvYOr7wsa0n1M1sR8IEAMvqtmyi
C+7CyGc2y8lgAGNWqIpOKoT3Ny7bvnJU0IXE/i07MYZVnWxywnO7g+tMHgOix7QJRlevUnNuZWY6
VpdnjBBs2S4x7NsjaRXm8uBZ6iHQgH04JzsNWtWjjY55ohQ7gJtyaklYZ4ewak34FjStC+jAj3vO
I9+69YK7vHb4XBDtFckU9WNx38kyLkW/EDZ0g1e0n+D8pcO/DGwxDyMdzo87mJjumK/cWH5ks+lO
ANkDP8PyVfuV2ABMusvT3Bf3uTSfYBFZrp91x5sI6MOQp45nvUTJ6awmRnSevjVg4H5aCqTB4d3p
XDHU4SwOVk5yVbDbCCQQH5KV6BBzEsx5dcZsnT7weEnoBLnpssxq+lpClur+La7r70JYESuWZ9Fu
Zrbvui+NgyhdVp17LTE+svi5cCp90majzAwYjaT8FYWrYAvqNoGvTznzbxxKLDan0K4RKyyoDjTN
bNY//z1MTKpLBd8dt5w2sNQIjeThCNaJLd5ZBIXKjFcgfquJVMlsCW+alI/QELMu9FHZvGxOokDl
84Wu39TvYYivBBxlBHEVEwaotfuoUq83iw/vfLd70X3+4ZY84l/DA9NlnvC0+DuJmdt3Kxe7aC2/
Zm5sFzovAGzfxP8I5dKCtZn3RjGM+ZeyMQLTxrw3KVl4b7OSe6hLGhSfhAmSEd0CENxiOo6Xg2gM
qR+ivIQOxScFzCpavfGvUNOD6F+PBaNJxPlVwpnpRMFNhmYXNHBvA1nR+2AbnBwFQXE0Ta+BP9Hh
IPZ4s3Je9ahhVZwABv3olmSkLVTqq8vkLSjR+e9mYoT7MU6bAsNmLbIGvGBAyDKzEQAuwL6YS1aI
Pe0YSK+LSR1yh3ApgcEAstcRgzD26Th4IvDtkfz7wZSitg6i2DHdnW5IfXm8v4zvMCgBXISCsxQq
znh0xntu5E53VMLYFtflX2iWkDshqI3omwMUaTwg9yFNlbbdzL/1PufcIcLjSe4qRO38bwyzvHYU
vUv8t3cgoKYbSfguWdbqgkSPgovmWSsy803lkifnyIAcrIcJHLCWM/DZsVwCQw43ga8Gl8CfRDB2
BERp14by5U9i/rVG8/pzPAGGgvf+bpTJoxZ7Huj5MXw+9fWxYZ4NDAUe5Zn/sExLgh0oi/R2lrWT
HXIxbBEIBHtWgYLYfGXU7tw7avzQW+491i4fNSyBVK/wCxxWKK/AFLrsVXIX6zyJRVsfThsdrTbR
GGu+m0AfpK8s6g9WYnv7RLcKRkpl6nC7wcCfEKUv3KWfKpw08NDTblLkvr+xoWfLv6aB3J65d6fS
VnolJqG/jo88lZrOMK/EwRNuRXi0a8HcvJGacZp4RhMX0Z87fRomN6s/SnDGYbqsjWeWkpsCmMZb
jkwTrovNJkgoLonJ4THLhR72PeNhRwN1C3PJRiDqMy5v1fn1JUrD5q4fWNCi1vBeJsHrkToA2J0H
QtKtH0u1nsdghF8+8PiPs6YntloFS2btEm5zZM4yJjOLdkmx3iV7V0MXuvwVohw+95toV7pZhpmo
XkrXVs5hpivg1blKwMgeEoANfDZzURQy+QYYTv0CNtwORePnRpFe2uzJVmovY5kGgBVIntm7WaDF
uwEkVMLdT8o+j8rX0NI8KPWsRc0JeH2H7JihlnHr8MY13nZRRx7gZuutB529LJehzVW49N/DYUg1
Ji4IcR9VA43hq7YY/sGMECrE5qKJB+TxDiw/ZZierpqdxZtYAdgFDNmtcWRB+S+4Km3dU0xNeTXg
rvpC/TOnxeH5SqGCgjgJG2xxPokKLmcv9p1nwUTRFNXgvYAh9uHqLiyywk9AznIDKpBEKsUAZnz9
H0eDgTMLXQlrQ4c3pnxst/HUwdTNIL+D7MzTLRxW88FtYDzMoSLWwu34tWYlw4FihZNri+7b7VJ+
BYiIBB7MrJhzhfjdtdH/kEYfYWm30oy6lMd6UvOKY+p9QfdC2DCbYF5pcErlLxs1UX46Dk14dPiu
gAa4ohXzQia/hRyCiGyg+qV0Kc62neGwUo0plZRxld087unVq2ut9r5ZGYcgbHO0yklRWgorUnbE
irVgLmsuZ+OSXiTimfagFUdHXR5UrkrirNMzYDmhv77SNGWwDX8vrc96ERxqylIv9hKvsSIW8qrE
4aVkbSb868uwx1AB78zk6TkClStqN44yBn6iqyQvmVRhZDlewzVwarkcIPy2trtifYMihTwQuwRp
s8aLuZ+4Z89ck/GfPSEZRjvYwR5Hq/BZi9XnKFyOWSZii4rg4j2IshL6OxNJYDjT8en4le4HyJQ6
OlZzsblpjsTxZ5oujEeoN4KxqwftaJrAtmxP9s50TE7BIFjgptnloqajGkiximCVBKFXQYgHiLE/
HpubqDDFVORduugBE6aOUSrs0E3hL2/+aTGVvpmud9XH0KfUgNoTfuiAHHPd5R/kdB4slp49euXO
Q5e3jAMF51nB7PVskIXHXYoTPhwttKbusaWPWUDSgv8FAj+k1qPEht41REyz6MRrGZxfhjXuiknm
otW8Xd4XkKrsXFbYHetnewWyTaCq//XWZS+ITELd3d0vauWELTAr9CTcnfzr9NJXcRas2MgNJ1Ah
EQEcGwYZD0gpwDoi9/iqwj9mhM6yAo3ZhSgRcDRoWuQV0nDmMTOvK+W5PWSB6hvldDGhbfA1/Pkb
KKpoYzayi4G4naOWMYxRhPN+TBMI3OSEhvyUOTLKG0xJm6McIbSPdVrQZj+n9QK02+W+gtAVV0VS
Z/YL9GH4BrEtUT7FuCvaPdILzQIoDSR7kliAuxbfZAvNE+OXJbPrhLLAybgekXZP7jF43dcOwM8x
wmwf2CZ0SMPlulkpPc5JZVdZU2CJLBllyQNEIFPntLVFUqS3H2WXBzH8rEQAJZ/++FEBCWLpXaqy
2Klp5gn727barO8/GjZJzDe4Xr3a42yyohYi7h4bSsyW0Fd9wbQ64SSncu5g/+xtOvQzKYrjpZ4U
SsgtwYowklbhat+MsTrgLnvn4gQ+xC+jPrQlqpphpWSGY6paq965neZ49w8NF1EAvuBpaNVDx1Sr
YFjYeK2NFjI1gMoKACdj0jO6n+JaBOHvM99igBEiEQjNL3+JEy4QGN63m7ztH+IZ6GMzRE/9Zy3D
XVAgopc21NAkIdtF12zZuSED8QzIK1GDoTZvJ0e/94VlIaL+xiWGTVJhaM5ZPYL2OyVHx7nF8SBS
bBgZnFitarqZW8VVZs3bj1urnlxaWLetIUUSfs4E6pyIpHrq8fOBZW1z7PHE4UrnLV4fZLl8uoNW
aqRxurIsMXk2RKdrwg/LFAP9xj1Hl8Ts9RgXRxBfz19hrbVh6yFwYhFfPq2IsWRBABdDZLR36G0p
s2y6lfgJ7pg6yL8hwZbJJre1GQA4htcty+JoEoSScFt63am4WrUUP3dVYdYK5r7VI/BWUL4CUFiA
atRPXyRkxELleDLdUuIooOhYe4rcqtvr6/SUjmXJBr9SH5jEAjDIDSgtmlEcDuKL29qP4n2MX1/S
Aj478wq1lcogtUxekCjaBbMrIoa4fR7p4TdUSgFKqWpu/FBuAhXY32v9WmrK7r/zct9HhLmF5Z8d
1pzS5PiYkOoM5xojccV7PNYq9WfWu0NoR2EBo2OlSOc0hsmjJ1TyxwQ2mvCyjoq9nEjuIN28uTyn
QZ02nYyWWXyh07C9Ssa2ZLAnsyTRL8IO9iHV08FyPizPRqBQGBgpe2AukdBYcjxDZ05yg3c4yFTa
Ku8rQ6rR0Gy8wUMA3unv0KKEOCBxv9Xtgdo044Azx64hxUUic3abMIEO6oLcJBzFYUYZTqPHuc/f
b2sAMJzHqH+jFDOxfWq2TKWORbEciCIQdhm2p/VTvA13lrs3vxGffZ+GX+kIK+AjsAWR5A6nVwPb
beGJPsbRpliZZ25fQbxCVqlEskVlwsPGTrpWWzH7RT523ckzYQtxSghxDThqNOFqvfasYHu5B4lZ
djRuNk/RDKemJVzbGUW5/lQSunCaG0/18Rva24ucLGVQqzdPb2Pn/99BePS59EzhFVi8zdYs/qPF
9k/H7jW8HMMFbUZSeuQk4JXJ3JSQpWdXI2Q/KDkpKx2ggIfnLm5m9a6bhlKfFaujq6OufBFoCSI6
R55J/7X8BbmhZRFmdiUkJz+Y2NRr3NgnCF9W7tOP8GziKpl84YxwjpnBVI7Mp3ygDQoce+ENEST4
jK0Np3lRgYw0SmYJXYJK+6gXmXUveRpXE5chDccyuqqTdk0o8cgWxQ7t/NFP/0NQVd2i7EPDeRFF
F89PRbSD12r/BFS0Lp7Ar4CPlPm0EPx0flYwNSz77LXYoD9cyy03fgWBc0cTl+Qtw3euTo88/+2N
zsqIlnm53IO23FVyMdK/OlyOTiscOb/UtOC/g5rFBYY/loTS54fS+RrrA+MONmSeAJW98FL0m9FN
wD7szAqn98LGAjyV7RQdwplNiU45lMuGmVTBWKL/XP8477MhqixVWw8hWVRmK7cfx9ZyIOHuau+0
WKq8mG8nkBcxxea5J3lRS3TIHXVUR5Xs8IVPFyzlkpYj8wdnJphjRwqh/Gw0VsqpxZOahZ843hpf
s6ZFAFs7J+dZDyRy8v0XXjDrg8xclxYYnKcahmaP5kSFwMSunO1IAfAKalqmF0XxqSrYV+3PBJRT
Z6RYc0HvGn+qYorf8XSgLkb7aWOkEqcj1bK8Ajy/hOOMHF6ubowd68VGJ3v7vBT8JJYnFTRIbYot
13hw9yQgHvAJDwF7PjRtXOoj2MtBHwYW7ohR0SoryrpAT00yblzXF1BNPXkxGXZxZqcofnfglgeG
qSehLXpDZXD2EmK6r/jTnUjmHZxmdZRLY2JC07kKcvJ7tkrksB+KXEVz+vsPtcGQnU71T2Bcs4Ux
CzwydPz5L4ZvWgubwNiY/HTSvJC+WjCzZiglbDLeEJfHUaSOEQpWWVK4FTRZY3xkxUMFkcL6j/yl
H8kt+mGZf6nleqeEIYnNL4Vmb0sJQJ/Y1N5rfi38To1YQ2m6VTKoq3CYJaw0PlNF4V+VX9leyyY/
whjEJESEfECrYB58HvPv0Jn1/k8+Ze/hJ76BgSvK/YRRkM1xd731kDMydtQ6Bb4sXBmWsBFDG/D/
QLtcS2frmIZrbXywhAmXwdvBb/Wsbck3eSv+rhRWn3FM7uSwkVgY6rQhOUiLjQ2+DWd9XNKZasSm
2X0Fv6BvIXmyMuVWSkcH9HpnPXPvo+u7ut1DO8d7/mQzurzBrnz2ADjiGo0vQMyb1Rzy/54FD/+v
GChA5Cm1838Cql7mxsdsCskwAHcSbTV77ap57qXrG6Kz9q7Mxip0tg0uvj5KmBNUwxMNYWBaB3uV
eYicndkXjoYXdFA716KTC9Wm1M0jIq7DtH5wkzr3VcFFt/gyOogj6YeczqbySAaC6Dp+gHNIfmfe
cWonWDkYG8UcRyDG85dYZ42koLq3GUHpHT4MpB4FYUHRwNoZdW06CsYX1AzdbaiNql5mhJ3KcGzI
Ito/x3eerNz26GG+QEkhYP3s1Vp02eJZ6sPT+SS71/9pka0rIqrLNjhgToPP35Xx/lXuhoHDSgB4
uc1R9d868uXcT0bLzyVKdP3bitxX9tsSxRj/Ze9FzOVjT+nnKwbFolU8kK8tVOQP20fYuv09Gt6T
PRON8J5NzkLlZlkl+Y1w4Gpq2aXIxocOcIQN9aiV6sKvCW18FapzUSMBWLwLBZNZi7YYtdkUUiMi
a7Tk+p75EUDO/S8QZ594BTwNj/5WZkdLxpxyyuLNOzFu9+gdX4Lr+zcxB0Nx+/IOxKynoHuFSNd4
1t7L0dGhCUfZjpcXHoz4s+RHcw0wDG5HN56xdQ5/tr1praExDRWKPVw3w2njs6JxS19LHwoPzRmD
s2b1f7AbuBNTU73Du8a1/C8Nf+5asA7Gqiv4XRmnIc4KYmoI5pGBNmFHLaHUbl020IRWIpt5apR1
K9F/s3+EuOz9lErexMxTwONQ0nvcFdM2fHdItbE7MWisJbRe7apJv34JooyYEbXUB1mDMib2os9v
phOTlxoz6pEk3JXcl3uJkidqu1JPlS7gGOS3KpGMQrx/8EJPVkkDglNgitJ8YgePjvkAHyt3/rJE
oyVpcT0fVgLm/wZExgujO+SPt7SIbkgzAu175gOnA94DZv8NjuGH1AWU2+HzGwXdDF7NFXVsoB0T
mzd0hgW2UtVZtHBruZdObovmL3wOS1TiQvtu4ceCusQrJkNbOqxkOHUAOwkD72cyJzKL494iPMfl
wlPzNbSpLFRpLPbkcaxgaieL0HYGEuPLuEqbigB3ggOQTd2dtomGsmq5irOciB2E+XtW7OedIwVv
yB5eX1ZCx85tI7gITnrJUTMmNMWEoGziIyas4XjnyA7mM9QK5mowUE6L1k2D4oy8SpNDZoNdUTjo
6W9eNLrz/+nKAEMKRt2UEKZo9L6KucahldFeciG1E8j5f+0S8LPIAfnQCZaGzgYB0OSQUqr5hHN/
6XRqw+tvICz8iQucYM+JUUTOTPI8Z4POZRM5Pc4h2GhrVqcCXZhfZDke2wFUbcvBdD6aLsw/D2Jg
lGPUXokR0WCf9ClkIzagJNKnH7b7n/drAFSk2weWtRVkfttbu7qlwOGR3CYjYiXCpCBfZsuoRTya
+w66TH9VyPWPmiFe5xEVZkRGXwDKVp91kigqq7BKwLTyh+C3df8pc42VcUvZ/AiL9z7K15A+T4ke
T9VsEVlu+rhYYWTEUJ8e/fmaOA8Zi3kTBNl+cbKm+CVeuQdbf/0PJ6ETp0zxXo+SC9lgfXsflHnK
0dRP+jTAntAPylXK7ZWs2TmSuRYYGJY1Yiyii4oc6GTnAxRKNRNQY9DPuUUM1XQW6uMhfP3OA9xf
mvNHUk0lGC7F1XpaxFvjsvWpvWMJFx+BNTtk8Sc/mIUYwoQUMGxCgcq3Nu6TDynC3IU1RpU3vaMW
JSI5oRyxqM0V3Ffg8eoSkiPpIYYgRqCDnP3AZ0kDS6asKMey2d4Dql1tu4oW4x4OT7EwXW/RYkIZ
sUXAEZXELiri4H8Q78XeLZl/+f6yfWxn9Hgkn3pVxyWWE2TxPAWsP2XyS8RCqKvqWK/UAf3OrCvj
lu7D4NRdiSRaO6z82rbl6kw7BtteytZTU36TRbf0vVRYt396sdZ5FyMqCfEoy3jZGnPPhKwFAw1b
wo1upIaqaWqRm4EysHuvBvHdP163fUMBhoCm+JjVlDS7KZcT8J1SpxhECZ6nqpiZpjxnArR1Y7E+
KQkdlPJEVb0txALcT9/FUApysmmaZoSNyB8w/FaDWO7GrvGkOQCvMjpznpIGBOnofWi4Djp6S4rE
C7AsEdv303P6O96fj7QVwZilmhQ6LIAQxMDzohpn2f5REVc5riIXlkS4ZiER8JE4k4Uy7XVoMAb1
MVBSUGBb+i8ionu3xGW/lovjuKWMtY6QYeag29I4XkFtUyatS5kSyiL5NIKMZ1KUL6f5V+jvHOC3
hXVFvEikOa7XMXyzJ2MTyeSLRPqbCXwEz9mD5mODLLfXUGB+MjVJ4atUVeVzSGLpt84YSxlKloGe
wBZxYKBbwvyjVsTxpDCM1XQGuEAy66dfFcXCbMeAAz2fhomEVT4eotX0TnEvyBAntzAw8W/Q2XHH
5aGkSUzQGbZhcg+uUHRkDzT7zOla8kkCsXfG3UTVwjw0BwCrDkqjqUKCvB03iKfQUraVmk+tQfVX
7tN3PUWKL1WPxRqJaXGaft8kAo1wY4/CClvB9COIdjQlOSyqocBxsyxBNeRYpuXYkzKWMw1QuV5E
T8IlCWsNGrKMTg82rro2koxLjVZE6yNYm6hd1Uak8PBm9UAvdlvC0r5aoS45qdKWW7oqU0eD7Eun
fa8/sJRd5OxxW4dqbWHiLcB5nq87GHtv0T8xhmF5BZij99aUhyzh8AOK+nV1FeX9zwMj2nLmenr0
V9sCOZo0em+EH4woGJVv/zmLkKYPwfu5ZuJnU4YG2PbwGysTYAFD/4Xkgi4uqhLygx4BQX/424x0
sxy80kvbwAF0pJgYWD9s9Kvix01+13jygASRKtKTwAI89xU2pXirDN5QMyttT+yQHlc7dIL7H+5i
dwWtFw7ros+k2KV57SvCjowGxGPCwn+p0LwsrXGZYPZZHXASCXqpfiFYrSGNIWWixeBrvBQUEQ7G
FPeWdDIj3YP9T5WsiuduDF1rWIpkzQQKQqAysyI4fXSg02EPP8syP9mHaaAPHx6LbfcY65mhWT3U
p8tB7HTPI7REkjV/+/TCbozhn9vPU5wLn7l+I58DufPaQfZgIqyzidfsrMmvvuALmE2bwVoaHFl8
FSgNbQEqa7jRWc7UP3+kNeuzlS08+pcinAxSHEcDL3BdiraYeSTmcFaeR6U4JewAB2acJt0NF3G8
Oane9f1pDGQnSfItM0GzSezl95pvDG/zYCgJNZEuERLhrvvs0zUQbWjGj83NMz46Bkt+rSTxENL5
xR1WO8ySemKIZcg3G5L21DrqkJDfvVQbZFDwQlfFo4EgKlf1H58vgywO5L0owkhm557Y3KxPd1cg
VTcCVEV5mlk8lawgPyI62la98khjTp6uHIKHAUvQtp+8VWNfPFv1j1O4D4Bx14zui4f/h3J1IVvX
7gD7tg8whdWP45ARrHess5P9i22WkijuspQDxzAOJW6r1quc6WZiTxj+Sn8coUJ6Ae0GupoCayg3
Y4P2twy8AYfU0rt0zz/4B2/M7IwFKcwD1CZ4Cklq8sx5+JjBu5KpbLwzfyoOwWAvkd+iytbvEsV1
JQUORjfs5lDqg9CReqLj/FQWevphUEfTqbMnV68xrOS6vPHWm0MLlZX0NiF3abEW7ivDVpSbwVJV
1PVvZFNRqnOprp0bkK6zhgCMLIJYKgsPNLSFl+5VsztfojC7i4RcszUIH9UM/1LfRpSi3Rh67xin
FG+LcADVuCm2Dyptd/kbZNGOaVAohOI34FjjMOTsIUwcG2XFVw5ToWj28bcKSThsd0ZDXcb+vfy5
svz5oZkdiY8OZp+iEyX9/WuTvnFivhXzwOLdmXmHrgvZG9tGnPDOXcjxQoYeyu71d4WGMsRZ6B2V
K3WndGnUVbAso1W9T8cJQQYioLkh8px8Rqd8S6X57mT0r3Cn9ImhSgsdWzDMqvH/6IQeGlXnu7dW
RgAh3Fo6OPt3ShjbVVpfVfF+cTjWPI7u84YqB7Fn7J3b/PYiQr7taoWo97wN2EL8x0k70pCR+KBo
EdkZnoDSGVRuOoja2cn3RhJJ5gEGeycfoaXSj+lwuCcNqkNY8Q5uA/ecLjQgQDGN+hPKFl3Nqar/
UWuFttIS8RtcuUpxGJEKb74CN8dE/rnLCoJU//jyIbfeq/XNZM0n5CM+ZwXOnEL7v8gL5hbnGce8
NdUl/CNIY4DF8jU+GRMw0slcboor3hSG4tvWZy0T42RlJoahqKZT3kG1RBXcEhzQAR57hYc15t6f
Fyw4HXc2jgYfcsUxKop3gtWll7CnzpcGT3YZmuuEdABl8k+rcGWPLYOv41CI+zgJuQ2rPo/J3DY+
tj18bUaBpc7Sn6gDvTRrJZAC4F7Y+O4NjibGt4vhGgYJ0OwffE/iNI9JNpVKxfXRFp/jrWyPxjOI
Cqg2zIZ1xKEwux+vN3P9o3wY/NFvtBlHLLvcPG6s+RmZaS9un4tIpFxzTZ2oiUuaSoiGFiH2XMna
sTkI9bvY2SWxr4nsJT41GOmZFQ+kt3mwsrMOb/upIQR4+KptQhx3DjjQwZ3UvPLSY6k5SYe2QLCp
4TVguuDqWqxT0XbhhEhidauGaF7Gy72Q9mf9/TbFgJZtY+Jl+CLbiDI8ejsgnitzjGdvLFVPYHRz
Y+2XDb1PHUcsFf72S2GIvVqsJbT8DUICnEBwCoQy66Aeh927BtYc222iKNXDLDGyR9cPCoOAp9Ng
4HlEZyH4NqNbVrnF3AFTWp6Ys3t6tROH8VVaOqkawxfELe9studwE1hgTgitsOei+CHyi1l27bsX
7uqSqPOC5heloFkY2ajeaytF5f5nxwq89gSw+Pyn7aQ4we7KnsLbzt0peMa4+eFLfSOZzX4obHFQ
+5IdT7cRsT8VyswobhqXBoo2cbYPufU93fWlvmdg5Q6EPHzG4yhUkP/EunOt9MrymIk7ZVxVGp7B
ZUJHDUOkY/MMBHLukxG91BeE3gAqWtDRdeCFUqglgV8fPgYwK9ftsIAz+ea/f8XFlXLF9p7xeIs7
eFfunYb1PDomGZCBm8O27D2dwFs1wVtu3SJGiOe/G/yKSOpoRaNGDpOh0oAfJxVTJ7ZbQTbwscky
uIkf13DCu0PaIUZZykWlJ1kDN2vLu3WmO4PcMi/aKxKA4nOUzGslPLIHPiHYiMaAzSoOXfvTjnWC
RIVftouFJrV+3WyBCTmsfBhyJvDPhwrIVSHEcbVMF6MsfCsMKOsD7+XbjDivbe3TpCbT3exQOIAE
nuxkfUwcVH/fCc/J/5vjVry9tj9JAmuG/EZHqKuOUqHuaYiSAaIS+++GcasbeLJKpwWfa3WAbvGs
UpQqouiPhhOMDRCcIZofBTl5jWfjPk4yx54gE3dNMMhbObo78Xe9K7TxZurvz/wkf37DtqAMq0I2
iMma3l5qmxIJBfR8ASVk9/sNstMavVIORUOc2ERnCExu3tYtfL3xzkLuwdISHJkDN5pzHfyc8+wJ
G/rRKDvdIk577p/JGzrXNxwRhFAy222/K2jldXTEg+BQjgRDqOR7v84IymP2RhHEkKO5CFvt6wty
NE+G++oOOK1/39lT6OHDqO8rq2j4X/9vVdY5Hs2NtfBhniarotcrv8DepCvFc0Cns5E1wwRmavGP
Vw6furHAXyxbgUyO+J157sjggGI8zP4aY2oxYjfqTLE2VrrcWcp4Rt8oyu4i/Tp6mqoR7vfTQwIg
p9uRnxsW0J3didi+8hvXZ88o5g2DaQ57AvPQ9Uf3/an9rG4R8QPJGk+lfgFsy4PX4nk9G56usgq2
kNIwh+fH7eSvyNfQYMn/xhL/tZItGRt161K4ny7tHfJ0uzpYS1pKuDvcnjoMdoNVVOF7x6YCX2KE
MPJgQP6/yOWLAfCVtqIbNQ1im3ePzn7e6TAZ+lrYXybSVK2Wf1RLwCStcf5xxeZc2tz7DilcbaQX
WG8on2NxFh1Rhryxpc5ESHuYstjwITZ6qiOOG1jEQv0FKETczIBuWKVgujwBCy++XVtdayjoiose
RuE0QGnpj+HgDXKMHCNWgUMh7VLDXHCTXDY3VgvwgkNJlAduw6aOnOwJG3PFjFraQBwccHjJRUEp
YWq+UvpVCVbXxp9Tg4mD0eNsl6eHtZ1G4hWRCGR7gtThl0ilrytPZJiOOjVXypP+9Bvh2RXuNtjz
H1KBnaZf7nQrQ1RF5GcSdyg63b2jLMUP5KMpOgaM03CLeFQRynEQoOoNrgARSAJ0qRUPTSQSzKdW
tm9iZziHHL/nAEZrPyp5K8eqpiorlEsUF8hWU1Cmf0M6YBhMPU2+1DA1eMQL4opLSIEcq6izOTcC
VA4v14hyw7j3efp7cW/RXIb/x8yC36OWHdx5+E+h8MyPsyeA0Tj8LUPK02v6jkdRy8Qqlj7+7IxZ
ZfxAoBO6lA68i4esZB7DusBnfPtsVs9x9X2PLVEK4Sn7IaIUlY0v6hmPGnE5gO5TsLrj8EDwgTrf
Rqa2Nl3pXIScIpgExP4I5g862t/uncqY6xJTCEyEZv4efaOSUdmYPVSxxlWj7DKspSzpFPaeEDtl
1q37A/JEcSuMsJCC1vtY99TuVN+vanUdOWnKkfWf5gk2E03wGb+llJ2I7XSVJafKunARPRQaayVt
kaa7VzPsjN5BVHUGsoNQVBzwz9xPp0C7WyVG94YPZIJNhgcqXErvJgzHCPImQFKB1Azyf+mJ2Pww
GYhMLu6xxAn+8hTEUCia7SPqXw09ylug6qz/VN+nkThW3X5n3ANpJMX06pJSDZmu+/mTDJ/61Crn
9zXjIOWxUgwvyhfs9471sHcFMX0m9n345rZ/F/diJWItmT7UPRlbU2gjrpkP8ZyutshS3A7UHIZo
t4O31HTklYgxAKdPYawj79MepJWRmlTtgJSUcmJLXlMPMPJ2crQ7Cd6FfVzRP8DU65DrZrJIF6dw
GnHX41cX51WUNIEg/Lnc/6kT1KKDb8UxjuaEuGLAvVoWdXLyJubZ4a3aTm5SKjULo/lw13OeYAiH
dJ2Ni8x6Oj1sfwCD+GU+J4GwNn0Z4lEIow8btH359Zw2YjXkOjQFGU4DXwJkwrc4baLCwVq83xGa
57Cks9vu4PB61htU5f3iCoczVBmR5iMDG7iMUVajPA1XKoiruu/QpfjD8++55NHVb9PqL3ImZMUb
XgiyWk3p7tQpqV3XxwuM2VVlB8xi6/v4USZAWldH7jTxJMGzk6ai1iearMY7uRD5X6co0zOk6V8g
Q0Z5vsobw5E65Yq7SRvthaxM3y/wjjURwW5ROL4tALSmU1OMPb0ofMY5niPT69W7+x9Nagm1hEKo
H9dJp4zD+daclkseXldIpPzkj+HPgBA8goyTOwa63h/d8TjgNF05lavJaeHa2YkkBupQdXd1OciA
+tyo4iMa8xZ911nH4940xPiLwPOXoHj6Jsmj6iypJA0sfhryMRzOFiMDa6y39QcRBVQaOuk2FG9G
k0UCBYtMcccKPTZSLprhVr1PRyjO61SaSBDPj9jNFF/bzl4LflLltBzr0dGZ2cB8YD4sNymGn6qO
tzrOwjnZC2i2QssNwWFOh4pZIScImrpZlkSftGd27jVyHeI7e+v9cgtT+GcRh07LsDVC8IZERRpv
yfVfU9GkmsWyRliZzOy9/m9r566T1efxEPVWfti/smh9M2JIhoqITQ8dQkDbj56VcDJWCjR9AZY9
ppAdWqTSH4ZkgO0hM81w08aPpVpoVPfJbbNOwbKXz0eToYixRPJE56dCVIKebJIJeziCPbRXmEp8
yXISFoFC2w6ErAqH2AANn/ZtQq+/ND7W3u6vr+KxNjUIaN1cUyOoiPcjw3Co1PX02b5l7WDck+KJ
lLMlD6xS3DPxZk/kHN6nm8h16xOAikblRmr3iwO/rerWknyTk97aM4Cl4oZjj9J3sncDWr5OPRBT
brgsp54U9R7rI/WWGV439ErndXHmdtu2giRyFkZLnlSG7G74jKHQcaaY6AfDqiieqbMiIpn4kPow
RrTsEpFTokO6dawM3WnPDHB9kj4DkGhzDJyNocHp2MOe/N2S8I8syE93Gd4Q0j0xyhRy3g7N2Xc4
mzXh6xjFw9fNtRzlCcUOhj+WZUpasT23XlDWDfNjbJjzADW+YNN4HWFzn52FBHTUxex8FxJnU+SO
nf5rY7KHHn0dBDomrU2mWIavLr1kVHVWs7/f7dxOuvMITes6Tksxr4OgR96lkU2XddGf1GULUgbt
h9oHUcel1sKye3TCIn78adj9CQdfUJ/Y1EOFUgsjvFA3qCC7q/+m87Z2UHGZp83kn2upTcQ30gQJ
RqqTzWv2QBRJW+1v9AGZ1Kw0GDDCTg5VEcsMx4zzdABxW+ixRwcxuawzmZsovNCkBe4j92Mj/c+L
dmrsmSi0hqi9qILRI/dIUzYdhcORTiKmwE5KoDh36FUsyroiEytPmQMHn7ndoyjZk1Pf/lIKMAU0
aP8vdx2X0vJgl5jWd6Y8jZ22hNpkn+xU62iObnThfW/J4BJ4hhOzxva1pJvblwLLAjIOPEOYT5uj
dqrYs4tkhjsU6uW+w77CodgrAwDABg9i6+L59r1UG6voLNPbmOkodoUvIXkuXwPXoe51cANKZVZT
bhXLquzxsyJbSyOc8IhIerQy2mH6xS2u7OR2M6ZB0ejSQD5xOJVREZ7TLNdomOUOccqDRDwVeUWP
lxAulHquSEZhWBzdBtiZSOX2euTj1+vSsTsOoFlzB4BLrcGtRLR33C7SqBQwc8FqzddcUyyQjT/S
khvTR96cYKtBdZXhu4IXwk7083Im84HTMmO6jmC9rajSrAFnt7y64HJ1CMJ2eedKesSSReDYkadj
adt/wlWBXSlmmXmTEGA/2rIL7Xz1i5C07A2ejvXZydcZI+7ujGg0elrQT554D4zgQKz/qxKG0aNm
Iwd4N14w2jtMrZYBpFxMpWRv8iBhOm96st0Ryw9W+2hGZ9NukLe4G9mxuuKafF6teexVke3tfHGi
UxzzS/+8B/kfbTJ3IgwqxoM3Y+sWKHVAlhmwNBZ66NXzNUpWa+iwr/I/zHUvdaU/mhWIe2xlLVex
7PdkGkGhhrrN1XXRrsQrVWyiWDw19QpUwWNLzsQ5Zvkbck5wEGvhyVX0TsNyD9HRlPEV4d3X8BpH
pDxz6nhLpbZWnkViYEl7wiPUfKFS/peFHmJbj6v1tyd2xFidvA1ky7pG4oH3j63wh7nUCAtSLSO+
JJWvILZHp1/qWODZ2v8n+HT3sMW54tVb2X2XUDBlwXxp/yxitocG1d/8nEDDu1GlnmU2GzhkqRA9
1bXq9naRCA8E1H/8gNMcjBlQW7hUJUBI8uJpGaYYqbvYYAFOCQPEGP7irwJ3hha/fSFMhu3Lbgdw
hH0HlcBzoMNT812PJXF2p0Mqq5zqqRaZzgdatSlu3suG9J15hZmmwGgfOWdtQxKkKSOp8c63nDRI
eYSMAY7jhOgHYlGx3An1rxa9efF1oNIFQv7eZYYQPop0Ijb18gY6lNyfa+G3iDgnNsd0FYYkhbqr
Rkztp/mKBzpy2xbG53PW75A/dbahCqsONgPJbeym/8hCWMmVYrcYg6K0SXCZ8q5wQm4TRTbQ0rQi
HS9NwjUHxBkEGlJWw7BNdr7C97oufvUbPt25qI/wEiGHNzFqkjzjW6u17xGn1cdVDCe2Ixp9V3IR
7OICoQ9Pz5OecdjbQbtV1dFlY0h9TpOsh7HqU8vohoUH7SnQQxyUywlNNBjyBlC93DQ6F4hHuT9K
VjoLXfTrabj4AOEnEJiz3g5E+qoUuFuFtYi/rBaApT2p+CzU9aeOX8Kn+8C6xzSvgqZTxnM08JAH
bMekKbOgazujUW8YrnvvRSGXJDxE2DT7xjRQYljhyBCJ1aPNc722v4/ooyManWE61K5uJMP0f4Ww
R5Wz75BXJ/lQ9TcjddJD1BuScxWR6CRRiH3Yd/oeSkRpiO3I8kISMgsLhQYTQldERwupOYrEhz7C
wuG0cpSZ8R3piZZgN8K/7BqpTj5BUhqV7NNOZ9kM4gP4sN1FMyZKYmk5nLVeKYhbYgE+cXWafDvS
eDC99P6MPNB6Zdj9ZMulnZCKPz+2tzcdwRhxBCHpwG3NYs1nrahQHupelIgYJgTbCUEC8FgFXUWy
1bsYXxtXOQkvcq1dg+G2Uz+zzdabOqT1qCjzHXBzHbZ3OSmldguLbFiZe+INNaMRmto8CReXB1zJ
lyJfDwAPdhtyMvma/PV5Yt1hehA3Rfg73NMQMDtha7AVD4iUbIDB5KL0u4w0ztkl7ZRBgpE00c9V
qbt+DUviIhl+h0sKrmFBMX8ca/E3bkyTEQoq+nBKbX+pd8g9vIJutZdlOgvLER+LfBYLA2VaPtMd
QzVjYs81OWGhlKm7PHd/Q9RuO2Z7aX1e8pJx7s56UzvFw159sAi6lM/42OCHKCxiHdOlDRaZr6X9
k7bKRXHWW1/bK7B4vwRxPVPMZC0JRc3Tii0V1hwJRoODfOSH8a0nUKYOUTmyuzqxQqAL19xM+dnW
X6Nh9MNVZELgPFYwyx7xK3XMNlnRLk7G5LF6+Q2bWZSVCG+KGZwQaUF756JKUh4oNayBwT3FniJT
loGglPvl0fJwdC82Lb1NyzzxSgDECf1ePoRXg9TP7dmMNmm8fVGO6AkyNwGQQ/HPfpJHjSEeDMIB
84PaR0A+YXLQWP9UN6UD0NgmzQ6jDwpCV7PXXPLkaWUFyyl2sm/7xLG9Hsx113P2P3fmuoXXGesF
gjACWsp0l+99zck0Tgfdr/AMBT8g+k/5dXihC04wM76RT2OejNc1z/ltGCXi6mEqyr6W+NPVLxZ3
7i+9uB7EfG9BD0CYuZ17jysdR08HTmErVPVY0Jp9BuHw7znXee32uoxfn4zhbmCzfUn5oqwVJlBh
BYJPHf6zu+jzw1ZIPd5fMpH4jwDGN3KNOE8MT7529e+7k0jWJy4VbgvaYKF4Gt4lIOHSHBCuHr2P
T2Jky0cD3F0AG/goag9ZKJz7vM1iFTVX2AoZFlc6guMBrmUCkWlr6UwzaAe4iJJMORl7Nzo4o7rK
q/pVWSC4ad8B1HZgoALOGVoH/Ko/PRRt2FnoH1x1J+yjyM2oVctEixFdIAGns+m2VG27pPuWF9Cr
qe8/M6c6UHDwac85E7tFWV9v8OAcw0/8bVvqCOqgo7S5+34NxikuhEK/0i8F9r6Cj/dICC3aTzbE
SvuYWN4+0cHJMqgY+huY9pn8DuD52BdESl170X17bmdGv+yaPAYGAXxN52RbxqLoFLRZerMm0JiA
O8oVAyi1JTzJDp1Xes8Z3jC6m7aDnjCNQhhg/z5QtIvCqWjPzxULG9dRwh3r5TpTphD6pZrgvJCJ
dY2KK0hjDFFRALPBDndZO7kjrnS3XcqB3VHz0tFMIIJv2r9dc9LMqJYMxZdzGe1uUOsbyI4Tsjle
JPko14Flk9+cTfp9haBRuEI6LrecjLaWC1wTfEChE7o6tUrG2MhYZGQ7ceuOhxHETFpQAiSmnBv8
c3hGXoHo5yHTeByTf2e0Hk9QInxs1piIfFWi0D3S+cSlWx7/XS6fqWex6KG+UfEBYLxqq/tqyp+A
Rxji66//yYSNqV5uETlB9snzQyUgYalG5fe02EU6zeAOSXLb5T7uh5bazSV+b0KJI1eNNJQFwhfZ
vlkoLJJ9kyUe3C1htqO2axPIjxsRc/hEqCUGnc8VfTKzkitoh0u+fzIGgLhg7MUjPKEZ/pNsxk9d
ns58eDCTAx8GOoWSPG17BpRiU9NMlzxvilDDg/RoqKZPebQ7VdJ4PekfMhJ8+iseQydH/Zj9Tnkk
uco1Mfdm/HhB1xaiZOimovN80c3Kg7k9B4mnpVdkfnvaspfxckT+b9r2Yn8GsrSU+L3TBhIHgLz+
6rqpc2bye9sqmKbcqsnYeIauAJOBouVifU6SxWVjsDV6mER1AwRV264eVvRzTAFSMdhPp7gtTcOE
X9VJLfmasdwCIABZ02hK8e9D46JBPtSk5q9qDEktKMtjEE5ASpL2qYpFZweN8s66D5REOj8E/595
uraDcujo6FtJibbO6Y8wKurPKVpXRvUr8mUdmt39wikMtrmJovNHEz1mHiAaP7nWDxX0fl3QJHG3
1U4Qooj0WC0MllyiT9GCuktviIDUNz05huz72DbZQcok329ciAIvX/xvkzPUhXasRrZ4QW15da8q
9Nzux01T/KPJIM461vPsZC/Z6d9tdcagH3jYHGh6IRKx9Bi1nNtWEx2dmvAFXIPDdWSU2KDnC49o
RqD8Twf2zm7y/MuBtn4o79XakaFrmWlgjEcyA/cBQbzYxGjWB2Cf1MbivTHup3Q0Pb2Y562Iiywz
aG100a6Hn2u+xVTLO92uOiLTxtc2NuTjUcxT/PDtRNHZ+Hh0xomtkyavJSCUwZSw+MoDVbpCSFu9
2UrLV6WfOyFHKAtUh4m0LCy3CHnS43rV1Ayi5+/HFROOZRMHmCDfgOwnoPtksiPwQvzY538PDKj0
NiFUS1+nei/d9d8fnu4Vqbjq8AaM981lOo7tTJHgGaWd+PiGqK1HpZRDi3T6Py0C+eJR0RQpByUC
Lk5N52IYvRYpcXPxxvFTON+8zM5oLKTJmqDiIJe03zp+FPIP5XbnTaAPAFX4Fnk7lNM5X1ZxdSmH
jopcFsc3vJlagO99OtANsaq034IBuz5WDS6QWJFapEc2jhyRDrSLEHB4TCl37/XFwv/m+sIV9EIQ
m0MIHeWi59hS7U8lz1RsFXMUsBrWH2G15MBU3Ta/w0naXauX7lRtGwIf3kwGQeUS1PxTltK+nl8N
DJe1ndtXxRdve7IGI46FjsMdRcz/3GlJ2nZkeuQyv/2VhW4Nt3/F+ySWqLwbQ7fGJhM9oKG7Mxey
aIYN+9+hY98D0WRJGCroT13drfvAeXBw/o0ENln1yzNaP3tHmfj23Zkx9a4CJEJxxhRcFGU1y/5D
lp5gLKKU/tjxjbMztAkzG5ONlATs9MHMH8e4t5X3WQQ2Szh7kjkWav2QO/gpGlnly7AbBKauekBk
Ai661fnYFaCcGcsbKTdePkR9PglFDnRBRF8HOCYS5t45RkIIJFr418gVZbyiwce3e9elalKsQhis
Qz5n/mT9RnQ8idGM7rhaN5CJPScTX7hMg8iomD/Fq4i0QRH7svzUWfdeF150B8m42DVBuWpyV5dd
rcAiOynTIxjwgeiDFPXcbGEQLq0kwbhPjr96TbjBMjOKWaUgtfN5NBitHaB8Hnv6l04mvl13msNo
Jdx42/h0AdzOUCSs6zEsUrHGNyJu5KlcXWnQyI8bz7R+Qu8TazMSWx22dUAONxdkyWiLLUR9H3Ih
LYSVx0JhVGqVZoL3xx2COC0TWs6w+yqFc6akR6qppkpNA/SWFkpztBHcyygY8Kk/vtQCsu8eiPah
v2smsrf7CQwu9ndgmxksdJiQChT+Q3QP/hHJwUUMfDKLVE2rHmb4Z2et9sU5tjz6BH58PbE6Z+R9
UNLtWKRqPxVm1ujkFa8DYcNQyQj2a1Y6LUhUs75OPEWMHVtghkQiyD6EK8eT4tYlIqHR4qPZO7X2
JWUygv7MPntVzYmQxto2W0x3HdKS5qszS5lIsfzj2L9diZGzGAXalaW4v2903FgGtUqYHSAgXYwt
m4RBqQdWiOQ+asFWtS+A6QMIZCX9b3bhYVCrnvHpXuou1UDNjEfSr/PRU5Cx6GGcN85kEtFRcq0y
N4cH/ahKqtbr8iC9gzP8MElRdpFqi5GU52h12/5kD7dJRnoforqps5V+2dqKCAGaPIKEyDy34hea
pbDmbsIbMEbDk9CrbXg4QZMQ+T3yX5m+dTAW9vjuMGJ5yMi9ZLShQy3lq1cPZKPfCgfAcpzmQCDR
t3gL6rd+8ILFcbM36QApu0M5XEHy+3QzasKNOvpEQTdNvJHeQNU19Z1sK0/qSbiJyazgouj9SPq0
J8xUSZCWEC4TPBhyEQ1RHzE6H+CK/HgsN6CRIVPR1/XOFRghhX54LiTpVo0VM3WrRV7JIsUZgDAz
OCsPfL9095gSqRLbKLFZ4cBvRWbXhuaOFIqu1/X9h8ulZ4xbyTEeyajtW/58dMV1TF9PNod7t3Lc
5v1O2vrVBRvpdf6aQ4HmV2Dm+fYxpvEeYe0CK8thWlv7rd4fgh3sMcRZvqjt03NS35mZxFAnPlEd
9oLE/NB1ZfJTeQWmZ46kByIMT06s3ESyNiURz7UBwKDabKOm3N4roxYiuPjwngS3ec/VHT5Uy8ZJ
gvV1ELBb7vc1wLU+0yr4nW+5mNBn4UuGQgpZ+MJWakzBUHofDdlEBcLGuVn3+rzLqViMCcUHmD0K
Ex5k9Ivew2vivi1PCAiMgIRs0ZrOr3vEizxjXCZWuru9OTutFjsNwwQ386Z2XFQIk8JLa1IniDQX
ZE+swW6EFRR6lWDvkfEo3MDy2eRxJF0IKXIL6NCEcIOs1OmmLhN1Jl34iY4mMoSMQ+nPTIY42/6f
xrTYtiLM3RJbatXpcC5fkD2tH/Bou/d1F22R4qCS9AO7SqCwy+zzn09xjbarCqOej7HbZGlsVxyz
2wcmD8GVlMYoh1M8rLujKkaohLCLevqjq1OyxD4QwdY8fjAC+PcjNbR1RC94p54o6h0pXMlUMq8I
m4dz5x1JqEForQexMN1aKWy4kE8qgyc6Utz70RuGeWPIQBNaoAk7WrQzhVdGHRClm1LHHmJzCrW3
hSt0RnGHcQd1oC3spep20qxSmyK+HtcpKCGvUUrW/sIGfjbL7hXcypy1BHs7vGl9totfWn+Y68xp
M+hPg5Mkpvd4Fjg7KTtK3txEM6ns4UcwWZznY66oi/l4lLkrlnyUUDYMfYNBw3H8R8GRUAZqeJE4
vmEQaTdDh8yV0gm8kqCACdCNhYyehbN6/PJEH3Z/ahdc31X39/LVOd74oGfaqncxy/oRdeyqd5b0
PrU8za4EdCkDbL+mZK/5IbkmUbAg0fIcb7otJgH0MNi8fszRDDoZdNqdRALubAfR+JT+TQVYLQpX
RT2cxwZLGvOBGjqwy/1ZJrRHLIVUhoaWvsOHprFGIyutpp6VebXQwWHqZ6VvnQ7fgczsoZgk81YX
nZKtoRsQDavWQ3umUXFceLdI/F7hrOaYaPP7siPn/kvwzulSrf6w/J9XvQJNggwGSQMMGvO/loOu
N7x9ANAmFIJ73u/FFys1HPtyfidpN/pa6BQBkdeT1d0DrO/zv9YTMWuqAI83EoaIL0sMkKkETMcj
pyJ2sfUTCGVTDDGQKDhYJDyqqDuZyDQaBcxxg+97K8jMkVXT8dCZeR/9csLdq8+j/D2AgzsYCF9z
R17dkCjeyK/gW5Gu+WuyY7E3hk5FoQu6/H5OsZjt7qn6LIZna8olTBzFQ7HxsrIMOT0kkkpNZFBf
Icm8AfmpgsHCZQ8vwww2I6ZUVfvM9fkLZaCE3PRMfTYjJVkXqrjF4syUuXmoIEbFKInQX4bMf6QC
Hx3n5nhN8yjQZMIbW+6bFJ5n/G8zyrOGOP/6hxEQPakkFvKPLWiT1xTZ9MjJStw7DKFUo8pXku/P
r/vpNJMfmwXKl/Fd0RO1YBQtEzXeXjN9XZA+GnuoQmtRk7zsdITp8VKk9dZbaijL0QR1k+027I9p
0IdFPO3OnCGn2zjBPqwPxzAkn6cPmBBthHiT4b3g+PnSdCeRzs9Ww4NRN5DnhT/+N4EbACSLKfVb
1UqLV0FcGgXSn7WH5S9fiGDWNU4J/SkAoWQVgdsQB4fZH1BBQnwelBZbRz4c0u00lbdAQVeK5vNE
foROI+l0QkD0wd2cUC4Nl+v2jRDQYyWXbh1PRnnyRyvqbLE7LoTwS9t1eJkBAosrDZ2MpfYXrrU2
X/8T4+P9H52I1aPZ9bt3q9/uvSy+/9Xnay6dhdUHPrvRTnjiDsBEenKnJO2b5Yhj1E9r185NDenT
yX/I59IIFGQWr/iSw1Gbe4eju3fdsb3Zq2mz1ioZV6oVCQsS18h+1aIXsemYgkJCeI7jjEdUmgeW
s3tWuYFbyFhb10DH7qvbt/HS28uaYBNAZoxREZJ+Sk17m7uJUMalFA+lnj9xSNMaiczvLIPMmvYW
kl0wFS4v/RPBLlVZUtj90vaEClSwHi001Nnqhui+SKUFg/9xPGj4Gr2FTH+T6EH6gaj6BihPpZmg
89YeexNrKn1tqbYFLWBIXlnxcySh9UqNYeEtDfpqH4/6kwipSJSqsFKDs+JIq5uHssQ228MH4D88
iuO/XzC5MPkjhlvoMBzHNmdiY/B6j8oJ7rcjfcNFXnE1N32ZHX4RYLzfbWGsYtTaA//sCLWfIg4h
UFwUgugQmwEwB3nUDhant/0lmR/C6RBWy1gTwPRPNzCrDthkOl0RVhFugheTof42ozyWjflCDkvG
8HTm26n2Mb+PaeGI7dGk/3Xm15o9JOkFBnXLMMTMK/jNyRruwmzbQnwUuSen3i/NZ05cKHZuiVhx
C0WDkM5soGzfEeDYgM+VRjZJmlsAJOTZCDqs2oRDoMHhBR6WaTjAHlMCjE1f7POx62bbb4mCfTMH
XnvxnBu9uz80plMjhjW7QKIb7xaFYEbUHog93aVBs0x5tPMnX8b9dfTg6aEDkyIb8au/F2oH0Qbi
EJprrCxgKP2D/SfAPYB9QPljN6896Z6jOeqHx54QGDnwdcFkX+Ys5btZnG+9hcyiL+kYWCfKOcXh
ol27oy4qUtcYgBbV00O6m9hrJV6WX4AZyCKYa9IEQqw4VEUJR3Sx+gnMf3VvRsw8ebxmc3TYv3dW
cBB6wDhBZIX0tMTxzY0meVS2moi2iN1gjbJEWu57/0uyuJahdDOFWrOsJBHwkAhAnbL9ct/gLDot
X5+rro6g2WUpFQT6pEH8Mb/IVp+QPXiZJuIladYZKFHzT+1f+e7U/PjNHB/xjC/2M7U5zcPfQ5ij
PCbV1Gv5ErUVB0EJUoUJSZ3S7b4A/nB/n90YSgGUDOtLvN54qAnWXIJZsfFXWQIU818yfF/21nzh
lBI6KA6/lG0HGA67r8s830hBixDBnsIsZaZ7VyAYhSfmqxs3j3QpXsOcdZGmSRZNYxhu+tthYDoI
x3nc8DU95bZreXBqMBr088DIHPsqJuaxeHEhvkib3TrU7bMzZTRb2/9V4hu5kw3MAdC7zb0RW0AO
QYuQh3og4E2V/WYzPHAeny0eLukbehfMZuimXxAmLwzu9D6xabAgdm+SOHlKa9tHUcGNw86jlwQe
oK4ngXmtI2V8XXrBfk7dMbd3E7JEG5lPGXgJSYoqUHTEBD3JUOqMiP9EEMBAuEsk5uq9QPtcTYwS
65JZ0vnECXsK0tqYJP2891udbqXmxdP8lePFv/oTe8Gc9z6nqFVMLrM26arlm2hyZMWOozrM4KAs
1ev18epx3w4QPZjjNAt13hUTyFafnjNGhA/YiI78jmZ8P/eCsX8DUYS5LPlz1Fftt/qIMrxfKJ3P
c1GCHG9KfwGX3pQr+xd2V5uUJRM8tvQXrP1d3y8D/Gz0ALrvNV5SwRqFg8TvMbIH3C3V6lSObtNv
wcWM/V/n3ScqtNqHtdTtcB+Bl3pBrWne1vs5hKzNCYnoxoKlqvXFG2Ko2DjVCfSyuBM0EC89YdAT
XWJM1YtgwXNCMBXGnIPuWIQSM9BOTfptQlLyTXyZyt1CbDVoZwSg47uNqhS1rqwwblTmakIsWpN4
rH1JCftcmUNDTmdqtX0wOKZN2i0upLvCW7U+aPs5CwxNPO2BJ1lhOHVCMg+2CA7f8ivjC7mtYPaa
eqgS1E57nv7VrCStjecG52Za9zF+KPKKyMBf4rYVgdVwR5BfcFzDNBYz78W1+Tj0NAUPm2v3QCay
2CZGlN94/BlIeK1QriJ93XsTENxPgsBTBUchvHP5VXIxG4MZuNva+jk2vn1DOM4KNKodaSkpzslz
ZiQktILNujsBjrzTRC0Y29Lo8vxLr/nLawCamGQdJ8dqtpeK5E6oAnPdJRLQGw9kFv/IKZBUp6W9
mJdS5Vt/gkAzKwpAhAc4KUxIf4FmLFeS1J08fNwlcblYEBZtHu25VUH4XZAiRJ9zCLVL3qmHDs/Q
PbCnrQQqCneyc56Fpb0fmp53lukSymJMXpMY16EFeoisidFoNzo3Il494VvrxvYp/11HP/gEo2Fw
dZtBt4Eo+Wg06cCU7CFMsVLpc8rahddKgR7NrUgOOA3SalA1UYnQWnc2HNxE13lmt6XezjqwESad
e683ourieBBMbMEiO+TnZG0bvU1ovJuuW/9T4jyPbGstjiLklfR1OTQgIZ2ZADNFGyoNVn+nwipb
fCzqv2JocJ4HfrTpxEiJZCHSbZB4aTKVV8Z4SY03OUtz6UNy5cKKj2LfcHwrnxBoJA8DVfVqElMi
BWTklaSIiRA00SGIDP0Od+AIfP+XhqouUjDwFysxrETbLUnr2g1eK8sSwhpUEJFRJSPozp5mmpYN
jtu2xr+9dIGNQySER4ImQoFy4yHRi5tz9qo64v9slwBxxw2iUQGb27auU1ryeZCDtMWxZPbPpkf2
nky9bIZTJasmeryLfrYkCpcl+aNipy8MH/CBudsEstSYPjnt7DA1hUWieo/1vnZgJHNSZfoeA03p
1zuzncm9SQccH4AMw1iL+2o97/a2TSlv6ksStnjWcYpNSLarxk3GYinaqG1jfrMAfTfBrFI7tUXl
QkCLyhV4usbqSS5L5K/jtkTHQ7PVVM1VdN0HZl2R+NE6ODsz7gptQn+G03K/jWMqu4atVs/zHUFe
bwxByHxbrsPFmiqjrU1CLp1s+1dziD3k0d7SGMrf8Kvv6r9fOGrv+IToPdHJKJzXMYsvLgHcL99Y
HsLkv7Kau+VaJQKQOukJhbWDCDCv6J0vBMBNU+lw1miq0sYmDib0iYg1y+rATWvUqGuIjkMFG6Cz
q/vmkqlZKFmONajzRkjhWGTWkrvdVf4JPEcTPr6u0qd0muDEk1iFWikOd2r47CKAtQAQCsHAmWPq
nWyhzF1mHZniz+yXGnAYQ6hFeWrBMpKF2/gBy29fLVadWJJubQguum9tZT+Dnm0p61xpvuLKsQzN
xY8NEl9bD0SIYfCHgDdyyk++s9j3M/NKErydl4oBD/Gfulsm4SJqlqwsMw/xiFSA2grefNZM5FQb
aBt/uvz/geKerlTFUOV3xjIE5LGRFPOAAvmUZ6F753c1J6V3ITtfY9u/odR1EnL4txiZdCqSYzC4
1qZ9reAQ9evZSIzIioAzTFME7fpSv0KGUIrLYkqLoIYJivKGcYKF0TyszkBSnpAlSKFln6il2sbx
/ldynWekFg4PQoEVSfU8KBdBSzqSFcj2Uvfn53Flhmba40c4UyvYVE9gRbx2Lqz7dIyKvLU2z3Gu
0W8ss3i4Y6RMTWKLTycenwIcFlChee/+TV8Q8Sya0PIFhGY5hS7hUQME86/JEPMN7uTCGzJP0EMD
PeeuzEc1e0nxXc/Vz8w48PCCdi4Ak6sD9gjdRHT3vUAcS6+wilBwygVLFG0zcQdqZlbwPUQvgxvw
qqLOvi4GJE1cvNIYWhUzfclzG8BkyaZ/yTlQtPVXFuRk3K7Fv3FnKlCMrpTtwFoEaHHJ0Ak7o8yp
Jggn7nIldwAXTKVuSsZQZwmFpGkY7HW/VSrlHUvprPV4VYm5KnSHnJRubJk+x1s5FU66KAbpwR0k
qms38Gpjbb0HlZRYUiZTvyRMgsyixNFIH6ICDHL9l+UNDXH5E9aGW7OqiEuuSsWu7RfQdGDskRgq
lqtIK9O1XeSff9+XzTHWUFiHuK69fpS3mhUT1estwsMjE5tyCMeAugezYUFRMeCT6pBRTQbnkVYf
JYcRae7GUdLjFscfrJlerMk8U3f1GFDR0EfJQTe9kqYhBLe4Xno/6s6k+McFXwDcSa9/58lI2/y7
GnV3vY+EMPi/q/EjbRSFGaFDS0X9hzkaeS+CBPVReSTCF3h0NiAW7HN2uXlbz9WhqhlwUTnuHVyS
6JDHYYlg9I+U66rxEIEWVrlZvS1hFc7Ne6JlLwZBv5pV/mOWMZN6zFg/87CQvrnc9ZnXdhZHDpNM
/Iq5+7qFTZ10j1ysxd/M9TuCHlAUmMMPGFdkZK6afySRz8IeBl+76RM9ZZU4nkbTnM9cgytMjhlF
DNdWOVb4xLZ0GcUBDER+KQOks46HhC4qEmVx69M3s47yb3zbsZOTEy6+m7Da7s/K7L9Zq1zk/aLu
s6PZ6rnG21xlJS3kxSM4ixieqVHxFWCNQcn64ndvfw6lJy/3WiA8TqervGOX4WbRa7gB5V0+x3Y6
/eQhEwByfWxcRmEMxJIGIXc6jznt9+02QpognQ/Pt65IzWA/fOEhchvMuZquoXCUGrmwEZAI+uqb
N7OWIqW9mPneZX1nSGTep5FG+oIVT/oMLs+pgWZw8Rd1a0rfyO27/skj3mLhtEwzPvHMwxONBTSt
YbWUSd+z8u/XmRWCniQpjgbMsEXhGSoY+9Zzt04lL5Ofjpa2ipNegHimtKO2m6My+AR35E80o9jn
yDhZsXJJjQT8TPEJdSy4YXC8nJymVpKu6hWbJDs+5fOvj0BzkNaQV6YRwt0tAdsFAH9cAIICAX39
YYBO6nVwkEI18IaTfh7xDke0JJyKy06CPG0p1LLSW9ZMkYqIHXeO4Y14cVBvo1u08S/OOr8EhOZY
FYTRZTqq5WYrPcJ1E36uzcjJd32+NwZKF45rMUsp+/QMbq/+VZKPxaBi5WoXZafv3RerWw2ru2cz
egU/TasnVzWVEAKjIrJ86XsHzAvuMWmCBkHf0gHU6abuGNX7x6D51dxNGIEp3iOfc/nsQ0izADUR
5hB4xxxpfCvbDcXJCDLE/Jt2aRX1EaJURTrxfGPu0/cBu4WCko6I/w69QLazlXCOXfQlWHqYbVft
9HkBxWR5OwlY/2+TrIdVFsy/DV8yJzvM52UfR4aK4yJEbf5a/J0BC5r2LsH9fIxwulT/fRYrK8FX
+8ql1O0Nr24TRuuhRvCLi5jzeoTL9axGhBGmi2csl/aeazp+ph4LZ2ViDSWsDgUg0WAXDU+hGIo8
OITQ7c3kCq964n42LnmZk+evz0UcQ43MCorzhkbb7Z5x2phH5JRuEy6udedGWsesX41UFfEx/geU
IZkq5xf1gLEcNKam+Rtt1QHydvnQNzDkdDldQfs17Wsq2jOQ0/b34lUV8LGoERopmo26naYctHBj
ZGSFfda0C+mgE9pExtpkJkLn8GpkKqGqHiFlqCuDG0+JlvTBGdX+j2AqXz6rJ40UKhyqlLnUD6ZE
7vh4ISeibIPvxSH+KdRUArkRImINpZt77u9v3D8m5hAJ+go6hZcNBfm9qjgrTiUrKY3IyGPWwVkw
exP3yg4VF6f0GP7LXS45Xl4Z5wlWvGZJP75t6G05IZXO2DaaLIltoLe5UaH/ruA1dz8U2M9bUadq
gR4gtIF49nd3AOPLdyk1mBosmAmqNwD1WL97E+gS6jTHN6eWtLKjgVQhshXGPCjpyKF2OXOF6UO0
2txHKUXer1uvMnbvSe1jkJTtWT2+D62xWdG5SG6CWU4RDj2RvO/fyIsWnWEqXcswChmGwQQEit4F
3tipEpytkoY9OgZpz2HbSUo48ZU7fMCOaAEsDw07IllMUeWg/rLyW94zDCXy5vameMM3/JzQRlZd
0gUyQCm99BVDgXR47w5xv6xA78EdFjB9sIHMlGtLSGcTr981FfeLUSo3GXYvkpvzRPAhnAOB2MhM
4AcA38k05GOHXKbNhBbGPGzWSPSIbzHsR1V/14YuyfZEoMZKyAZd/iFZA3hAQfZ+3aK//VIXnGod
hVvkyiV5rJPqSzEINH6ii67RFVdOwNgqw9s3dc311jRvy9Tu6TGbQtVOlA8sO/KKTv1x38WwuEqp
4LaJJbhkybresrNP/xekmW0InDZIAJfImcfRRqI38zazx1KeulSKu0NWpu/SO335OGF5HZKczhRC
do6vhDtjCGR64EI4XOQAzsa9o+swUvIKaYvHe9Mvf9z9ABFC9DKcPaRBPCLTF4it5i1H+vY+zxfT
PD7/2mxTmKTpALGriaNoE6xBoAMwbXEqb2n4gaNpxgRuddGpZYgHZAlZzDQVBSdIK0hIEav4LSHe
iwSCWH86P+5exCp+pDpV/xwSUIEL9M4QAzEdOLUBIZVVlDxH0kr/S+IZYgG0QinuNHO49FQjodLd
sD76XaBmBktView6muqtGXBCqGwScwrUr7IZJaTPS3SDc1hAoZ7ofYnRNHcV1s2ONOzQjyrc6nrZ
7PE3BChSNnqNSB58im6VnFwxw6XJso9m/9gnPJ2Ky8wEogd0RWysCs5bgzKEINgCTyXcyePVE8Z3
dTusTwjP8rtkSTFEEAMDCNTmiuPf9oajdu57lrLE+yAt5AGAGRrxqSGXXXrDJEgStD/2Dv5ENDBI
gwhBhiC7v52ncM41GmuidVMebMZnRaQqMF5hgLpyrG/3MHSRjAlBTr1flAngeY1e9TputNg3xlQo
pgiUOtuIDBEqBTqSQ+MoF+0AoTsQ+O1dnFAfTxxCd43em2PHvvqM3TGakrPOYm81FM8HUh7k4jD/
ncrYrGw74/h+soQB9S2ARbjP1nGxhXN4nHy86qZ5LeCaCHhWfs+vKMjNa5ACbyQkNGnX88sj8zEz
nsSU/tjLIayC0Yu/ZxFNqBn8N2vasmguvuenY+017CHE3bH3HLilu55JA/JR+ZXvUAQVDO/zB23D
qP6CIzlLcTpBRwwgCPgOll3R+4NtPczC/E7yfYbJy8t6BcZ4DFfjOcztDKojDIuLq+8X89WjOdYi
t1CGyXtrNEcPkNc4/fCmx43MXe2c5Vn762O8Ahg6AsVmWitUDuE0UIwjv8jrYGxIMMgDapV7Hwye
mlYwuTMjlV/Z9jrROFtPlft2tWbalOn/CDySEtD0JHFnQIj2OVNuQ1MO0/iVXJfgXue6K2oEeLI/
MY8EXqrlhNf6/IejsjjWuCj3INeUAEKSiMqcBD1xrW8u70OuXDHabU+xUYf20wXz9Wqx9l/lerZB
NNtEd1St299eammPg72fHDS9NXAqt8UlwtW+7/XVNaoifCFUPLl5hZivHkYuAKST/2MdXNyWxzJN
E7NdYRoxWd7R53BDnppdiyiuaoCgecmhFOo21wEU42B5e8u/tRfHNqjE4T5053EeMjdJ3z8t0f6v
o5Y9Y0y5bF15p+S2QZb+jNUvC+BPy49dMfUbYkD/GgBEmS/wAPBNsg8ep+zICQPTTSsarAmdLZ5Y
upyrIN/LLEGwG67LANDABXJbc0TO+XQ/CofIOZTLVnyA5RcmuKaIUoAOdpgzHRI4AGtEqIF2Wnt6
hR3AwfGZeyT9MP50fJSivPePrK8k7N61e/a6VnaqPBAsSacS9RP2DluDaoMdw11sHVaxV0AVHQ0B
JzWli26b21+zY8ZmCjBkjPYRce5eOwpOrugzyGl0q8l6uEgb+lgjcbBtrczEwqb5f8niHC+J5esV
Dvt4HeDQTxf+yuCj613yiUuotVF6JT84I8Ha/8qmL1gdopmVrOlRLKCFBlVUcNXupjyqVAVx1Giy
YMs2PnqPfcI+L6prCjICerbOnEl2T8/kWYG77+HowR1JoEx6OJrTufpbRc3j5Q1S/TCnTdVIGzbi
ul7Jn1qRZTsBn+hIP8Sw11WRQn4L+6dXa2KFrtseek7UhhUVrd16nC1Ap5jDhdFsY4MwPF27keTy
nas//lyOKAURoiin5NxhC4vX1x2NuitUhINM/XQdPIPdbepJaBHHS6Ovjiv3t5dxw9kQSErDpRsb
k+1sN2BacwLoDdlut85oC2lcwNdBokH4f338RqTjy/hefIRkdcFSLcmg/AdmJHW9QyQ64EhGLX8w
DtsrInPDQNcNdnfxrQ5G5KfexbyFSuJVpMHRTxY2pa7rPh5e0rzIWVhabljhPSOrckN17lanbOhF
7wOqemjRJo23fymp6yip42xV8lu/oKOeecJ7g92QeeKh+bjdyaXQKRJ8CV6c2HBU93H7pgh7/sKY
qD8djy+rpnXaTj/FOh85KyhY7qp/pZGYvmoUF/D1bCyuXGXPfJBNKSmTgqsRE0pI9b8Npl50MjO8
d61FIb+1wMxv+Xi5ElJfHeO8d1LrNOPLByWGLFFWWSM5JCjOUEy2kb4aC//L/U4oI86pfsLmr0TF
gt7dZK44llmQIRml7WddgnO6gpBYfT8Uxqz0xysPedkCLbVC1a9nnMSyGdq1O2uvsT6Su7ZXAgAa
RVs7hjgtgi6HQ5+kpTjea5JRQ8dqfM/5/TPhTxCG4AFBafHFTCDHT8s3g45nli2TkXZkGJGWst25
fjV39wt4bzixfbJVtk/bLwwYJU1+FGuvTGY2vU4a8VvCPfn+9PuQyOKZi65T9va7tEXQluBYv9vO
mh0/CvLFCaQlQRufzW7gvjXWPOXZ+n06DIM5tR9wTQwjrVePm3QR4W0p1+2qqAo62W7CvalHZ0EZ
lBBNcfB9PkXqBwUk61VIkio9apeLG+FnR2RkAmN/W72qFKmppNKiwATsoUTp7qAakT3SoWds9pot
+QYbMQ84kiI7bCGkCjQKJALHiYZl2sxYLbi+ty4KVRpJBZXefceFKuS4ovdl8r6Mzc1o0ox9LTPg
A8KgNDJBTGx4g1Zm0zzaVzIL1hx0bqhD0uvhstQwK0xOiHp9yvYUQM0qn+CIB8farQWY+0FW2dgq
BnXmnpIvWasXen7/UIXAdHcNUI//Wxt9MEYq4N8WVGYrXCprvDtHNDQF1CrMWyiOnIfFiZFDxotl
WIDUkeTeRfElMH5PQEftqi8qnNulRotv329bN+Z64zExp9giwhEtZVwPpcS5rUIeAXlkNvPekH+R
PieLk9nlsXjOEtRvnrEedhcs4JtB8Yn7OLQ+d2CVTlDK7N2qo/tqL5ULPn6YMegDbMAxGgjiZWDI
Q16UDBe52Htkq2M/zH074pd9ERsFFE+col8hrDJG2zzia4PxgTIz3NSqUuoux4LmvcV6rQTsanLs
KeSDntHOlUtuXyd9f3Ehcp+CRJzrkgAq8sMTqp8SoHuGLhOo+L1u9Aro5YP+r2pNVoK1FEgAWAXL
ppaywzac+dKejxbCwIBk70mrLKaMYA4QdPLonPllplgRvvpsCtWZvseCGmHXLlLI/n+Fvls4Yarn
40TcggKUpSTQs/+m9c3XJ3rqOngC4L0omUoOBTDc/mDsrK9T0VHaUoaOUB1CJZvvD6RnoAzd7rad
jRGyXYZSmCee25N4UU+4Aiydm4dRHaB4ZzZZEGWmntTUBI3M4SLQePLWiRlPdPsL94PHCkQrAGty
GA3yS5XcmhO/0zRDAMr0MOtfgvHnJmk53IvrCWtzjtApsxkdo4g71p6gju3X95Z3ylW9y8eRTP7h
bV+LQ+ooJTMv9vjHZTJOjaZDgLI8jxkDsXbGuOQ26szFg3AV6Cp6x6mttB/EfisEFuSaldHpxsoX
jKhRGKm+hl7GfaIUp5tWZCd5gdP0sbXBamx92w3seRNdzv7d7v+/MGB+mYjHiE2+L61QQlu+dXav
KvCbf91OAXU3lCW0F4EOW7lJAp8yGGd9DgZpkcDsTB6l7d3pefWJEEVs6/f5apUt1Tb9qDDgEaTF
EGfMaVBKRnqm8HVmlCpw5mJmtiZEEDr2dYfsioYDbNnhT1QYXkyBQC6A0zCDO8OwlECYN0Sci+pU
B/B4t+3XCFYI18xP1mUfNnv1EdM21Aq03/0alDvhn5DSw+7ZK7NIVJE/r1nMMnu/GFwaK5Wzs5Br
gDIR66WmM7Ui8Q+ALS0N4JRiiylyJ3VvggdrHCqI/V9hQEcQVWVwMtzCfiGcd0/WxijiJOQjYT81
zepXeptyy7afcBezAa+KpKTQ3pv5uP0ZEdZ4DURWV75Cu5zs4FRFRNdGjFCuwvB5RRrFrTR+vc8j
GwlF1exuLe4UViGHHsaaIAnjhJfWvrt4WC6SIM1KkZnXvGzje0PvWXwxCWQg5qQmLCEPFFhRodod
sTQhEYzR9g6Adwwq7KEahhCNJp30SwgDAb99aAMoJqfjPObmY6CzK7qtciTWg0EIInKYSIV7QhZp
KMzFf0kH45OqtUENC38qzEB82XJWs7a0CnGtUAhCLsv01unDU9ZvPecT6y4EPCZ62dtYQZP7/LOP
k9CFFmn924MxINrOOUZEdIVGJ4Cfh0IxKBLOopl4iki/a9SMAJfgChzkXN57LOog70WtWfqckFDt
N+ra4mh+GPcf8gxFi/oqExWtARAOPXk7B6HYvk1tXZtUqecOdI/ZJkBph3BE4jxiJdN5dTCz49FT
dPltAzhUKTfWPg6lPqr7wIUQy6x/7HNU/4GdYjt923gnqoTNQj95jzWx10lvKqH0sp8ZaIfus8o5
/KoAZeo+BjS9PLy80wBW5W7/O0KezYlmeRU1hcpqzNJjYLgwLrGWqjUiBjCgD8YNPLNCdZMk1+Rl
4MTIhQqptVFfbPE4j1W5X/wng8DLaOUdJjiU2cf/VCeas7WQaeFb+auNM527r290lw2rBl3/5XZp
DnJYIerDshm10uF5eTmX6Om8Iuc4FnwDAtN5SInki7AF+Kzv2ESfbqSp4izH5RneZ/ZbC8JGcbkI
EvcZP9Cc12Qc+85kAIwBYzRLuzj2pgbOcd14KPNkChhDNC6EAIA3m5MQMfmLtQxmPO2xPCDaEpA+
sUsO6/7fEnpqY4dhhJpYMI+jCTks+YWLNdcRh+WyfXLZlUslgOIGODM0XwistNZLmRBaFM5T1BDb
XEFioWp/3CT+YRZ/cRR15fDOIFisaWKcznD/GCW1NfXDz1IAWqXRDkCuXA1qGSXw1LtnyZEiAhQK
0zMHIgjYYLvFn0BkDmAK8QM4o59I8bsEbUFQYTXLrTVWDu31wPLl8sAUaF/Nrgqsx3Fl6x/foNtt
zw+f0FHrMK/p2Kw5izabzdWnHaju+KCTYpj1jMuSkH5cMlp8gUNUfOxRBRtJ5nlUEk5LGSG4tgje
rEHOs5ZKBU27y5D70DZdiejmF/v0CYpFg19klpsGUx2MjxXYWU66bwwzvqOJHo7RImKuQJFLkkRf
yWUEbg/ypjrfcHxYE8e/x01rrPESsRH88aOnNSRYpgznXZqB7441thDVNsSScZkgqYBD/Q3MURI/
nQHSyA7HK/+222B45T+IxqTLrYu7vNPTQM7bXCVt6cOgA/jSnKWKwWcR57jxW1yy5IrwstpK10z/
wpDBg88jmbQ+QXTUq1R04dlx16hgfRVKSzW7dDcMHtYCB/F3dq3ch/2Z5xAKLLDZ2Md5JSAbibCr
2WvM3L4gVsjSl7xzQZBJ2p2Ea9FkkGofNnFExrprqxGCQunanwKw1Rx96ymbjed0HqW5I9NYsFvq
LphXWyJxGkiEWgTdjQC0Xkkk1dK6aqyMbdjzIrIpLnX1VPGjLvLQePUp4f27sITPSUvIys/+VcH1
01YRD3Z1cZPj93QdSiLyj/zOfReOHdxHRN2YKeZ4XpGmBlXpvi6muMR9rJRh4LKdNl0CQf6cgWWd
+GM8VpFgFc4vEzhl0/aDXAu1w3M8aOM3c9nhlWo093jMUldie9i9icxTbFbi4yKQd04ipT7v+XXm
EtJ7Zc7515b/ljU3foMqFfTwKznWm6XNKkkytArNoLLcHdQSEYrJxr8Q4QcrAIRmjWRHLgFBeIud
hkCOCg5EhYtFk4VHP/9YvlaCkoe/qX15qpqON7PsxRZyEQNzCulmOZoEdUuTCkjjuCCtchsV5ErM
TGZ9bPuXQDkzF4AzF53n7y7FmZwdRdLednf1jT8T/uUafap15wHoWOFj7y7P3PYbgztf5X4/sk19
VbII2qj7kV0yLd/fFFagjzfzNY+4bSfFONQXNuWZ7s5DZfgAseS/SMFTFbebP0JxTtKFdJYEj73H
7KgvOh7maygBZEEV+bfT9Wg5NqtiaBB7K0PKUb8uL7BSAGkzzszdkJn3BuJkHGMUqddE14nySrVf
YOiadypT3NLVh56qsj3WDvzxOrEkoauXQ4LiJNwd4YKBMNjbeXgkBDM4zGpWoqL/t/kNc2HelqqB
26/CTZjA+kHCMUdE3q3iIUzYia55umNcmx+aeaTRCDlC2H2aewsLtip31d2iKJ++QMxH04wQFkam
lYIvQhozN6Q3YY1F8BPdic+ZnIxV+ucaIxZDTjeLkZ6Kw1VDaUkYHp1JTCo7+GFIe3K/yYiluvZL
Nfv6o6Q0r5deNfb7+A3r0drxt8pqEW1lAfOsqNJcDtkm25eylVWzc247RaXKJ0rj91m0K6v63W8/
yCFt24/lpLpBQ3ay5/T1vYF4xiiRPtwbVZHrV1ljgcNB/aoTgFOpm3WDSLGoo2NOhg/ZGa7vM1wx
40qG519UA3al/RWN2WThLhzYQuQVwLibOZIyOe9l/qryvBAJOEJZ6zurb8+FAIHw/NU1cBG8f0zc
plKMorOFCtEI5SpkmNH3TWAc1JV+GVRJnc7nhFD51AcEOzJZOssQXsEWC0Fq+yctz2tapZ0/o6Ss
JJoH4e2JUbPTZtcY3wG5o44zNs6Ky1/fMoijxc5Oq7vgCHu9h6ploh0JYrZIWh1hIaa55Z95uU9e
K77YcF1VJ0wJLDxZIGMgjiE8w9ABpLlcovSbuj3mGu9TiLUJXkeJ4I3WPlQcd81W9TmSpewNTfyT
9fflKXIvqm2K+AwfZGyJPftgPm/2tkU2Er3a+XsGJ+1leK0JMHxT86KY7TgVa5Egk5N5V9XqOXP+
q3gcovskRMkyIrENrdWYdVhQxJ2w1PwV798KU+OquNC6qi1pPEtEhnoqc6E6iyRDqQ+RPWb++XKv
sVZKn5RX3Dppv5nwTakBvzamvDvKSksttZ0iNLBcQq22xKuU3KDYi0lUcGOTKS2hkdR5KYwAl0XJ
mDPF3mGs31Pa9VIVwHoOA/tdeVuIPq7zdOxGc+uEK1W3YhYyRiackFXFmwZkjbuj6jbh2FMzmV9G
bNrONu81Q+fp2HFPcPogy5iBTJ1us4zYIghltPrxPO1/UHN/uXYZ3q25ktXuPgZZmGckmLTU0SZB
YEpAihBcdtyMNEjqoM7vlb+9xCCpY8hlnrgp+QKU2HZQiWwnEruSoSsswEqzo7zcKi3ZbtO+ARYl
JcaDGOWXmSyCGFpg5manDvPXUaebzSyJay+2P+DEVVACadzE7JOGmyYAjPb4HPBM3zmpVJSj0KE1
4sWr9OwFlh769LMeP6+45p3yPlL7V/t8iXVJthWfFMHgrY90FrgUCk/KUljJDWDjQy8gzakiZJy4
AaxBAs+7IdqXfDETZtTb504h+5wMgbHoKYGqhPePZMsPLyrp4bLwbpnCkLhLl477u1r2wrEBjT7J
iqQOiyXp38u1lo9IfgrXdxFuOvybaq4q6Q6LV9Aex90Z0fqtCwdEZiX2Jz8/nNpecra9NBE/d3Uu
ByeCcawUpYk2B1G+0Mgt5pLNHqs5n3VqQcUs4qRl3WAOICj/N9BmXrGQjFjdZF7ZgsK23xhtd/lx
xuCpGImyh8NY7xNzieAcJY8Bv2yX3ICDlyNyAau+oH/7Q97w52DYu6DO2ZGiWaRI66mLgPTywc7d
xwIcQKE7xgcE+4uDightqSkNf4mfSSFQxzHZZLBrSlUoifPP5E6JYPeuBylCuH+sTTJvB6quv9IQ
0PHtcJa7sFAOOKcYkKoDWCG/l1h8lxuB1BXxORlIdBoRQ/0h+VCwUdtbDDAtiHeISHZkiR9cg1ok
745KFxoumTQRtUjcNoO3bmdQS2xpk4a1DiPItQnc9vl8WWlMAOuvcxq6vGkDl/pM747QtDHsaw4n
dzlnPjYtYwSEDhsT3N+lxZFfpU9XHyHDAhRd+r2gZF+H0nQTWwPzCP3KQk1W0hM2pb/WdXDr8C6R
e4f0Db+t+Gg5a3sVyjBLiOY5fK/xtSKcikmP2LwByotSztw0peiupO8WP+uZRN08Ix+wXW+9nvL7
gbnEMBpLFyOdHt+P7hqUeyZe4finCMTmvoRdjXAk+rZuvkhllgJXpOJrUuW8tC73sBpEfGkEeCCX
5NwhBkRJ7wdAToIZBK0XVhBYKRqC30GsLrAARo7ScA5iYm4EubcDJwFzGAGQCYNH5GKDV4cetu1n
u9NU3xUYzU/vLHqkvx/0FLQZ+tRmA1clRUfL1TU+Q6V7/leL1joDPGmaZEbsCWIqUy2ZJeT4s/uO
4dfsVGepB8LMZiBLIQC1qtILA9cHZEsGTOJeygiJv9WYS4dqWTzZuJdtU3ejO62alkOLvhHDjGKy
ow7o80ZU29jdG6vLMgBQyhuQGQv4bWtqNdD+juy82vNs0M8m7Bw/+xTGDDE2gy3nXgQJt06ZH/xc
37VvOsMpFLIpo0uUYDu7hyfObto3HkRJCbyLMgL/HAPk9jruhv52rmPQNuIcMAnxO+ynA6MXvOuE
LNIO/neE8WqR136sLuetdHH6m40btwUBbES8JR3IE0WlHEpAkFal/hUCJjBu+Bj9bW5nFIS9VGJf
r0FTK0vlo4KFHIAfEkKB1CGW4k2HmfUu65D78bJ9jajR9BKnxNguhmQrh8Jw77cAIenUhLst+58E
P/YrtgCUNZj3wkgzqqxU8aoVev/7QThueJct8MDvBEybcWt1sqbgAF3b36v1pnQZ17GFIfb3Hqz7
kQ4oL66AjubPov57eslPT/7uExgk3OWpcc01Vat0T/VNDYUu8Z3RHzRjkZuNFLOe8nRDEm2RxBCA
sfTyFhII/rSt8xmS+Q56xuPO53X0QkGHH4p6aalGdt4AZ9KDlTU3BJCqJDjmRqB0ghGVk47WJaoY
4j+JJTNM/kh0qeCHur7HVQnajo2SVSD5KIO9fZ07s44svqoA6bsdq/rtTc10UVTiOIJXZ5LbNpdJ
NCyD+UL14Ym1gcLaRRNfipSXESXQUcC24tSZTgjDHsj38krzOcChynpf6dk2aTTBZnneIQnVDDHo
LetcXCi1gpRIoS/Shxchz4qiEq/7XDH6Eaj55s1ym/QvzN73WViSNwKxKy5FUaZKp+QfHWXTJOMC
Ov3fwHq3l82UFtDtb1SDZdd84wy3l4W3sZlpjc1/lcLMnp0gjHIXxM19T9yPP9x8Y1PoC6rGGx27
3f7QPML8YmPf1wt5w7f3y2m0VO29e68eVcgnbrbT4s1aqpsh3LgANYwShTqTTDZfYrrofNU8aH85
mZBbrG7pKkgcgJHyDSUHpRYTJrSJSW+d8eeDDHrGHukv+6i2NixnD7gKtO6x4Q2FcfY1qZQ/6nTi
lFikJzHaMcuiX+BclYJ8XAkhegDpWxX93f3o9Zbd2FUCdzTW2HXcOgjG8DbfqqyOO7B2m+dMrYnp
Emhgbxnccj+8VTbxTt93+ErlfA3jP6p1/xNtyQVM5lPb0ntVIt7iE0AsMroEftzdNUnlldkHNdIS
K194U4KUTbsGdN6s/Yk16rnvpoz2GMvlRndT7wX1GsF01U8Znx1TKU5krX6zpodZv5TM4HMYgz/c
L1d8G+WDJchxzoAYTPS51KissyNgdc3qcHnCpYrDKZR5b1oNzWFDl/Ix657XO+CQuHeMNbGf6Ekc
mfoV6lrF0PqmpuW2h3+/2iDBnxJrn9hir80JX6Jdj1lodmmp5/jJhtRc6gDP3D+QXlghB7DNZ5SW
4pwuxnStbx2Wq8ZVFJhmwN93yh6RMcXsd2TLprOZR6Qe6M6lV38L9bcrRol17hn7lPd02lvj5CXv
WiDJh0IaFGTr3Sfp0dR57RpmZqir70tzmpKZ4vvGSotrM4kT6HpS6UB7fDL3As0g1mESv7ApbULZ
jeRl6pVPutiq4BGsD+mCPOQBLHdkydFTQfysD4o3aeg0l9j888icZsVzxrlAoncImOiS6i7zN1au
mxzFukJj3DZRFwY20C9jVTOSiDwYzrlhNu+CTr2f5wQiBCgDItWMH91j8gwLU4ao0swAlTIqd0H2
uEuQuh95wzXE9K/rtYHJ6A1E6hjpWc+wjByyQwtfLsVGZa42iUAPxKcUm+1s8vEis3bKGvX4jx9S
LS2kxGMhQJ+CMt0aV/5v7hzjgGiCXaL89dHx4F/SRG5CgerNo++/QS+FQXXRYgqmcgnQx0M/R5nS
D8yfBmDXNF2hWYilH1CcNuwCPSsF2OxPnfnB3cEkZ4a9FQ5poPU3F1/8u4cFXDqWFMGGDskebdh5
SFzYMV2gEkpBCI0/6VZhjHmKyXo0r0mwrq5eJmt+HuH+7qh6O9649Kq4l7vvEiHzxtF+MKDJuRiS
IzuVH5vjpzK/Dr5fv7CDPSydhMaLkIeiIGZIIJ5jnC4UX90R+sDT6+En1Fh/Ym01cuWy2Ouz0qOm
nJMM3t/4sgzhhJGQUqoXfbEpodt3mLBCBKdXJayOA5HkzYTmeREpttXSxZ7o4dwLCrxs9uuTqMsK
hzczYBuhUNXwwO2EgIgHkL80Aud08YcaGN9r9Gs56IY4ppCHUwkcK7o657tVYK76cCIwilVd7np5
sMJaS5x8gEebuxnCpmg7wCyj1BTwkbEvetYFqjPUFVEE7JGW5WN3v/SGkfAAPM1ZGF9A0jhOWvIm
nzQWD5KDkwvigdD3LfbCrZtQwqJw6VG8YSWc1IqgrxoepCWU0GcmzDc1lxJTTbcoaQVu0SI1PGxd
BdJnASsLcfCxGKBUJOgEQG1ugXbrw6zx0x8/FoiF66p2xijrHi0MfA5WgOD14nF1QDZIsT4hxaWM
5ippL9OWySwLfnOsC13Wa9YzxsqQMyva3ROPBbGDwut8XGxrP5xlPb5lKOQTjp7X0aB2Ljp6j68k
hQ14ap7QsW124dSMn0AyqbknDmziYAWzJN2Yo9WLZAQSd+cL8qz80jGHF6SeD0vLcMiQNqWneDfo
bWmrvAy2lb6z37WHSqn0fV6TMzObF7f5tzPzYLo5AOdYl2v22lqSPmoehuCAY0Pk1FoUiMlQsLI2
7bQESAo+U7Adjs+FhytzC5zn4ZbknEuWEb1S4RLgFVvww3d1bbmZtqjefcWmDajSHgup5CKkf5dD
qoWMVgTVB9wtgwqx5l4fCJNE2PvPeM9cdLwbWUi5HyvKqkdnlTV2nL071qlYs3jq20fVApjODqMv
dj1bxF2o/rmmssZXZIg8l9sex6N3QaZ5CCB1dAtcby7kNWdZJYqMEiZxPTyyJmYNf/bEoiyMqW9j
k5DpVds9wqlz8HiZYDMT+AErRL6N8BQMgEleWssD2PrLdlRGrRduSR6og9O8wLAoHxfs9FUiU4vX
SqUDABp1ghWT1u5IPEVO4yO6jq7Ur69fJV1gEgjrOFmVRBoCKyEZrfWZFD8IO4jFDvt8Yu2LMk7X
uKuv0jkll7a+PN1kN/iqzgXNvI0Ni0JfR5tAcEGxQ8foIZDvCquwWnUQ0dzobfBEyCe4TR94c07m
soh2mWAiM/SII0G/r/y5XdPZL0zTbRYun1jbq6cIgJYxITnQmrGKj7k42Dg/GFGrGgYs4An+/+0p
wr0sZVJGK0fE2TAl1Q5KaIDQQcybbieS5EewyjD5aqmJPlYNfuWksBX3i3FwO+yhmAR0rhCUTI2r
pLrCnb/2UZdZwpoVY+e9XjdU9AwOA2i8HAKbPsEcqf8+FexgJmezexs5y0fQfnu6IX3ha2ilzDjC
+qAmlc+3nPSN68rRfhESzUKQC8l6cQKCD7vlpSPBhEuF0yRe4dA/e8OcxMeHwWt+z5p5JLlvGR39
hVSz6uSatrXc/8PUnm3Z8MEaXbu8Nr6J56h8TpyKCq7QT2Ld+lRR6e2HekL/4FjlalQmUtGoDPIr
c9xUaf9NAOP1UUyESvDWCN/FLEBiujV5JleTK9H1kJiC0Sy3wtC1KIZNjYE0k7NsXfO414+aLhHs
kpOl3/MOOAtdvwffxhTnVnUu190kA6sA4BVdFwCLL484g+Iox2DlT+2yVaOvxetMqBQUGdGa3H3e
kamSs0HDPUGpMxzQF2tNnqxIyxSQ6aqqmlK+JZx/D4brcT8yHciX9AksJSzsQte5drLmbhPqTx+r
IyOSK0MbZ1vljfmwHnEvax4D0MO8yzD6alYJSC6PkIcULV83XtDWk6Bp2yP7C1KqhURgoqCJie8S
15gYnNuYRYAMhKQSld0kJT6QmLgLdWrM+/vflWtYnZiYxkOCTg4fnt+zD6qVb47UtAFwC2GKCpQM
MtlBeqT7UosofqjyKPH8D7JhXcjhimX0viLngQukWMiHZg5i4wCDVqppczAjxt7xgwGqVS5QlZ3n
WbDnLvJ7aRDBEVUFjD48oiexdMkFCOsvAEcT+rJE1rtwd+VCFaSrTEAZtZhgG3ZAWkwucMa6sCb/
SKR5PdetvzPJooal3rLuZoFqDLK2k8dJ+Z65st9PGpOHHU9KgFTzoTHCHiUC8aITSrePCn8zjPBg
oVsHd00kuF2tBChvQkM5deK1TUhAD3DEpboisKRGyJKX2Rk515HKeLhockZPYRQQdzL2TTv4pk8n
tfLOB0Y+VYcuULcQUaVUjg0Tl7gK6HJPl+oMTH2C1ynKhzE+VsOEvRfkm+PIm9Fb1jFoIiFRlCSC
aEJz5BzvhxkfZNLOdKYoMv9sbsEPEZcG4Yl3JYcooSFOHi6ig9xzn/ClhVV5udDcpKb8PfIX0e9U
Vm23ycsaySVY6rxzysgogcEkoxPvCNiIBhjHGsv+s5iN20pDDFc3fkjvcmJ1S9o0hfOrwGnqx5a6
Gb2lJSBQtSrAigJgq85dv9sYtxe80A1sAEY5r5NhzKHg5z+9WXhqXdi48qvTTTx9z4hDK2da1hud
pYixxQuOEiW/Bx0XIYmDPH0aSfpbcUv/+SCKI3t0U8DBtYUTKy9MnAXgT+tYrHZdh7NvHL0xzX6G
GX2qF+s+gnZKUaSaxEvko5xezd/brCsXPTa/hxfFSfZzVUqcEasfx9qSTgLd6g2QvMfz/+FmKsxo
sW+1SrDvbP7+phrjhCj8FFZznaJe0VcQZnyrnUYCTKV+oxbub13pDJeIXHXem/73M2s51qwMyM0k
XMquYKhqcaFY717uIxAr+kX4KyUNM/Z6CXbbBXQHj7Tx4ZKLTLMWN39daL696UtseWGqRiC4o8It
c4CIh+YDrXqckLOZyNYDjBLg8cKoCJY2VLfFEipq20FVZdibJ7oY8zoKTuSNP5A6U8uuUrTC/S4R
HFhOPkMRNTNiTls/CPPOHKEdI2Vz+ECuxsp0UiUCEx6qFap7m1w6hGOOSh6yaaGWJky4JOSsnzqh
yBi+PcAAWBarrF6btXj0eFUZbheBJWS4jrbJ1q6i0R9Ch6D7wDtP2lxTJh8sVUr5s99NB3+ejREC
J7QEJOcUSmk1tzQBgoa1l4vQ0RyUiX1MlNCdQK9N0LDr4nF0sFTIf+f5tugIKR1ElTDX5RwANa0h
FSODw8uMeZoN0+B3PmxIR35zy6BzSEwi+pk65H/d8IpaRE1RaaSsRymygF800/IFbZQRquAvGCvf
V9VuF6lie6mIsHONrkHbv182sSFahp+ve8b9u5B+ex3POm2HN+x7aDCvSQDZ6/KU+avoM2qHbnMA
8YAEiGLF66xFIf7AcRZvbM4a/4youBpJ/vw0226Dm3T4f7ZMc9wDLK9q/BhKkX+qERKWyuw1uB23
hldGevcVK7N4tdmjuLHA5t7+nutM/yeIY6Aus5/QfHeWeDQZ7jJwLy3JhsGdisw2g4h3Phi3gDwh
yksY7X/Qwr7Hc3x+yRfuOpclpm7svSu1n2eo0luJpxDj+N40d7b7cMSiDdx2ppb0oYLGMXpqwNNn
1jzQBoUvZzdbPgqp42iga2exQiw9QpsmU91zfoIAQAOK3ub0ZkBgf8KGamZBN5Rno8E1HRYoPwJR
m0VsufASTe/4fSiQfRYgsu9NYilR0msK6TagROm1JURu+mnfDCHUEio/7Tl1YGjhg9WmB8Lk7idp
m8uYLcce8odcRePcC5ci1C1LaE3xxJCTqVaECH8ilAa0YflkoIWBkNtbu1EAC0xB2NFub+tcR5cC
+/9S7XNHoWsPIMEXJHc5xIIJEtzy9dKzohHCn/Pd1eskdRadIah8xWpwbMg41efkrJr+DFczNp6b
j+ZCoCUE5+3kSPSRTuIVIpRrU1QjFEMj13MNhIiacLxZVbqmjIWe7u2LJZSDn16G44Pi1EnWBy2B
aSYr3dRAXenLV4hFPJGTBdxSBq4TD2p7mkKnN5gW+10t7b/qma/pjBTHeS96NgLTMlveZNi93x+G
Lk8ph8C51Bcew2OC2dbqsioLt5b1o1fc6RhJYOTakJ5gZqSXXSOpl1vVSVjzm3eJxX1FqjM3lwQ4
qVNMyAHuydL4IZewj3ryaS+gI/3Ka+8xSrp1ZGJMgpdNM//LZoJxyOYM8wZZPd77T5U4kEkfDQM0
2bpjd57voKbVorGnZVdhgFsyO8638WonxXVtwLv2BoJbbcKaWmjA5jIZjCzMTGtBLSSS6KYNuczw
tNG+notCSRhRhCw/vj0zTWUTAKV7BkSqDM/aKKEkCxBxS0yG2G27sqlDhrry/8tjbetgYnGC71u1
eqTbJuwA1HVnmiwYMO1fPoRWPp7xxXl88svD2DV1bezp5CpiVIMhEDEYTiQtu9bBy2KERflNkv5A
XhzpvnCmPWUPbiJkecYoW5Hdocaw1vq26eNPPUqRiEk3+G+EtQFXCqhURAeYFDQL7kjf5DUw92MQ
wlqdJJSvc1GLyNk+g4Jo7qdO9XDZVJUw6vFkDmi2IvzNiFa7AdTxk8fDtgyNHBjB6ZvLjZVVGzIg
TMqnNWAsUh2lRayfiAsrIzxLF3Ag+ZuZghJL3/12nQtSL5R2MHFM1wBx1kNcWiaNZ7hDcg8F/D3x
gnguByseQnFIJ3Q8QCqG5WiEPbStIj9VCATjti7jTs0Cv0gCd+PJ7HZ38Mr4J203zo1MYd68ZADJ
lnOBrxz1tBnphE4azQtiAysU4kGO8VjonyIGsflps4GFabzyAqphnIvQwpOWUOuy+x6SxNkmmtBb
Y/s0ZEkbp26aXG+UxKaZJ6QyeEkIeOfugzApkn0LPtfFAOunjanIVj73kDpvv80kNyP2IcArhxzA
HNsfo5Fbg+S0t1rXT/A5Jyyu0MLAZx8AhN07N88CjcTNrcCpIVC0SJGs0HBdq8V+4VOT6mS3RnPK
sWW3/k9CATB9i1UTlqEW7xjD60uzpc8JxJm6u83pLAFyreCWAQM6J3C5LiXnqNj6PZT375ve3FME
EOzM98HfRdxRCgZNtIAnBRQcKkVHHBOlVnVG5i/LL2bh+YgIsOQeTmQhJf1W3+B3nOaDHaUEw81p
7NenklKRUo0iweALIwLnW7Vz0VTfS6v+3bmGYT7w0BWsbu3i2G2v1pjSA805qvnd122Fe0IATZSq
0+YYu/cihInl8XNTyoOX80ZWpw04M+PlskQlXJhcJdfi+8L7+b28tCuNKi1zJQEv9gz5btEM5SKC
KoKhWFn7viKZ9BerRGxuDOt1kYlhPrRF6JUU3X4wbFCGYqczm92Udc0yNeQf2ZdQmkVKXhAh29mV
bLsZcOTc+scrSseUVZ8DK9auWT4/CuCD52867slSfT7Zx97mwxXmX+LMsraQBo9whSw+9/Fcwmgo
hAkqLTUGdrNIl167YxNtAxAQwlS3mLkfQzdMlyc2OtRS9QlhiYaFPP2+ppbm4eM58F2BZckqyn40
niMgfDdcCo7wsA4hnWzVHD2O8vtHG1Plznsd3+mRa4LkOJVeeKVGRKV+Y6nE03zI5qHEYyf+wwah
hWn+F87BGwVJ9b9jyEw+CpqIWq+nVym2Gc6LjsA6R4IxeTdEQRjantSsfVKhnNWAb0ajbnFohFnj
2/ZIOjsGRzG4t7qaRCj117uRbBdnHH8VyNSMSgqpP3mlmYbDGAL8kDCXZ2WGVyCv2pCOtwLFiRcF
eSnDgtB7a5tWwFshUBkBnELeY9gT00BhH2PJWm/y8cblnUm3SwAksFYELZVr5wB9TY5OrXFfD/6k
cTK6BUbNdBs5aVGBoRrBpAvTyusUwTv1bCtuiK957Hmux2H6LjlFwtCAeGY1N/7GMFZwPlzKY5Tq
XPP+jqUIT8KXstYK24eB38orxuul/nUxpv/VZ1D4C9N2muBV0Pi+WR/RMEbzu7JwkOwGP6K5bDbW
XoJZ8LbbrrzBgu45RM7OA66tnLkmHeuqBbBuj6jDFnwkpU1i0Q1PfI77ENq+adkCXxhGJbrtC1kP
ma++UGL8PdY9WdeLRMCYyAxp6S8g44di9U3AeaBuAednTE3xBJy8nHKgZ9Inb80CGJ3JLfMbu1/F
e14YNZIfsz05UDH1v/DvJGTAnWzthlL/c64RsPsK9EGmJ4OA+TQ71poAvOLsZaM/+nOZXU5KahyN
b/CXgVn9NDdIBAXZL04SlZrf80MwF91By1rPb3nThOoMLiOzJmXX5jC1NQ2cVMAuENRynFsoXtc/
yHjiZ/ncV33LHJnk/81qL1er7bfZrmZsbiH9AlnzvWf7AH9z3wT8CUkhsH5w9YHUD0ho98wHZhe5
WOWTgUDHRPExxOoR19NFTgq7k8GX94mrAa0e/oL+I2ddbLFR+Kigeamq5p1rZUTHylYFNbi7tvDF
d3N2UE1cRqiFGKWRMRRDmUy0FJoMDUytFLT2dGrhLWET5uCWcz+fmurw+HLml91Bd8i2pa3EnX1D
McqyEs1JLMs28YQ5WRztUubR8vSl1z+45/KBSfizt1rEfaL72AtaQnltglbEXSNec2il7FHvWg2A
lR30Sf/765oHuTA9Zmp6UU6t0+brmKn5R9QloY6imOlPfa+UH0uSWqid69wJH+PEpDTPMKWZvp+l
f/gy3eYYRdVuDkpsM61YRQK2tCuE4ZV8OAKmL+5oFsEluOd0C1r/uIJBXg5+e72D8Pf18CCZvQLb
FbL1oUlRJqkPYAk/bjRBiJajOxhTeziKHmYTqTjlOhLJDqmCNXy/BLJ4umtwM2iWM2K3M8sr+ZsZ
zZpbBOgevkbxeWKIHG3XbCll0cEKABqs1T6Z5eNmcon+J8WDDZL5rAYB3HjM3qjeIN7UQDT8mgxl
JVkpROFuN7c6xbGmGqc/Kk2DcnaXKEEEZzrUXYWoDnyDisFboZ9cBvZAAXHg8x4GuddRljKGalbK
2p55fKJnu5u26ZyVk8Srwjdcpwx9d/MFAabWOHLbdD/ib0Dj2IJVb51xEQ8V+u4UbZURvw0KmIyx
VnO76xZyBIfp2WP2aIT1/mU8GBM0dD7dMMona1wtd0+cKqtUEYwgsBQPTCPUjt8IO2yKNVqj/z57
+YKZ0/noOXbHQpJggdH+Rb+rlAaHNL68PFhqMsXcJcl6Tv4jadgV7NRKnrWqdGWoVVYiaS/JyhuQ
6Z0AA6rm5hF1cPLy3QByn9z2UoVeBAWsBCNnRQT4gv1U6XBVPT5d8zIPAW5S5nna7ZGz8UVv1pTb
vaqwS+G9JcZNzDrm23YEOqvbHGWKnkVcOGTsX/bReWfzBvy7HlOPbQ0UusvFNe8OFQkvKn2fMtWw
pJW/+3w6rIX+r/TE+szSdg+L6TpBvJ0Qkm4L96drqb4NgvtCw+ViwZXw3Oz+lNhz3fd3yojDMMCv
9mnK4/gE+7cK7VCMioypZnsrQNHYGBQFDhfq2/xVRayNlURJTIbLfygPzSr5P8CwB8s0k3VmmnHK
Kxrg25F5e/icLpU27fav6Y6hwyzoU37KI3Ns8scrl1ljMHnqfjhqhLmZNzZA9DLDkUmePV8xMkGP
lDAC0RuNaf08Fz4tHnHqub0ovOl4PgGVu/z2G4OvHPVbmY1LpRFBSENnGCeDx2yLxzXhqSWJayGx
FQ98aQJhLepd7kDMMFeWbqFHzt4vx5ymHVgfLqdA3LhLJeJXTkQi8g0dRpAm6TrUKH7qh7DRY4Eu
51d/79Ftj2biBVqVabLEvXy/HRq9Qum/hPa398ZSL8ss8D/GNZFYIiG72g0uWxmXfyU00mwpUATP
UD1JWb9umqYFQlzP/SZRI/f+0S07sMnPWddRSryLbRva4FqMMEOR2UdzoSGgSZf48Za8ZCyU/6MJ
lir8ZpNhpLOHCm3X83u3DI1wgFTL4oYlvyB8fHGhsikhpR04zHJWdNzam+NLr0kIL3RBvDvXm5bL
GouyYYiBekx7upV9piDSPPEBVFkIgjyCDJ9mY061Tm9DTnBUjbLBmBBFj88sj4Twr4V1cv7j3FJI
Zf2wYk5oCZ0bFHMU9x40Oe4/dQlWuGk+x3VX6j3zOo+wJriroYQrrDMlHDFqZmkASkMXe5lGqCBA
NZwfSu20pOtSD+Pyo3+j2hN+RQSsu0B+IS6kHSB3QGO6yERqFUlDO2OjpDccMXhpfs1ZcEJ18FmM
GLgg+Rw6l920ollQZ4NED1YTCDE4KJVC/0nTF5uT5PLN6f6onX/zgBRjOnPUCx5FS7XbLRHawg+P
z/r7x8e429jI/N8q6SIhhdSky5nm5JL7PZ98xDH3+LvSHwan2H2++EQ0+JfEyBLRLg7QQedOrOiD
65GtOQ9KZ9R6Q2mFl2/vk6XiqPoPTtDCFulFXpmAvY9jW9fj30Db4Q5N8Sf7vx3y/dHAxwy18j15
IYB6eU4AesJEAynenz43tPBTtZvdqH1p+QscpyrDbmEF2qg1Uf2E5JVLs734t2EoVM6fe2RGpA9F
sOdf6T9H7vn1OAb0Mzi5cNvlgDsG1woSYO3ZRJWsF0o4HTKemAwa+OZmVdCKEqGgsW8OmhXMIBqI
N0DgrdaVedLh5XI+bR5fIOlt8eBoj8+Xn+96MIO6mc02RAZf5udDiLIYL2S6+1gnq8wZwuRsAyTl
hTXSCsunK5dvOOE/Iu6QLV/incrrppb2cYuD6rogVxCFLH2D6t4tDYtLIn4Zq3/mSmtgspHTww2y
IKKkYE54YGrQLD26xHj374vCP4jV0jj6k1iyZn2Wia4SGqtz1+Y846Z8DDx7WfAbLT3AlAN78zVP
Na/gnfV6YlPHwM3OqhE94KRxhvuwC5OkImNyQKc9c2uyxeR9yH4MRn6oH8w4U+jl8gEA1lc+dlXv
8W/0Sg0wMi9+ym+DGIzsIxSWaYRgMvdRBK/kz7kAKiZ+WY+NNCxPfSsyhUE73lUkMAKiAmLQsRSw
q/yxT/6aN78W8QI29fomkblieLZbAMY5ShDcOnmIeBujpae0FLNwqw1IptBXRgrFACFnWaWnOXGq
IYQK3lCo1R5msZZseNoElr/jjJ7cIJdlcxr8oiNYJzCshuhtApJ6AXp1jj9ZMJ22+pkT+EnVeg5S
neyLyjsP3Jm6ddFYc9RRu9+yBDUTObVpTWrzHNZZOT0qXkahjpRVX3GQwdorKPIPBrHzPW08t+XR
j2RqI5fiJ45nDF7duqu+qkKK+TsGsLQGuhtkKvPQNxhpYyjeWmeYVC2ge/+kLCdhzmqdYf63KvnU
KBXZmV+/w1fdBmntn+AVDCQp5ZyvlCh8Koi4lzD3Z4NfXQJoQPrkEFBBCRr19yytrjkxEZxeJN7w
9KJSdks+avkoRUEsLcC9SvPqB6TxXAda3tgj0E6MRiaLWfXPU56QYtylZlO9F0hiUHAs8U1UUAol
C1E0LGtYrfbVzyDIeU6x2PeK1pl54y2c5RBUIfgxkcjEOzebGXp1CJdyzFUa0/azLAaHn1VnZhv7
wy+tnCXq7YGLxG+7A5BR07l3pDN4jPWhJJa5zvbhi/DY0bvG9RaYpofoxtm+aaFVlC6Ui5yQl2C3
s8WOyHiHbmCtdPta3w4OftSqAVlFhPK5vn0eTHZADa7fVnw9oj+ivW0vTeJWEcxm6N8yhvl8t0B9
afmBpxp8fY6q6jJApHKCwo164LuOrWTVUPZCx3HaeoRwASsJzSljeV+It2e9404vyekEQmuAQJvG
OeVZj9SgQLc9zxeoLjAjwJfGFxOBe0yTn75Ejk9nteFVd4MtnJ0g2KaxV4C4FZaI8puAHJ7W+YHl
SQRr9JQ10WqlU2PzxxsAA4UwY6zAPefrIct5FBYVwsof6K2c3+jPevNydsZS+DTOmZoA7mogy4Mc
0RqTf8sGH2s2voSThJv8qKRtM6wDD0t6V4/pBUVAX0W40dS2b81CjDQ3PeGxG1THUurGVC+FXAmP
1tUFiGncjxTZ53wQ2oToa8zOlAmUsGDQkZmcZ4pGkjTw05SqL1MbEaLBzmRG2hMxfBOVeNkv1QZf
KmrgxA5N1mvMbWxBXNSlutDIWYED/wK2B3vd25l4ZyMhiBEv8bvAdi3EZ9NUOcqFywphkHCZUXjr
PbMaQJIehmHQ9gysKtCoLu54iD2Vm9ltgn2kYvGvwT6pAyLm68GP8QlSGcRDgx4ulJj94asbHUXL
VusukwT5vY0aH9XbV6G+kgcMMINisdJ2qijD29mGU+XGzEs2VZl/O3JbouZvqVBs8dJon2vC6DZv
DwtxrzauaoZUmG0buu+5btTsKgjZdPXreihp+hEbn/V4xomJCMahCOvs/TGPZZ4aJphn9Zyi0P8m
tGL7Hm3MjhwmnxIJCuHkM+WjraBcVi54Zsvwm0JgI7krJWIJMwu9LorYl0pY4Pm5tN/C29Yj2Nyn
yBR1Cn+WiUWdKn1KCeBmTcpKIMRqj1plvTDXZXp2pVjRWNNvcHWIBos/pEOomkHk86NalDwz8qJw
UudNxfpDOHkb3YzzcbWzvUtuY+2wYt9oplMZYkVxMF29K/PYNneNg4JPze4u5bmB2AqXTJyPOxaD
AdsWNE++6zORMYf+hnikFXXpNU6LLaTq1ePgMhcOQTWwpr2Y75HctDnrJPQIZy9yVdKOC/mSeKPo
5Mv3vCoCmXpSEMXNmf1sWtN78pTr68YsE0wO9woh90DkmpC8CLTxhB0ZPcOY8tCAyeeo8FPhy5wp
HTUGKpIw6N0NEDs7m1w85ZK+YHstdateTXl+z63FZ3quMOMaU+BHqvkXSo34EiBVEoeHT9lFEkPX
U0F4S7H4yhzCcQmqm6BwZ74mlA0S3URd+yA3BchuaqS+GvMBKXuVuOokG/uLlq0o9Xy1o+/fZZ/I
e5+W5GlQx27Xt8iRumqe8rq8ooaxseuBw+Ld3d0zOZxH8zg1gVEChouDS/gNIZoNbxL7LXWIsw+h
KEg98q1ZepkVIZ9zHOqz7dazZsy5r7ejvbd/q5fatXUdGXjHLUJoHOwvV+PMxiOXA+4YJTTcyzfk
pSGyGW7qyB52ONto1UQP/9FzCJ+qiKXJfD/fXekL1X6DGkfrDWYd5mJVVYwYWji2/p32jZB+nB8f
Y0oj6GY9dt/gK70RUkA7ocGiozxlLfN8xJi9mwRzDpmbxfHXYjW4mV3mwu8yfEhyxyuWz2+NwAXC
EWkzar1JG5MxScLRwAXAFigf4gv095xKGb9Cx/eOa1cUNfH39OnrvO9Tuadmj02hhwIJAYc4WoKY
p0ZFtZ3r9pJTBvrNhbLDsp2iEWqXVvLTNhdX3wa8sJ4/s89sz0E8LKD6/EkoteKpyiruOUEOm0kQ
0Ds3jj1GzQSEDq56HfGxvIDaTJHXk0bPnjpWJBnHxuAgRMY7GAdchE1xtUWZK+6aA3s10L7y4H5C
XOaWE7E2wNzAbmSpXnz15A0ddQ6B3OCEgwpj5Mdzy7XRMd/xynp6+irbFXUASE2r8AGShV2MRAkW
jQ1WOvvcZyensLsRv0ubocGao5VmR7kEqOg7cPXCvB/RiCsLJda+XxhiaWzguwpzWfI9J/wL3PrC
G1hNICEwFLrkdpJny8lLb9Su9q/Fa5na9fu88cOsN7K8vK1vY1/tZtoT/Z9LPd9BBqcjGvrAi9HX
Um5QpNZlIAYPa6KMLbjgbKotlrZhxajmhZj4ux0zQFLDP9ffrGgpQFqQVNeFmJoWxjlUPr46U9nK
tsXMMzDbh9xOAV0IAO3ALG9sBdTuR4HgBeQM2Hh3U3rTaDkjg5Q1VX72Ry27SK+BvMJmwqWVyL3o
1NtwYVI5ml/tXkd1DzHRkQ300UmFcJ3PbIg+iegrh8qLnDYb1Bp9Mea1+rSklpBcRCTMm42PPF55
2TzpSzI3rQpGOd2ROakt3+NL7gkYjDGNGkRdtTvbhCzMugyZ8D+O9tkqSbtznpZW9/EImsqWlKCL
3I8DSlJGc9tdyVqE0Y7/JhJYjU6Fd4P9zlmrf0ENbigDfHNJsHxayA8ZvIBs0KJDvzwUadxOe7/z
RWfHT3slRJiREXa/qkO/SW/BoumFgulnvol1VuHG4Pltl81NtRrT2Z1Tx/GCZDkiixvmhNXgRruB
Op8TRQGgS3RvoZs9yJbyQwdL3zSs/Qn5cnQK5JUarBNYirJ7xUQurKqJzKcLEMkMw42KhXyXcQTj
w3Wm5PQZ7p8N3CDAcLvcVGezsH92/PvNjQLvZkeOFGhGEdg4LOHEzgi/xIVrS9PU7ZYiboTGL9L4
HiFko7UKKMhyzQIDwMnYuxeMLkIvEmfGSoM3XAvFwEKzvm5x5AHR/6FaL3OGkjiNlAiv/8/aFFEw
KfVklOgKgPYbPT0eE5QMu+7rq0TUXsvskg8A9240QMWxyHVuuYvaVKGkknx4qC0MI5bYNhnncNmw
w1IBxs1qL3LrRho7Fvk5mt/mI1zTJyxx52ndZ/ZHEjBcPcvevRE5TrKwFnJRZGCIGJq/Q7q4EpHp
f2GBMv+OCMfWRWVaSEcmT7og6wR1AMXF2D6+I9TiPpwtVxE3HGrsBeS/PtEZH7OP4CjVWsMJHuGh
DpBs7eU07hky5kzRYi9sho9Lq2Z45FXX/pgl4UEgK705kShXDV0cgToOkMiyWbVS80J5fMyl+c/j
Mhfm9RKKOTvZ1BrZnS4o5U+JN2qEXgu9y5q2/3pQyzNi9bxMzIDJcvhv6WTfl1JFgsNBskSUYocR
/URW+FhwAroBdk7NsNvAYN0FCAkU6sLsNtxwp4ruBCqXYDrbSi8E3HRYEngeG9R6QkugO4rfycMY
57JE4vrgoYBhTugVN6JOln85J0wVcI4vh+X7CZkwK3Ms0kQYd0dA2VHc21Q9jJ5O147W5Dk1pgAQ
YWK2rCzGdBMgRllmdHaX8auqhN5Di7566NGkfOvWCQu7BPPp3dypjnyvtySDXQYNQd/Cewu5gS+F
KrH7xjhE+8J3o41KQ+59kEGJOE3b4fWMfFKeTPjZACttcbYIyppPs9R4qoJiotxc9k9vTHmqj4Qi
pk784Fi4pFJ0+iWnVLcxk5z5glgYMSczZyLA/NECw/sHLPuce6RKsQoCyqEVwP3MU9Z5yvPiv80j
dW8eW06An16djbgrLD20mYtmtCVNZsas/v4IAvR/AeccznF9rdg5EsMtVApUzfYfRX2yD5ctTh1p
SYrppzQ2i9c2ciRzIDydrNtnLu+ZD3rKH39/7KjI0Fu11itOmZiNiMa7aMGQEpNjYHTpuEhsQM6v
tj/bk7y9iBsHRDXB3a05/sWtSEC3E0oPdm57boAOYC1gMKfHw5L2j41/4/WKAeq4i1NryCmcU+0j
nkCQl2vBaNa/7Fdopbw/MtWUBC6At8bd2MHwAXvqixcsRjry3EIrtk1+fup5WkIsRN1cM90vaZo0
u2HvyPVRXkx4iMtlfhIOcaauZl+Z3h8tmxoS/7eL5j0Lj/AyMfYQLRIDpyxi00xdsbsUpGmCkNW2
CwTXMdq+qBqr9Tmw58Lp9KlxSFjspK7z5jZZgt4ePO1quUZ4WuHhQGnFnuOhWSMKFrlQTt3+oS9k
+9ewYUkpji8cawN6uCYO9h+8o5vE3r1Jt0iIhIZUsyEuA2UHvL+Mr2voGwnOB8wX9yezWTB/XdiX
DtBPFBPrOgNf4re2XxSDKKOC1rmqINvCm0YEDOh093IQrvNPAAG7wlK1nRcDoFPcFioIRBwEO5Yb
SM7or0OfeSv7IRyj+HKDqjWdEWdV8fxs7HObu9vdAqFLwYMnkJtYDRYmdsda9rHTSR2QeZw8xma2
t5jNGzQaohbrEGbgod3T7YX44kVTjSJLa0ZHXmcgGvQhsowlt/wRfeXVMl4yie/afgycg0v1IFaj
vv22tm7cbykeoPTibIOJktaegGc1KdFMp5pt+nxCO6VSCz6cwKfcHXrI+KO//ri+Ta7XeNTKQ83N
bDn/H4NAbmcA/9GgR7FlBb+3vFH6ScaRnKfMihR0ua09sG3s+3ihqWUZPEcbSHMVOV2u8qsImYI2
HPF2UNl0RDVzy7BSZm1hfwO38ga4tPc+RVVPNRdTmYQltFm+GKmnfjHgjVNMY+3JZ0ymEZbTY7Ms
F+cgRP0t9n0I9/ZqHiPUVkaFeV4xdAw8HhYobXjLfBU9JpUWsls+Cvz9Vq6elZKRr02Vy+1V/xEl
tgmd/tCuiMv5808UQo018/QullMfFIDZ3ANOEZrAvq4a7UCTNO1zoPoKxe2Mk/E962ybCjMZqWFX
83fDiR1pJx2u1hevyL2Zja0dyKtb4KCLdBBFOv4DYWznRg42KpZDSHtMoL6qtbTkfyp8P71sp1v2
PaNDOu4v0v6DgVjiuSsqWf6pCP2DMAfOXf2jrkoC87tU0AgZqc59VnKv8v8aVtNu/YLqoaQ4FE8a
AQwUfClWikuIp/VKPJgdcbcvgY+N/P1CGWEXnleaWWX5Pc5YTVPK8AQqBpNU0TSYZ47lxTPwbEdu
MZVaa8EhmQdEJAQ8gJneQ8HNM94qNwh7r5EinxAzwe9lIWvT5CidI+jonPz2jmQAu5Wms+1hC1I7
JhCUsj2rSE2GTNyfj+b+5d75spkTB6ftypiWAHRSExp5HZhzYpJHCpW8cSO+W+I1Is57XROT7EWf
8NtB74bchK11GwoI/v9Gr8c7B4HKXwSbAwizVO/KjeQIhQ6pvvg5PYOesQrfGkK+7PebkI6Zw7Ng
6MtHAmABsElS1qcteTvsb9ZMlDPeu6TVP8XjM+RXP18jVjgTQR+4ANzHcA5fhq/xmlNMyYD0xiD8
oUI5QkaXlNqU5yL9UDrSxH2vvSnfjjBh0rwUNgcPhMv3f0JxdxAB1kyGcrJ1PGAlCoSEVsRQ7qiD
nnq7oMSlNhnVrxki9PlRV4efau8l3tiCrwri8ROMeJcEUYrwtykHJhfHEDoO6ZKjPOwo2PaOoJYw
hITRs4KhgCenqzHqXoCdOWYzQCl8Y/z5bOROAc5AV/DRtavUOfl7hPgFsNcR5wVg+FCYP+GfYBJK
EYqg9qVEl2K/W8+wsP0IrdVrzOCLpXkuxUqnxD3Ug1/AZX9TSiCV+BnTT1woIYz8jPFlckUHfqCJ
/2puGHpU25aX9gAGtPZ1i22TZCO+xmZV5h6zif1Kwndt3XnN1qwEgaiQAPem75evzkYtU3tM47hB
NIvA5nUOCr0Upr2ZG9m9Ol0SA7XnYn4fuKu1tvmUOSN4agCAxerBnVXEF2/gTP6jvbGMIwgD05k9
U6oMBkWQeF2DnyPedBAApqsZdgn7TqLqj5SEVvd++x5i8MwEiXLI8FoGGCbabORJVASzUPKW+VO4
eFiqTxRmg8zArC5Z7LgxNtKyU0lnu19+Fc2uHDhvVGAbUj1A4s3sIKhesrpCg9GY7Tx7iqVUNiBj
RmVs+CtFMDN0wqV+gF6GJHv/KYZ07Xm0IGPAPkAJydWBTWVSGZw60jNjzu4iAVAIcMvore3Tc5mI
lZ6it+IjmyXxGscuPZQuVKjtWpVnUZI5nfjrOS5HRvMJ2YEyvStfQio6Qpn1Dh56QzID2fBodo9k
ecAZmGN2qYfjQ5iHopdIFcYNFrsNf6HJVVIf2Ns/afKky+mSmeTx50IsJs+gq/N4ymgLAwJv1srv
4H9Tkh4isnSnj9OUna7svae22aEc3UjUAEnT5X9ldkYS2zC/QEvJraEda3ay04gBBkPuL6/5e5ov
zmoMasPHw4CPHCTzjtNOeHRFh0t/zMMf4aCHzwIoJDEtApnv3mK5OA48VNQVQIhbeBulvFYPOdWV
wdftdn2sgFLLRzm9OoPUGRHRNzLLZcmC6BSeZhihRc43ZCi/KblvLEqyeWh+oqh/a5R/ExuGZPM/
HuC4kESGy8GCvDYdupKDOuNwsdd/p5i0tbWJikUTngzL1J6iS9vNVDDlJulqXAnWaFDB3diXbvAs
220sP4OnFKPiMB7ohBXEcZMMBn3CT2IPY9DzQWT1VUgNryzvibrCuYEuHXfuNDNbY/lWUNs+K97V
bq9mS7cDpRs4A85m9eq+H54Olv2HJ3gtsrE+K9qtR9SAOerxDxb1EmZj6e9+vs/RwwAXrTcZFUjt
LsFc7skBksh9OZTV6aoom/SRShAeAxNQzOcJ1dlXLB4mw+odSV7nD84XyTAxdNVxeTnJ74IolFHr
z+7PRLwR6pw6wbaWM03AZWZRtAr9B0fP/m6mPf0iecTzj9g0U7t4p1NIOG3Q9kKLqpbvXtDV2TQK
lsbytnStK0eIbv99aEOzCrFGwrsu9uXmASNyExIJcZHmqdafGNZfNl4ZBuu6hv0O6q2M5b4ipbsi
5wev+KJVFExOrPxrVfe2zPWFQTu7JEOSddNW05y6JZE8X18JzWA7BO2cKv18hBpOWNIdEKdc/T+Y
5YmjbkVP2htMpLeGUssRyXVqxq6EfzLIF+M/xKplOtt+x/JDPsWCLYXSjWd7vZqV2C1EZiB4H1mT
z7oUcdHfqJf70zomhRTByuC31OccDcvHlWmn18YNeyZ1Az5/XvegWRb4gpZxpRCS34kfUW5jjseu
dcKbrp5kekF2DZBoLXlJoDD92Chgyj1okUv8wG4s/gZuVJe/WMgqUcIO+V3eWNEinkLTF6M5YEgo
WuomU5lM1VNAGQj0EtTv7iUy1Muqr9+OrKBngIWserctrMqC+ekU3ja9YKL98ZY05ClMYpY3Do+X
oQGHcz6c52IclhnE0EkwXF/rhmkYbGdTP+tUUId6iuifVXSG2iGppcrAfjTOdARJwYCJtJMYdJRJ
Djo90QA1kSUMXQlBrqJP0RwuM+4BWWL0Hrx9v35CZR4H0YU5bpISmFYa6tvGFp7ir+Agaez0KBZF
yeHON4ZvunqyMWTPc4FgNf3VI2lbtACYGU8mJd5ZtC2Za8c3oN/QCZyqyAxq7epRoKoc+9UP56QD
OIP5y9XudOmfgOtrYQ+SdqqZ1r8N22xQdIP2ska49WgLXNTqDzE/a6T3GcM507YGh0PiMrpONDwX
Ae3JkETv5YZGXiIhVPsbBVjsiwGcpOimfU+OIF5tx6k89hIgsIugYGoLBMRfprY11Wbl4SIz7nPK
3prmjUyPMMLakCdQXolFeMZs82fRbXa6bW09dwJmA2nHKeawPB8k1omuWh2N109yXCVPiPblkg6y
LJP1Oh/nmrSlYXrJqAVt3TAhM9HNmPulbuDyJ0/vTQm+EEV0bodpvFxRcRyGKJ59tzQuQ8Z4Fmv/
OU4k3eT0KvZqyDI/5AY3SaWkVoapwB5pgweEIF2wuzeyiQLUOTS8LFNwuHz+WFQP452YX8EZ3Nyk
sK9W3dcVR+J/qJkaSvH+W/Li27+QqpqL30AysZbQdk0jsAmquR5mc5v/Jvx174YHVoeS5+ypFfJI
4XWxpkF4wkSj9Orq6izx0FIbhvGbV0I+l9fESDQA/BcNnBPfU4rlzjV+1iHWlBmBAJ2DiUA2gCHs
nKSUEQXaNt67ADbzmMQisKM45gYcm7v689Y4HC3DrERMFIZ9Nl9SZCbLO+RoOCBNam1qgDP/SRJJ
ES/pfXEVu+dOLwIpDf9Frke9mG0qBdHZkf8zT57Q6vgZ7DRYK2KMeYxXn04MkXs/ReLQOPGw6a+s
8UVC942tK+jo6+RIQcdm7F3FWEquUWdfGA4T7SBEe6VVq9nHBjR5ozS6fKjtcHJahdrvzLsq1OuH
r/aRBd6ZzLo9yGFNDtldNP+na6bK2iVoMY5jaotOPuDwxERm5JBEt3Pqg32eJMSRkAVdeC9eqxEH
8ZAr0ztWoZBY904ghOSB5M6MsRIWLQPfXgK8lbyHHc2QIXh1/7RHy/VGgkGEkaAfGfFRXjkWnMCJ
YA3Z9Lw5aX0FqL0XzljawR3+I2vw5TCe2hCQz6Ew5Wm3OA5BCeb56tWM/ApCWPRqTZ+RIwbp0T7Y
CRvZNq9MLd1b+BqHjfgMjYz6TzVJKT3ugJoQoRxfp/Zi/ntVnkWwIQSvpigw9+9I8ZGxbNz0J/K3
7wICHZr2/HJ3C1uPuE/O0mLM/agACqcWxiyKuWPpHeX+rUwPOMy/GWbjE847NeWK1ulIE8mgrY7w
/9xV/jidlqicmUnMMZfA0GCrbeUnQX0J/r+lVCwt7zsRRQ0qCyam4VHL5XNx8sVV3Au2LfEmYbh8
yE+7sMb37ES+x5UNZfehLLINDmAgFSWPrNI5QqhW1zl2b3YuHIjfFGA0u9pCV3BM1tundcBn+H6Q
i2dW5vA+l0oheeUay6e/r7H2OTTxR1Tu5h4xW+CnpTpZi5TSctIupr5FJ58FCayqGTgqKwUwfNfw
YAwtr6fWv9i+lLzrbkVuLI0YwiRNitCKZmulLd8A6UksN1q4v+vOudHxccen/u/4YZENnTv5cpcq
GheTNg3krgtxraRPUznFipUS1NBiXQ+o0S+I6/qiBvpskPJCYXOJ4pEcUDmeuCrH+6bCoGzhVXEP
7HouiLSixwb2Yrvt0p1vooxDU88KGMMf67KiJMy+jc+ynMQxkgr6qyI6oa6xpAOztcNdnqE+VvV9
b1QNkam3+LYYAj9G99w+SSWaXPP1Z8uqlUXX8WUY4WG+VlKGZIEMtuiZoZ3C0xTBKwBaZhHv1Ve9
BxmDuf5kMCY5Bbfi6jfyjVAG70JsJrFnLpBWJPb4Gj9I/vMT1YZS9T8AsB7uL4kiRH3M1Sx6zZ8B
k89iwfugdSrIiOUEQDbt05GnP6MPRsdjQntAwgfXPO3p1LtLB4wX1UFfH05+5z+tlHSV7xSZxH3b
7jVmFYG7FERAB+ilSltU1LXo39CduLa9pY8koXGUoVHsnKlLUWO1yB4S5Dpdhn668U063oveYbUj
gbYjpTWC5GeNcLwyIi3Uwqqb5ynz1nV67ReSs3CysNE2hZO4EBc4D7DQTtjSIeWxJIDeboufe6lG
uajCpKEe3f+BeGm9VlEEHss4yY7wA4vaVZXxVfUrvbxBpmZZhDl/fz4pWjFlo2E5x9Mrpy03M7Zi
BNvq5b/DIGh5uADnfe8n5DssWVLNvnTPgKozr0W49inUmWP0SDVZXxaQP+iouSGqLFCgJGfLAgml
X4jWjn5acCXZZjDxkgxi7ySj/K5HvIkpiF1JBrphzwxKxLKSJwMKP9nwV2jvThW9m/BUApatNggH
W+f4He3EX8dSh5uHvvtV8U07aUjlFm/sbAfZJQSdnZo2kL0Sv78aRlj6Zy0oj16XBJuyZ53X3ArG
e2mKkREdI+LA3qhmKr6OB30AprttLHOaM5ZWlE/blkHQ16RFZOYE96ONxVJkn4G0/vJQ/b12tkX2
SfGvX+ynSbaC2Cq3n05/zUx/t8sPTqsu5BmFAcQQzPsF0qcu2c6PDYWGOedyzb0NeZjP6Yecp+hW
CQXQrdNCIBD/6jthn2syGt0oEg4d1cS+sKBmYRLryPpVIQu8sQvLXiNdwUBOAGCYyJvlbLSN7EvR
xs0LoVsXThyHmWBR8QIaESyJSeQ2UL8LM/zLT15r8QTbyaHtOsW2ds9BpPdGDznfPGfnYWs3LYQN
YY5W8BRH3FwBIihp73W3BwnCOZ+3fkjJBO0ewAig6sqJsAztIm8mjodOXDQXKY11IzlGL3z0iWE0
Npcp1/+t9kqu/Ep+gt98V+6fb6/2CJBGufmVG25NkjuCRzLrtJoBcDvAMzbh6wNaon7Oq9060ZF/
ZSh/MTPW6tANQAKrmLUzO3vZBBJT50iilTuQjMg1e56lCsFvxexUMERbU5hgDgk1/J6a9Kpac6xu
aYSvyDPrfWXPlBH/X/7+hId+Hq14KfjipqAwbD+R6la/QzaXnGHJhtfClQBOLD2lr703V6itFM8C
3xC7Y5OXapbZnn6RJD30QmxbxbIE+mAcRrfZJF4SqGjq1IO2CuY0Jb5c5owBwRth6/j621kIG3OM
egmc4FG3UcMdC469pVWs9VlWk7cZf9DTxNcC6iUlEsouH5Bb7PD+llhhsEEODMzcaNKOJzigKcf2
B1QvrpZixC8c5mlyIFHyPaWiQ0SMqL7OSUgUTfmdW3nku+8xflz44LKzKHMwQxByU8z0aSJAXlLn
N5Hf7Ndc5nmVXzr5sQ7ry+EzllWkTcHjqHkf7WZuTPwgKTcRFWFeguHepZOd6oiwEXLNyAt/RiLP
KE6gOiogEpmVba3FHCJJka1byZH4o9XZGhM6K1UiiZj3JihPGTmmih4SSwapjgIKyhpLRk+XM1WF
sp3wPKxhFKzrIUHyjxWAYx4/hpFGcba81W5NX2o2EF5lepBP0Cn3Lm7WDVhPkynJOVl5CKGw9zHl
+HpTuXqmD/mXD8N9rvpP1gD2aV64Vpb+KA+/OaVpd6eci7jyJrQVAinSCHBqU7ojN2VXSo6HUCPR
EdW0z5vOzR1rL4GAUfEQzmMbhamMLXVPpJ1zqdcM+XYEsCoHBT6MLalo05mfNjMXJgE0NgVcLcDi
hn+kPvy90WyyORsczwcnfud6xs4Z40BrhCMCSvDQLxPL/fGtfSFkCrtgvvOZKq4+eWY8IggLv5VR
kWcfTO4vmRw5TZ5a1K3mqfPsIN1RUxq+BDDbneADGkaaia9/110Xv5h3wzy3IYxfljX2gGDp8NX7
gVPCpSVW854jlfGpwKQ6AmQcz3YZOhUZLWS8vlT8Ih0ZTCpeTF1qfGqn2Uxx65hYxcl78Eitqoz3
QAaVwCx7YipcpUZjmfQ6moIb3Mzt+nffJyNEgIHzPfzYyK6WP7j2oTTFrX2Qa80gMkuSSwe/+AT5
qTcA2E2MY75Uppc/IIpTZMSn6AKMIjKLE2d3za8Tt/8ggVkWpJP0FOletHof26TTvUr8iPNMVaac
nv0JvC9OjqBHYXD0QwGo+tREO422dxRzWsul2PhEr/PCuu+2+YIE+eE61Uo4HsHsWr+poSL5EVgh
5SYhwNgLoC9K2pvwVLFzvGftobmcZSZcolx0a1VUGl9tbW43MPtoIRMKrecv9jbGwxsOUzQmN9ux
3fs4lmmvs7wC23jiXhq6aQ7+bvoJJcyuxaWita1hMfMqTRT7pFvLzZsl7oCNfOSUTJviErXSfsn/
9aPVbugGxKz7HW/ki8lCJcGfGC4GI9caUPPVLLinlPyv8DeX6lOEZtUOe+GamM0XdjvGzIc5/8+Z
oRXPQ5x+6Il2EuA3ntqQAcW//BHFYwrq2z2HEcodNUZP+36h4RGG6jVoHSnN2pvQ6/uTqq/dHFGA
A2wSTRWEs5vq94Bw9Gly/2EOc+gP1qpAmaUsjude5toKqQg4E9iGlBQ4rC0JnumxvAOBJX5xojme
PDp6x2uNsM6maTn6pb4a8efYnCVracr1VgK65d1Aq9NN1I+PSADYO4BWVfchUm02RdcPAoNw1Tjh
/WneoMLo8Be2fOZSi8fBomiMIeKPYuTPCHDbHLFVNl+Z3AeOBsR7+Y6iRQS4GmH8LuHmX0t31iBT
EgEJVQm9/Xl1oPIQhN181h35MF3cglRP66RVoS5Lscmk88L765VzUuuCisjeLgqllxOpF4ugkfIH
yOD0/MPKLsG6l7ezvpBop8VixVis2YJ6DKJcYNTxJw4hkUdJiNlPKf1R2Ikr/4YkFpr8GkAvOxkP
M9FnqxJ9jk8G4sqRqy/2YB+V8IxKs5ffFIyEb5hzT7FRNBL1sADade6cpfiEg2G97mXnDnjXAd31
4WX/wAbJCvFrHxuOg/qldvA8+6PpVPmNrnF8pxuRZo0Lh7F5BTaRWkS34QpfiRlTTeqmNX3if1uw
hP4ZZvPd65eRe8zkSHvJTejlZ1cXyiDVtwxCq4AsHuQJni7PuZnA0L7WRMRvhLz96n6yMBkeQbit
KtpJ+Xix66Ts7KUB/GtwS3AU5Of4ocO44Y0IuAGuP2l7Gl3h0yTunfbptSutqfHHYHmni5i2qEwj
fe4o21DNCiPJE2BQDK56XoPtlECwJHiSiNS17JHOR/BERQfpe7SWzvRI4pGaqh2TjP/WNKs7qYCO
l2PYfSz35RVeym5CqwIKoXW3w6gUHmhn6tXANAaBRATGEQM00JvIA82DpQEH5bAkxib21iGWRH8f
sKhtHQODRh/bhji8rpepP0XkBsTEsLwYu1WgVSlbAgSVJzGeCQflCwCVCFVlqk/B66iJyloBYMWt
be2Du4CFXUWyHdL/oq7X/oMX1GQ3dztHPLxUnLDNAIKOi68WeHTGFIVpKI0aw5s7OC7c0TXJY6zv
++JlOeGrvralUaHNhAYq3cLZ7jC4MSsn29EMLIsdm7IBtA+9fiki2ebuFvIECu6hkgpUDbxPa5ux
aiqROdPrUB8Npg2tG6Md46gCYIcI/6Q3xULptKFJaOoUDtSNFdJQmgAI0javGQ6cesDfcHJ9ceuC
lj61QUPp5/0d1uEF7CQgK+WtrQ9dTLer4a4HqrBSB5kAKI7Rjciv88trabe/UgbyJoeI6f6ML8UR
iL/B+MVeI9RGMlxydF1Ydb1yEEGsSxNTTkIz/SNnSejv0zHvhxnnjNFFiO8f5I9xYrET2/Lzbm4d
vMPx57BUXwl+wrcpLRGLTVOjms3JZGvsJTts8JCMDYyWKsiDL6Sm4GzxOjKK0HzTMu9oOUP6qHyi
aOeMrSY5dH+sHdcdBJTf37XbmKfybwn2f68sueKh3xCtU8fGKfYGLMxY1ouIop2tW1MmYWrMYIaD
Sa1F4dlANeD65DAXC3x4AfhBatyZunJL70S4gw1LLPI41AZyJwdveGoMAnFJfkERxO5h3UB+jz9O
f0GUyJ9dtWIDM6K1YJhO3NmhDJ98b8P1PkBCDVSvBsvlL2KZHdEkji3Y1VsnfXz/7UKLVco3SkPe
4pGOvNhxIk3Ymqm+pXPulKUpv3mJDjj48VYR2ASBT05IJiScwJmCgH/GpIrj5Pf+9uFCO7upb/hs
oX8lpTeblQD0i/dBPeoV+SgSFmLkbx58EkiZLFsroa+MH0qm+S2XOYn3Iq57m3n09pI4of1EPLo4
NUmgVkfvqw1Nr0lE3SQziCpu5ybKOJSKRvAkMvNJ4cQgkQ83izjKgwoWnDmmS9w+5ITy5Cqgk3fs
+xakUovSeG+P/v4aTwtsDjQ0SJQ9ikGo2u59N+Y/h5DcVMwZm+3HLzT4N1hz1WdKhDLTLJop9OjW
PlB6daqh48H3NxnIlKhlIGV1B8w+x5pR6hrnV9xL1jusV4890HsCw3y8pACb5CTokaM05qI9k1xN
tC5L1C984NizJMp3t5gHcw197QopVEt1MvmOA7aYoKHTGliRmDLCICdf1FYiGAoWlpbZ/Eft1/sy
3vp+CBKOXenMPlrySen2z8+vPX/OUjRTOimKa5KtzhtTmDwOdO6ivGUEiC0DlEkcHLXG91Fl32lP
wdfG43KzNATA5kjMIdBS1SlkGxhcbuRlF++JMEFu3g8kmF83j3o5OOjv/60ygis1gR1gxKqQDTJn
0I6t2p3dYy+AkWeCUhGiwywyHrlDUO/rW1q5WPfZOp/MSO5tRTrNjNTBFxYOdEAh1C+nsVS5DweW
WoaNEu5lT6cw0Vva+vXwWaIznbEndo7/0ORXqPEY6vy5m4BDL4jjzuyKds3yaMQWl4BWa6bgRDIY
b72DyzJCpvjO41ohvrft37/CzkqCKnYfnsBumcdQ40GmbcTIr1/VMhC14GRwURmHBeOt/sbjl03U
LIhOJI2vURUNmQozQyR+cH6/GTmkM9SUuannKRfB4VKAjJxYs7SilZjZiQof6D7glEW8DCRq/8CR
a/gtA90qELxJsUIiyqqalbPK+LkJudPyzMbrkR7nTvnGuK3au3O/ePe4jh6SO9KPT84cQZR311Kw
hKlE+S52QdLC+TFVIlyT2xCg7U6xJNT1H6FXCOF6SUoUym1h6kxYp6gH1qpegSjNodLiZarvq8OX
LLlnCvgTcPsPR724vz7oMWxmCCFDZDerwT30+PIuZB5jWVc5oyEOhP53Yp4m8EEcyE7l64QHoGe9
bIE4Kbf53fozrHShKZmNm5c2pUI0yPTiQRCx5TyIBaxQOFpWEUEF4//2d9iead4399EHyCtG1PAM
wGokGQrlxfm2obmxiVnUHsJTjtyA5La8QL9TFsypZPE7EG/xkgtaqj4IIupJYB4r1KispoSeYz+s
7gROhpuR2b/GTJb6lzJ45PMfHEMow6MG7FW/RdCdVl/fHD2Ly8vMhtx0TfCfzBP8GApgwHkNdUC1
hZvt1Wjpn1pKMVvJDYdOOLmZffBv0Qz1/QQFfgYZrSAOYS4L+KMSbHbKFxOMZf06sHywfDYwDAfl
MRBNhsvQ5Gl19sxVBubFgiSpOwtVUYFeNqMUG6Y/m1hFznpzq16rrXJcFScFhZnJRZSRie5MZKlD
+yh47qJwJQHnC1a7sXufojbwTeyxybrADxXOjyOjOvW5XRVbTfOSsscmuz69aiqwrd6Iyfaip3KM
jgQdf/318czVJBEbqIGVTFNF6qD19xIzxDQfo2jSOZq4Loa5j3KDtCm3hZb5P/CpjITWmgvvabTe
V6M8rqsG56Cpum1Q/ohiduvPpa5RVAdP33eWe+pUvCQq7tCH22tM+zUsrKWpicsec8Tkhu1ixtwY
thCCq2g/TZXuIM+kOhjWXBWLhmcaAHPP4DwYVLih8IyphfyXTm/mGlPpoSbWMQ//hlTktCG5643r
z08HMZsrV4I7aAHqvPQmljeTOZ9a2WzrmyId2IrG6xN5g3C4stBcPnX13gpBFJBCRS1oiPNTt1AW
KIBaRNgHTraY8btJSUQavXkRpFZ1IG6hugiOSaIy0/MY1RlQmHIjrcLtFd6JmMPZajD5CmHutLLy
g822Rs9U7x66yBChbhNytArBpg7Meblful6V4Xagom9ydQX/QXpFjkf9cQk6X7XlhSql29bQ1105
sWGjnto4Uj/McxWUVExCSHraN4F+WFtug+qK+NNspdQcYrW7ovgUGo8tQYtLK5I2Hke2ym9at+wS
z5Jyxwm3YxeRaHoNfv/ZXH977j94eTgQ9tOUA7h89OUxvvaevxGuxc/IFHHH4yXRWyksJPcnZLc3
IH/zahiLcyY36vQqZ497jMbUjMgw6ItaaCb/Zlvm6FMCsOoppOlygsKax+8BH3FHme4HRvoKQVgB
CbRkUTpPXb7EAMLcy/uwC6ivH+easZT5YtJE+Pz67ngZBqtzPisMsxfUVAexj2qHUjbioJDExHj/
HWmihqxDgN6c81ZPr8mC3OPZ6e4Ws3opQEF7PPMqKXsdJ2h6Gb22qKQPlthx6t4HWkpuV3iooNi2
KmKWArDrSloEwksnyxFilhQxscmKJ+xyEHc/b8t7ugZrJyCkzY99ZBL3exGY6EisXVvAgi7C1wSz
W8uTkbo9cRo0q6r5JhJ0eZq5w5ASBOSmmrSdIhzFeSTkm1XBjKbK8PcM+EuAMmn4yIkGsGzcpJqP
TQJp8XJJoB/e5FqMCbVfIpvWAKXsisO1chpOSPLJQdNy2QrMLCU3yPeH5HD6r3lC3AJFnR36oyoK
Oksy5UA/Fo/FGNKTkhPcUVwNYy11zKKB5S9SZcvLT1/5+kDGCEdx2aNVA6JoLMgqFvL8VE0V61dY
nCOD37Ub6UPyVsdv3juop+j6fAUEKAaFap1Iv4+G9VOUQBET5qkn8TKk0I2ZcTwWWeVvC53JHG2D
X3B5U9wSjwUEnv+ZRUhEReY9rgTai/nQMGr5U6D0SdsbrNIlgUgX1N6s4y4P/DMeBmwU+JtxAfnQ
k/uHRgesP1oO6I+tYNfy3/ETdCn7GzqRMaLJbUZHYghjy5oWh27NzuVVzNmO7X9vcOAuLDi5QrMB
qY1458bMFaVPMvZ24dO2vzX3MO3RaTCmE+g0Up9vvSqcme3YqZg65OjSNNVykKiUjhkqXP4sd/T8
UiVsvX0Wy/TjmhtxNV+gqEfdV0iYrvHjFLTHE9kWzmVrlWBhILhBTsi2bzaec8JiYw1dUqSFO5/Y
yPtPy/YtreRvA1bcXtAhp7S3Z7zoHf/EP8R667+g7R+IgTywsuITMlkWU/xib/8bxqmBrn4V1s8L
gYwsaTDyPHs+ZeXQ3TSDMi5coadYDSEc/5OEK1HEVN9UZfUzKESD5IBJnYWfmbFIoCvJERX77gqz
H+Euh0s4nreF0eUiY6pGAS9u7g0vfc/Oqvq2hVkqJjaIjWof+jcCXAK0RgGyrFd0MDpucKn6EyYs
maD3vZ4AxoMVV/DbWSq0Gt6foiPT59cH2Y4hswR1zTYVeQulIj0MZzmZuLBgwuSTJj1EkaOn5fwD
qwkSj9HefSIOBfTcjLWMm2ZxBpUgSgFXzg/domV/mhdl8BqKeEd9bQdLj9nOiuAa5Y7r+9XMdd49
yQtTaWKMCATLNWltnDiXBeRbW5FVOPqvbVBu+FY5nazzWttblXJewIV8UCaXd8g7NSxLCc5uWbk+
5rTed5wZCFTSz2O5XZAxJMlQf73AIghbWHZlUWjQGMVK2qO0XHDx1H5+n8zK2StN//323Mk/htV3
9ctm1RvMXbx8jjtxpFfm8iyVRvm9RszRLNfcbOlG4AaAHu4zdHCLzWYx2ulbgpV6PqE5lQU+6YsG
FZPJkhV6wz/LIqgv5DdOGabJEK1RaCb0AdFV19jYei4Fo+87XHcp2k5Eb31mQOUAtZkpVoLQSEHs
FomMBFe0mK7+0sDkOfNCIzg9SHwOcURalxgql5PeSmwbgmPEVz169a3HY3ewKoNv8NabVBohrr8e
ObzqvIRv9j6mCRvObMtpTz8pezi9omVl0eVUl2VApLzrhjATyB01MZk3UIfFpKftl3K9mOiZqKpW
S/KjXJHnfvkU0xx9dWtHRDeWO2NvC3JaN9iTao+qdOWP0nH0ODiza8hxFmQ+IRHCGObdJ0LGyVP/
yw2r0EoBTkInDL/YC5Jr65wxtEHXOQ3D5GHnN7kEjT9Qm327fr7sMU2lxW/JOuT+JAgRLhLIJE1n
oHabAqVBfc4xH24ygO29SJ5HQH4Y/xvobc/9w8D3Oj8TLyLUOTRNprUk43AXGxRrTox2KcBwswyT
VVSEQG9oHAm6pJjAKolK9b81wmHp0v9ewvZBvvLkFMydywL6ee7sqz4XZ/RAUQbiEa/X4azhG1Sk
MPhKNRv4u5hHFCWp5SNFYx3ON66lIqQhJdcd6uuNT+HBg2wxhG4QQjSzY8IcY0NE8OVhP3TXu3fY
8IQvUxZ+fmZlXqXsafZ1OXJsJlOHDsqTdwsHyYZYjXm229zjRTUu76ml7QiOBsP9lgV0pVWSj3fv
c4L1omDDjbJYt/w5vMApvya81StJ+mALUTqvPOB9OyaANJAQlUO5j6vNplAAkwz5EkNKFieHnP/s
LEVu7G3Io8w4yo4fhxBFXOPANEf/tuTVMfTphIboPQvPgc6sccaYmCXd/3+39jayFvO1l8qWYKvc
qvwATMIJIXO58Ok9LGn+ehlwHdC/AgMgdjeHzSGhRGt9h7ib0Vxab0dofM8Tfk9xGny9zEcRVM5B
abhcFfPUa/jT2BJEMdU3UOYMZ7XmIHI9BF1aY5r0g7h14prlVT+apNiw6CBtDX6bLN23PqcrlbmM
XdEPTpioIMKSxeaDD9Y1KESqI+HuS6jRrBW8B0kzwaibFS0egc2X5Apuypk2rMTVwz/+MKRBTVF3
vS4DxvG9YX9MRj130amXnUvLglzrdNZDN50fDY/IlSUwy6iQCxoJAqGKQBLgGpZRNIID+Ofcddpb
mGQ2OYncj2SE3BmVXaHDF1d9MsOoSOdicSajFTjdzZACXIyqZzJydvDvbXTZmOsPlxqt7FCiba0b
cpREuySFLCor2A6FklwsfgVbwRIL3u3WBM6QFpcCzUQdY2omgVbSAnb0YkPVUR6CrFLmvVuYSRWo
RJ2BqFWtF1zs7Nx4L7+t4KlEmUVTwcKD/SM8t+StSVDon0Z/YMHwUzYVKbIGsq92US1vGG0wgdxc
RQDszIjUmsNSLms7IO/tpFphtLJgIN/Fqs++Ax0JkVNfoVnrc0P6Oh36XPfCZx8VZrPO8Qb0EfoD
ByE9AgWtiy7HmEpY1oB/u/mH0le+ZBm1FEP7QE0hlSgIHvsmaYpEwWqtguxZ5THepF0wjcb7AgIL
K0mEgs12th1HkZZj5rtn/DoltbeZ4CJ+INKosW7ZubjzutqmrGbXYbcf4VtCDSC9voUuHplZ42g5
pt8LGtoIHrSfeXml9NJTJge7srW1DaCK6MkdGfPLmr5POROKkoTefeiOu4aOe2OTN+cIcKYgreas
j3dumuYh46ApsvKNaI7nhcTP0pxmTVmLbxsAG0WEgkrsRjbqN6o8FUKndhxLw7nCNGJYfpuaRDWO
sf18I+S0sotRk9fcOV1bzH+eEQhKfkWskRJsfF/yONOGMc8ahKGp35a7qsV9pDlSNhFNC1lUPnvJ
yru8dqWXvgLkO1gCxfsyP1oprZEuHKUTy7+zCsJ9OOhUt8pY+qxOkjfWhorIWxxEYas0wGYAL+OC
UQbWlpzqOfDa4BAk4Ie2l8fnGTn2rPaAI+k6/g8o3DoQnmbD+FQWR5C1ixIm3bhrd0XU5meqjCJW
Z2wJ9CG33vxsKxbCNt/XOjKCdN0feNTW3AauUrOlNNlWPwcARjHmRQRfhvkJHjbNRurWUX1y1az+
99bc8YEGUG/6aOMGuMeqDeN+9mwONnKibZneiHu/6qvvlYJaz1sVgm4ON7aoJWl+6xAl/GGuf/V/
6awIT6/U3hZ/ckAvxWebb/g1RaCzHkNw9/O2fzHz5ZNm/UkGzeYPT2tpSkoF4EGEXJc1sJsYGjKo
AywG9mt/cmM1IXiRhzt2f44ygXFB97S3sG3wc7ipuHAyxK35cM1KVkGTfJ7uiEO+8zFOTFovZmh0
bWB4GQayOvOiA85dhm76zGdADxiBevgloD/qmaEzWy9vzsOoP8iaqZDZHan9YTuHCy4Se2Rg32w/
w9EUrh5K6voDgkL4ev3sMIUTaIANnFvsS2VN3rYKKisd6suKbrdlKTfu73yw92vIuVw8LeosK5g7
EZdHq1R7OmGmqet2/EgDERSMQ1TV/uuUDO5kGJCscBqPvh/nzc6qZEUdGUYzPAJGJbTMPjI75XaC
z7IAJB1RBO3Twijq6YB65TTf8TlVukIQ1eewUzNwuW8hsEPS4vj7oF68xIvBEFkepR4X0kXRNUz1
NeviRobbXTtS15YV1a7SJ8kggNMrbOjSxky8BbxofzKdSuHaEK0gUiaPP9JB4pE/32K2qHGciyof
CI6F1DkDE1mwXmTB+IN6jdiCniGiYYGZlzJmnlireoZxbOIzy+yZAKqIJs9uKpAcPKMfGBl2C/dT
Jrx8g7qtxEKwbGxplalCJzANFn1ksOJi1uuqbnnGzhsAT1L/I8PDXzIUxO0nSe2WHUfiojuDlDiC
bb7WUXK77YhQ8IAWX4CwiJl6/wTP08EWjiTxwJedlQodeB4V9W5mOimyZ9BVMjfYPioSOd1lAwVr
DvD4vzPugJXt2DDxO4TZmA2JmTlJP1D9ZWYYpX0TMAt4vMUdiy5NwRjHPcRFMQQFexnLq83vn6xD
cRqoJ9zJ3pggW5AQuRLinc9ExjMUE/n3DM/W+rTeyzBstc+Ty8Nx/y5hH1C8gU8qaAvuimI91ng1
zYWoHSX58hr8BS63pZDRyb/CumRa3yLrA6f7zWsMgnjonCLEU23z9FbwZ9BkoCt3AtCroG1dYA/6
WwhcvwGsmhuNEi0D73nxlok1Xovchuty6DrdoOy+JDJleqDPorhUZTsKNeHYjzoAEVGZ1n1iC37X
KnIoIGno45w/jdthEFMkyKfsTwrRav+fKXf9Q+1vfAygqAyxfnGqCxwl7n4m/KWpM0wKVr//VuQD
aXDXVDK+/U3r0iBITs1voJH2X0zp8OCBK3scEPX5oXqoADocB3n2VB6ISFQzNxOuQ7lRj62++nEv
4mCA+PiYW7PtRrskPwvEKX5f0U3DsedeZTME3Rl/2uLaLlJFLCTQRcJ80dHVW9TXQZLgDsQm3EXe
LfKup7fWViduQNM3RFdC84VihrQhn7hMXp5AM95Eu70IudHv47km86FHFoY7IqUji61wCsB1FCn0
rTJ66xwBIZPAL3EJG2cv9dGOx0cMqOO1faeU/rHu0gUmL0BeqIgq22gLBk4MBDtrEum5CJ1IPdHc
0A/dWpB1GF36KmwnX1FoXSxtT1MolzRllfG6FtPBK3TE2Yzs1yutVuuk6YiTeQtOhA9ViTrMf/EU
1CpkpBfZYavcNwKi7e/ouR526E24UtyG6CKYfivVx7+juULrUqrD/8mSAjPBOQHKDUgIUoCyVdn9
jZxjvrRbajNnh1HPbNElbcslf3JD6VDLGTtBC4yVBg2Q6LiCTgf9n6uq3tpAKCg6Fx8nikgRmBl2
gklrNeZsApYa0n3anIm8+G32kktpScaGGPq8M5vHJ02W4lAaQC5xo/JogISsgMmYMt+hMkRm7Sg5
W3Njj81JcsLcwSqXBiFvofDxd03wBvrkbC8GPedwHIedRSQZp3DsFzV/yOofFCX7i6LQnU4UXp71
dAqbAmN2EnUqRygSfq8E2tdRtZQqESmZSFlCfbr5pP4aB+Oxb/nRg152OoEmRwNYajMiuHkMQ4cf
gWJdCJlbumH4nwCz5XSGWN/RgScCAAJDSOVMiRbyfzGBQ5dR5QwBXRckdlAcXpAe2VjdiDiUE6if
NKuFYOEkY9vn5hZYHtZ8ON/TqM+PA3kHXlRVZ3zTk+xEVRwg1HKeFlJ+zIrqX75+UIVQnJDChxLq
2WKkKs2M0VaPnGKJms1AD9w4dA1mKngwFH6g481EOldLQsmuU4GzmGgWejLqxtDB5vhxKbZZQEAo
Ome2We3QprOX0X540RLsm6padR21uGcHXiNukYSO7q/WvgHQI0WBZJeZX+vMyUgy56JA7a9Il8RO
IhC3S2SP0cqhB7AJiswFL/lATGPuMUCl5BKaxKOe/2FQMk1QnaGAinkVjZa6gi3Qu5SjHkjj9c0q
e1w7XHc4aKL7gjKtxKFoNp3pIt7h/7uaAtrIEmafDKOFynbXGpuWg0KvxOviWPCUQqmvOtTxvvIj
paCbGMnr01rpMkBA2AeQgbPq4fT1LuU/d2bl0E9UW2wXUyOUl3JokgqhPTIgQSeHp/dN5GxxtLce
S5Vu5mM9ZFiIv+cqcsV3QfKgWNdtDewKw0pqiQADkSlgMY4aKaOfspOhEZ63cw6W1OrGyH3EEw54
6WWL2h/s2HmXEgfbiaBncGupWmp/lOESvStkg8NJ81Zws8Xx2IglHhb5sg7FNqVOj10aPfXfrQ3A
mCOLEFQ+zusWKNppQFU/4AeiDrots0Pv4GicQolqTG90xXBkWti4dX+9JuEWr8Stly9elpCT7YWw
FSB23qpKCkVy9MoSW/x6bdjONaJnePvAqn3zWfy86RibHR9gnw1k4QK6kiiR3MEqNolVWq21Ekos
cQPY56B2S+5t+wU9uZWXqTfbD/F2Yi6qYb25fBoxGZzbtCEYGon9coDw3nP+duA9ITEU8roXTuBe
GAnqVbQmO3izzSHVGpYk5KbNZxW3ewqwSBTQ9ctiBsiBXPPycV19r6OrGw3qpOS8J7FlGndpjEO1
eyWmzCFCXIHIwmsF0W9Ny1fqCEdYp40LLeuLqE3sDjP+zeQyTBiWSOOkWTkPLrgLwLe/UuJA9LBy
Qk2XZAyGkC2o1PoLcHMhsIdhAr7EOhv8srjcm2NJWhbCtTX6xdIGPR9j0R447umQIOrWqLNV9UZU
Td01wa0alwY/M7swWxFMezJs4ng3ARSAovvckwJfRAwENWxr+qfP0RHpYiOK/REIGWhASD8nBIJJ
Y8wdUp3SEPu8mJ/l1T7po7utEsf7QGaN8cJrBUpv3/NM+IgUWET9+WJeIf7NXxmYMPxE2+UdIVph
VtrjJDXYj9TShrrtywb/PsJyP/rFW90uh8KiONyryF0a7LwBf6fOtc6Ae+UUeX1yuzHevbNYpY1y
0Fke5NgXCQlzZu/g+OPperHV6ql1+5WnhYOKjf1PTQW0QKYj8M2QWHEU1fWXmrvrkOhfgpV/hvd7
oBjzbuFI1MQ2r+lZ5RMSu7yEaenDKuLTH6xgmlKjChusmIGWb9A9+mLZ2UcC+CWxzRFj1UcVY/Gp
HR7eMmNQYVIgaW7bpXIK61w+YbT1L8v2KX0eZmxPBg6qiYuYxh2adnhRIguQ5BXC4/BtBs8AmTME
Zw9JZgqdi4gIJb3pdD6QqY+n271fYjEY+2NBPYu2Zpe4ZN2TcMDTJh6nRheLsX2Xy78nsYrsTpKo
lex5LzN7ZmEsCM3YcZ9y0u3xKhQ2iqvMtLFCKHti6noMvF2DGfVCjjFjD7O3EvJNRwx/cyowoHfo
qY75WxNe33KOCuobdG77dHa5hQ+Kmzavy/um8PO4LVJyd72/Q/Pwem/VxO/tSa9RMmNOu/KRMQXS
bOi+gKLK/TzMA7uevZT2/v7WwKcYymtEqnDx3OsSDds1nIUqvzVEnLRzBl6Mhh/uYfzVPCP86zDR
04HpapbA+6U+hap6FKInx8O63GaELVlbxTPZy8Yld9oSmhfclC5CwDe0tGgsy6wXNHsSXS2Rn0Jh
V90No5hV0ukZ/bIYd6MZTDEuNpL/W+Y6X88XnWgmQocpGwP7NY/cO9kgL0/q7GwYSOEHAkJZ1fZd
4QIm59rhjvV0uiTiJEhUom/Bm7e5tHTTZxdwd0out1c1V11GMGJskgf7k1e+L9OAN9ZmmH0IeM/k
yGsgvczP7v1teHriiF2mfOGl9s48rABV8+tK/SdGqSbv8HhGiF6GFOFn8yMxm2NPO90YhzCLT70j
8H5q7V1W10Ytk/IjRuYFlNWqwBlA2gE339MSf9OsCpKJd//FfkfE6C+QHTfULcBeSXAl/KHE+f6j
0cv/D4lANmbrBHIxx/E/hWzu+hL/zFl2M86Tqhh2+HM4ZWW8j21Qv4oqV+JeqhHzEZfqJkQYZC0w
d/XqSLfvMw9cBA9imkVqx/tVWwuBouIHzyCqtOgNo2NIQwiciz0MF+EmkTlEBXXs7kCL0bWLdHRo
hJfwX54qjM3N4VNgoFqZGpdEElVn12KM2XK1dGSWat7tKawONuKxVLd2aVqYxgBM2gvqiPO7jQEL
+KGRQukkTmh3tCxHyP7/fW4JegnphKPnIyRsvSqgQPO8eiO3WvQnF59hTT8t+kGRf7hrNVamQs7B
FObvzs2Vd9c1iVrg/+KtKmQZw2STR/oFzq4bjl63qGPJvuosX0j7EveiFk++Nqd1Q+Bwd+/lsrAC
PsPdQNfK12KLtU6acLynUrpcFYvTFN75guVNdcRjlUDRFL/hBVMmGVWDPG0cG4MwuyqRriWhuA3P
ezTylTSTtIlf9Fo6zz7Sl1xnCygi+oEYJfWacOQqdvG2rJFlQKZKODm3no7yRbie3M+njT6cvcsf
8EosFkJVi3fMlYamFDJ9j1B9DA/8LjP6Kr+eSOVRLAV+WEBK7pq9xByzx0FqIPvT0uRwtQQxy1bD
r9XWKTY8RSRrR+PE6Qg3Y1EzO1LQMHohW285/sLeBYX+mKorBsMZpNrP6xNmog5Q7W0SJBwMH5GF
1n+ZwBg/wl8m4+kxAaAP4dZjAygJ4vKIT5jmQSQVQdv+wRkta/8MS2t4VHytW4heqxsYcwKt3kid
FhhEPqkiL/YWa6RbFX7GKVS/8mmO5+ZDzAz7a9pzBV1qmTdrBTGr2omkFIxQ9FRs0+WConHagAOW
k8B3d05ToYI90VnSsWmUl9YzcySVi4ByhQS/V9zsQZ+LQLmiJ85E0aYhd71AJ+cGMI0nxOZy0E5i
GG7FvB6y6X5fNIdrcZ6MR1wxVX9g9NzQ6d007o31ogWM+w8Btonm//VCUJ1dPpUlzYQcC9uOkjwH
J4q2iLfQJsbLBV1JD0iglte1pyLyo9SZYj1pAgaFd6X/ukQ5uNyf5LO+leqIQfRKmWQuafaBAD9V
umua5j7ukL5QAn5oH0IMaVSVGRlJtUqkJZAd5ED0tIFj0V6estvFEesaFJAMUF9QNB4hrVQtLID9
sbXn3L/+Vse2J0rifiIe3v5eXKZ+G40Ea+6l0FeGb8RkDKgnl1asH+dg5HvDZjsDCeChQCISJOnV
8GRloRvBMc7b9CvtX4SVs/dkZuaY9a8IaeD/nw0Tew0Zp9ZTmIZM42n8KnSonT4cse7np4beWKAp
aTWjwUz7G20/2emyiKog9K7ioqsUKE9sEEx38TI9ocKxgw7g8pTWGAd15nyD2rcOW35J+bR+CvqE
8TOLI7mAGN8aR9EZ+enC3CIoJqft5emuwn0j0MQOOMqpFRcX4zW4+T+5CFcRc2mgKeJyVGpcyaI8
bU/mia2F6c03AY4HJPJVaXHNEK+zugErasutqoyghTZEBHFVSzDLdTWNaIC9+dL6vuOsCRpXQrZR
hss5FB+bzzpgkuPj5CMC9/ZI/m53csXFvhb8GWP5EYqy6e26Lq/xajEFprJWAU77gxBC9fx1HaI1
7yqgrPGNULCu+YqQAvU+QMPocmi/NFEq/bo9tITq71KqNiYPxVfhA+NEwsJMjVFgBMJ4PdUFC3iM
dhnxfpUqwobgg6oAclA2W42ozRkhy3koIJY81AXn3HfVaJSxW1fOqE+PWQqIzzokd3M6hCAxF2Tl
ywcbJoICF1qlrBYFk/Zq+XJLYVM9i9T0sc0ougk5dQBqB2o2o7yc+sFp0vuOg9OuomwrBCBwU3gD
iQ++iVaYBbllGlaAt+6WDIrxW/qRwGV4Qfc14XlT7leBEkMlb2vF5zTkVjnxArVFeIb/+j7U+q4d
VSdlcqwwwJ+cuOKUUX9B+g4m2O/3TZjO0eY9Sru2ZSZ+YkK87voQ8PnlmP+d7AGgdSj2pTt8IgXt
I4Bk6m2ZGNWnq1h+vo9GljOGR4Nj/+yHgtEzpJr3FSEz0yMV1ieXKBMPDi4W25eYBF1laE2htVS2
OpXjXtc4iLLN1WTneOPJtMPmqZllxhnGCxvWK4qDDTmQi07ZHjV7xQUIbRPdOwxRUXUpTeH57YTq
gjO/eqD76ru7lxyjKSMmsQhyJLTQrdQmLeqHC6ojG7XjQNKCLwZjB2rj17jg0PGWkM/2Nb7UIX5/
ryoG3JfYpAYYhKNAWq37sgQ1vvLvadRkOf4F2mq/9B8Fk7zXORBxEVrj9vC6/yDGGD0RP2A1VwkL
qKAulKGTRY0dpq6uWSW3apSp06SKoEVVrP5z/g4zxJZ9bBCzSf/rTqa+iGTivkFY8rhweFKYsrTf
l2KZu5igkaQxbtrnXWmkfpP3mcWRlEEj9uXluRqG5sxpnWUt0OkmV79kaoGovl+/u7IQ+rOuHvdz
8zXiyodSAlGS70DNGo2RYDJnvyZwtj1wNXjZdFCYUFNGRNMaawmWMT+Kkr8xZoKJiNBbHV9M98XW
bFOE5KIfEv183MiJQUFEt9UiklUJZ0Zrg5mLUyk0edCSra/hY0O4RebfeIebkmQtMbsmKk9QqIF+
+CT+asuTszNPedKOQRPMAc7+V8n/4Np+cynuIDweThN0B+rv9xYGSN+vKtivANxDVxHorfaVZaTr
vPUdmuDYC6BaFvby92NUTSCvx2Y5DQomJ4unhrnPz9hcGz7gxep7ezG8WUMI5WFsnppfoFI5TSDx
he/ktABx3X6nGT2te/w6XDfeaOZbPxMlO37vp0IkOaZPnsTdas44nQ8UINA+Tb2eiMFCPd4aZcCt
89QBo9WxfPp5v2cliBav0Wc9ZCNjQqprCNg9ACMkiF1R0+0pa70fYSQBhbpsgpsT8CjOWlIArtcD
I6QrauMKnbCEhvMyWT73VwoeT76GYN6B9Xoo8+R2oNtjUd0CVzywsaQenVd1O21Lt/7lbRuHczK9
uhtE50jbnZKPOIWkm6nv9QRXfKfUCJgNmbuXBvCTDDvAfLMOZHOADANXO/w5gHMO0gy9UD8+3+9m
uPhXt/lXwxiQ6ZxjFdc3HhJHHcWZGlvmpxL4ko+bpcLmLkmtSpXNNl7WlPLPDL4R3G0wtjtWTLGt
eErq+i9pR5q5CvKeubkkuo/x/FCqQw/DBALaXpDP//B7ygKVk4GLcLYGBVGf5iMnH2Kg0uD3VKEq
DuWzKZeinXvFEep6OnH/EMmoKZD8U9sWwmiGaKE1EfIMiXxGSlnecGjhJWkXJsaUA4v7scFeG/II
E4P8kk4nF/uwa3t3TiyMKu909rc/KQUY0NAdL3E8+2WlKF3RNgGF8DurtvZ4vJCa2prUPOT8WuV9
E4Hq3UMJtyhmetKcalDPAkUznBv742XwWk3RqlasDZYW7sFsmKHVXwGGr3uQ54Gw0A6KiyOhMBIY
hR4PXO2+7eOsBoPAem0QY/ujN3uI0BRg/pa48k3OI5BKavzeRI7YyhEd8c1JoUnnV+UH4pJYIJMc
FHrwuFYfY02HPbBOQZoFi+Wyp9M/LSoEm06GhR4PK91zL0P5KlvOjDHtpOGye4jb4lqOC5ME+u7F
e7Z5DLB6MmTxZ6if+JnmJzqsOQv/6JuIgl284p0IXV0AOXsRLnaSUGXbbNgNLy0YF4+DrqWi6QNF
G7DNKx8gLLNeBzhy5RlATrnWZmxacHSIOueCgWGKqpewtcnt8s0I2ml7oYtNPyteHJ7BQmnR4az3
Eg/m3CGpmT5d4++ISN+adts8HonaakbhKmXIoJrtdFip8VUEvM0AJi0sAHDgyWzYOWQKppbOtc7N
srO0swVgl9g9Ko4jVOe3eOp5WC6Y70hTRhUIrGsUwkxRqRnV5Crqgm2wNL3jarmgcGUjsOJqLv2g
pA96H+cwGyBs8SAgP8wfxmaYrQhh57vDLucQH7bB3hA51etC21uJ0BPaUpMWg2lOkUGsD0BTfZlT
Hf7Wh99YeZlm5TexJNdDNAqGFrBDxPiDaAnSabH0r3fKiHQ0nWdy02TRaTmr43rSnYg4cQ7kpU21
m3bzQ1qJP/Vs4ebEf7Qpd+xYn2hmX5qsujgTmIQGfxFMSOeugm7uQTwtKk453LzoUQzkjJ9Qfj8d
Jlmk0Y1OdZKsxti1EySVenmON9lifNNnVXoSSfqqnM/ZEyRAlLBm0jTh6C1sU37w64ST3KUAw5rd
I1Em/Ef5o+p8f2aZcKzFWrYppQgQjvEPxYRcB2rgRbvvMuyveHVvUOXQMJ5dP4OxTG98JqfpaU20
ETKJrxInycU88CJIvolMtqwLVev6643546nDAbMOQq5ARSR0Kf0/TkZuZQ4PUp3De1lKj7+lc6yD
Z9eEGguytR6fYflU/htrn4/GAw86633ZVKyzRzyabwi9jHgIXsLBIRLnHss/LW8SC3WQzcDQb7MK
vTbDGX0JKFHsdeylr9MhUNnHF6u4DTkk7bmdm7iYWgB5zhBfdV71wGrlAJLIW6JxqxKpe0vR1a9U
pCOXarhWNlINvKR4tL2lL3b1flnkRZ6duGnMOhIayZeV+MSu3Fe9fSBn2Kl9qNTd72URihyAwPDg
j5dvl7kAc5V14E2BlKRk6j0D4eNDtxesz7Lx6gy4Q2D6H0GNGdmZB108LkCqKvtiLoyBSCVRdicy
xh6XpvvljntKMRUEL2Fx/IU7L3noNzswHToESeHnCpOY5Rmp8WMGI3A75JL3BF7iR3qiT7ocmJxL
sn3EhdovFU8fJzT46zjBC4EerAb45qLVInGvYd1HagNR3IOa6BL9J0tkBXiWlbFkty7iHTxFV7QL
B/DBwI584lim9OfhiB/AXm1eLEpPsiWWgpVElOTrKpj4MgmAN6LtmHLAJk540i//0hWMn6dQcszT
oWvP+QDj+umiaQ3m+YWyfqVzklx/AMVN2z1fCZ+y7/zSaTdkBUxRyh/yRCS/lu4PaxEVLd+jIw+i
srgrCC/ebcKQBKRErtr5DnDTvECuWhETmApjbZm8+hIalh9wf9/HddrnqoseBgFPJApzYH8tqwgU
+dnqkHPe6kjvmYv8nqM+gDaV9NqqUpjdXaCkE0LXs9gD/4YCXhhrhei2RVq71fmqYinco+ynijxh
wE0k4+1X6VWVS+KUl9wCUmaQaeQE4JLz0TOIueKaovxXaOpRPizafuRPrebyLEwikFAUwOZPR3Fp
LyuazclG6Kraj4FcuPwc1GG98BBn1m/8uq3LTGBjEHcJ+FpC4spwdhx20NOfvGnYaOyAGr968Cq8
LyO1BeIk57CZQ0ovTK2CkWyAxQ5yW3cbe/sD59rWJHtV4ESiZRD9Yzh3E0WLabdQG7JgQx5Uanhj
8jyxTorzpnF0yvb+RNEUlRaYh8qytJ3kSlSn9rMmOn7UpT3P7xMuUQzmZJTppAPK5cBo9dsDfKrL
kVgV1vTCS+DZiIvQvMtMprRBUvYERnS0xmpgtswVyNBIAXIH28BUalKA8Oj3xV3wYsjqLs6xHifm
SEuf7wZjn7jyN09t27iEt7V+hT1YPviP/MD0RIWVJF74QyXNm6bUGzmmfKaS+lMLtBEqBZ/Kf1Sl
66LFVupMr4LVQvL6hgXIahXKqZkrAnWSoEufAwS1LBqyeS+3mXaDwNALFA1AFc8nakAwE1TnA6Wu
G91d+oFLmMQPC+3OayRH2x4qgby46Wttu5SfKM6uq99AiSzRSYd14hD3KwRHudjGvv98XIV5yji0
4f36M27iTIWRyXGdOtIA4VPpEMLoyUlk4++cwHo5uSDp1n7EXc7chuubjLxc4T8Q5srpyklCSyjj
h5SUgVQ/USd8sEfNDK7oXCZTIDVD4aouYxDOn70ud6KU6ZaCeIiq7BGGoLhdz1hQPiUC0VgtXbJO
d2up5eQ1GprzCc69rCsH0c+fxphggcuwh5v4QrrM5tsEAx0VtWxpRgB6t+7dqmkCc3IGC8/r5UgG
5p1Ap83JoawMc0ftNDvvVxffjTnonO2yqurxDMbKakD4YqcI18y7CRDu5xYoxwjMG/e0F/8FOftL
bYzXi7YarG4tpriBFfgftcy/HGSRyFeZ6bC5QlCgNP0/t1vqWAzfPmc00Gb3NZtvLuZEuV6wZHuz
7s1bt0y2NspHFSlWHhETewQo57Uq1Q/cNcY88fzAtLU9vYTTxlx6LIIfbRhk8O/YILl3hzbvQlD3
WWPXcx7HuUS4wOWCG6yywtF53uud4oIVOCvHL4b5r0JKOr7u35J61MRcnYyNyDUdSJDMo8osIpyR
galr46qChWlD1xiXv8BiawGjVKBpbKR8IzlTFcLWT/rZsISwAqZJVCEenS3EpI+xn/qBNNy2s3Gd
TzMVC8wfrBRnq7ojt/MMyLsCjCWRqs2u4A3nKhfgNZyCmPQfgO91hJqJOr0Q48yJtvGFGEIZhsQw
Jc7r/zBI5TF8In6q64Rt9schF1Znx8Dw+NZuKRI+je+eRLCoclaDHG2glUCmq7D2f51SQEaEUWIo
WbW5lCyjjQwOp4tZDXHUgQl5ylBjanmPulhNVlHK8Hmdw6Ww2DYYfOi5s0KLqhKvY49XCTIlZPbh
XZz73E9HAauOg+Rd5hbAGZY62CujzfPdBqCGeGCdaqcp14X29olgdWTdNE/8i5p5+iZUp91nEs6I
pRVtaDK33a6TjbiV+VsCCLy0wdo0zvNf9yRkaxgMVizGXAWM0J7G/KReoBb2nNT+uxRMu0kT0ndH
k0cyg4ZNcJpPTRhCxGVtLPd5ZbSqrT6JqwE8a6t6h7/oB9pEnXJkyG9Agyk7AmXALrdbqLi8gPAr
deQYgtKZZQB/Enfi3gJ5x3nzwEkWdbfq4zBKRSqvYnunduhjHydag1ZlzQbty1qDPjdn+8CDhk29
E00QKTyA4NdwsSQlGSJqLfUx6i5OrZk2QceWjYADO8oT+QlNF8kJOJYulVILWlE7bKQ+AJjC2p4R
Zo0A1tEWBLIzD2nG/Pl4qqtmhSDrNHndTnG9/nEJgg/B3RZ8N0oU/o3yXbIgUHNuAKDAUoioqDDF
lhJTLfy382vpdNhY+ILu1w954ZFXjFSlrKKwMB4EkjAELLe/SEDY1DJgxjoEZJSUO4iQswaBI6+4
7BiVKfFMQ0G+Ak22B0det3UW6JdmMvrfpoEi9zqrelQ++qba6KKjEIH4fnd7pS1y1gcNAITxmK45
BogjM5FjI7uKDEuo6dSB0ikxvPAzr/fhLCFCL3CKjdLYQCFnDkve/Df13IYlA4r/WpF0H71S7MRv
RaVrO8yVqxpXZPkxL5/cVtw3PfcxnTehOc0ELsCpM/wRl8rB8A/y9nVa2bdrIwFcGO0SZyRaJmf6
uEZ03xw4sk5w0haiO+ly/OJV05u3eCRkbi7POtlZ/DLb5Gq4U5TYka3fVjU9GiXN8/t2ECNfb/Ji
2DSJRdqVBglBw8T3+1I9pOxe+ORt2VnHksMt5RZq5xjoAG74+HH6G2VUiyksChm0tOPBCAGTafta
aD9ibofz4nVTWzCXB9E3ASb5uvXD/QfKCPaMHCOqS5/EtiAJgX9s64R1PUgJa/NJhWOy1qKUC9tH
+fEHnE89ohYO9sa9tiGoogNUO++W0pppNAgTrahnnVjbYIdencGw3CBMwGObySxNhKioL3zqYVib
D1Jr4GnHKmckqMKLxLEbi1UYLDO88aMt363+Q5GxU+szQbEsI5Tff1+HozgX41dAqyCkARrAoIby
5NdMbKQAxa9UN7FtSlB8LJM/ysgYy/MQvzEh4LhAtw97yJebvNCfAbkSbIEbcW3bLUce+Oa7mTzL
CCAVGMhwwvufqUNa2Uskay6xW9i8BbtehA3+0tlMFqsyTlD0xsMsnlNs1ZCTG6ArlbgHD5a8VKex
iIZNNG+wbXQ4UINY/BdGnH70E1QmaDXvTTDspCqxkQwZDcCwb0I3U9jSiUP5zXuWAD5HAnv+2sWt
7G0H9DGw6N/dpVU71fXSXE1s67gvRZX88y1TOaxM4uJ35d+/L/KTXrob6U8v27GzfP4PQHzc2GxO
ZieuWg5XVgpzVSbbY+jeugBkQQRAK/thxmYqESXjNuF8P6XgNl8DHMVjAEgej9ERI22NNAc6FzSh
JNdCEEcr31b+9WRmtfvRzzBoe+WFzyP11QmWTri6yhe4J4KM7psxRhtw0ZUlTPURF1nJhghYaSlB
fxATBzcbeMp2jz3z4lKDXsV54zDuzgDRflQSI4Xb4BzT2Qn5PBUWKLG20vld/yENn+lZ1JFrlQqQ
e/oJO3KOxJUPUNG3vBiVzsmrtA/IOSZCDPXZQY2nOKGxuXPcUY/UCAjT4YxTFnfCGKM1k0vrL+Uu
NAmzn0r42Nm2l3wiJIL8eBwSSXLmek/aPEs5fCq5D3/hFf8L0zK74q6WNswh8MA3ZeM8Uijlhwam
v5ps0EACkpieZrF8GDWP4cNLHCoBIMVZ5FtXUjJ2Ey7QLtO2HYHZ4WafttwohTviWQqCNFwyjlgM
X8F9k6vEezvqC98qPe7xd4zCcAsQDPfLDeRG1DojgZLpIB21LnTXjxplMZVFFUxNCBLRNNBK075b
1FPID2P1uFG29DAeELwq4hGSlW4p8R0RS3SR87Sn7kbKs+IAkRLaVnNIYzk5LC6Lj41jJ0qz0kvb
Mob18cF8XnLeaoqht28AOAg2kXfRHIj57i0P6e639LacCrJEal0c+2vgdfnDBQY627lGMaVxnKRH
QoPwJhQb4XYQbRU/MjdQ1CklPm+MCD0+sJSus9IIQ+WONBIgDjDDHTq2cYGn4Os5/ZjhRY2E/BXw
Pwpgo9ncfeBCan95jfFy+E3HFme90K4aFEZCjuxplsFwkeUWaULoPzDTtU6uxVkD6G5pAXeFarMr
CcDobg2Z8QY0SqMYclgB5a9qQKuY6u/7wtYKsORpc1u0I+SaqoRIcYrknCpmkh/WKPDtVMZ0//Vx
su3ZYGhBWZWs9EbQeASR2+BOECE4TKAJkXIdpO6JYBlpEL0AMguswGztaClcjiltm+u+Fwwmax3B
Vgmj5lHOMhhvcamShgJiXggXGY7X6zkn8pgmP3klT2nMn+YrVPsBLdNqjDBCgPhjK6psrH32Z09P
gKLWXqN+Ku+hnbOKtr3aPx38OzHN3LD6GXvPVNMrPxlXfVzQPhrqAGC9kjXCPya7P/SXJeVidOHa
pJEhKOKbKut3npU7mYl6e+TGhEFI2nfQurjzmBy+8UdMia7j5WNcEG42ioel9ts8x4IDGTdlyA7E
czB/fkRVWxH13t84UwnBiS1q9+zom4tlOQsqAB497yqifYBx07O2VgLA150XrTTEESkYlxdVSWfX
gPSFH0cqcOTsnt3wcHpeERxn1p+QMT1lwYa7Ry/G/EdMyLVB9TXz27lLdmVh5kFJdA8opYQdHQ0q
BLu35mjBwY5T565LJti1UA7eH2MFV1mwJzrkvv0No6C7VmPzcEFivyQ+jkkIJGW1o4UGVVdYYpTK
rM//5X8CffLTUwIjtYVysp5HPiafdkkJVwtZFqOf9TNSnd0/7wKmez3Jzg1I9LSNnm1cXNEn8xO/
pDaQkmaIHbU1I3GwCuHB7wz+z+/oh8lPHg+qdZfLMaTjj1UITjTY7KruDArRzt3ns8dKzZamNA8R
fctLK8t1bhOCcG7XJrAnQ+LGzE77nIr0QwsYKXWNaLDgo54+06e6lNF9eWC89n5592dcEDZBGVKn
70saLRsH3BJpMAWhuibGeCZi1Ym4taqwNVJmDvSSmUgz44UIxnDCjeXu81jmDP1Fgl92ibEGz21p
yGOyBGaiEZG08mjbKKwc8M3ct+CmIoHCI69WOR7Wf74hcG15YupDHfsEq1eOdDXpQeTaYDFGVQyE
R44tZH1Ia5H6AHRwYPMniZ/YqGb0Nn6j6els1lmIIwsQVlzk/q7hhSCC324elQUY8RjNeOBiYW4v
rF3dFpytdasOn8ppJlSQ3sXl/2x67aCHhUCc+s4q04e9UdRDDR6iBCfzXqbwb0gnu6KBv9h7R68M
BVjkSRLrWlGLnndi0ZITveWum8pfHPnJzJpW88EP9aPolJ0fGRMUDT+zQ5NXN2IHrSDnhnftGzMK
if8nZmfuyvxQmFdrV3VtuDop4gXBypBdAY71bShIKihUQrfgUR/F53ryBAxl4YJZ7hso6t4vMtL3
JsSpvYKLVK4WGr8byFCIoDsNBIBZmRGgCjnR//VkDuelUr/OdPKZQbBr18ElbhRIW70HgjBJ84F3
IlApFwz7gw2XztyvIVeMXDf4LjBBSWXi7mNJ5BAy8o5Cr83rGQbFDU1OpGq67AnT+a1zOJrqUgaL
mzurajr6noRrAll/2G13bhw/oVrnPKrq3jdYeoHNtjb4hL+HAP67zfKsX0y6TOwX1CDZW7max+8e
KRzTtuw7H4JU8EMBnQYvmCAjbeeU/Uo9cahdz97p0IeuPWS6QeVePm4clj21Cp9DmK0UcinDgZpy
Eh3HW0E15ASDURgiJtzfvoVozuCL/l9JtKiYN/UP15ZOsUzair5ja4jSYvLO3rbPJpt4RLt6TzAX
QNpBUoo4apytXZ5NvEpvqCdWG0K/uOubB8/E+f6vKnwfaJcklu7lLFFh+8cuiUtR9eZ+oZmZrG6J
c7rDqDQRMHJiM7r9nYEXMGbvH0CNI2Qye/McJbP798g/BBCKcA2bcTJsCKm/yRyMvBb/NKg+rRH0
u7jOjazu1mUic43qlodMpNNtCGgNs5O8UO2pqESBwDHiN0MdgXiwwBwst1y1FnCsjOviyOHKSqD4
Ri3RZdfpDHRHvAjuQPjSNFfmsoCedMDoYvsxDoOsNlbLLEeb/fnMi0RSrK1u2r1OFmcpfnW0wBVy
KUHmODTbv7sKQ6HUGrGNMKgC+AuRB7PjN62cRxJYcqNpvNi3WtzLE3FswtwVIqUAFHq04EEh3AZ5
YKFDht9B9KDJ3RYrVeS8ob6orZSA2O8/1WBqVIhhNc8DSwj2Wa33FqBsHHj9RI9qa9106yDAh310
9i8jFgiNTfCXzkfXFAPHTMMwHZRn8B1LYoSkS8Bz22PbBYeRECsvzJK6tlEw225muykZUPCFT2Un
XG/dNGWApSo7TyXXawLVj/n+J59WDE28q+HY6jbmEsetvgJw+iBbA64AAUdb6+pS25cvCfS+qXfJ
wfiC6WGQNqeLFB2bQT62K/PMCLgpq3qY/Rt6q7IJpkPT6F50zbJvWM3Z6tJ4vWNO9QXwDfqj1J27
/9iqKV46MIvbvQ21SCm+6RAL3SNw2xcl1rblorXzNQhPrX4bJc8ReoE1SCCW6XDy9CCsuTcHx/Q3
TFla9jN85YM7h5LdfjCtak0trVP1NsZbV1K3uLinXq8yvpRyzTrSaAlXKnuJQ1QMv8UaiIc85zVt
0WL8x2hLPgZUH5UKQJwCKOeAJooAFWWNmxAxLnyr0ZHAAh09hLl4tKAqvOjYx49+by+C3n2sYtpv
wKXPX0lypxyoctVfZtaXWGjA2ow1aYFOA7ZbXXuy65ydnRJpEN72U4W2Rqr/0DO6DAndsJbL2Ezh
PiUXX6S6bCIebWZPoGBrmzk5hXkVd1d/6ZEsJvFBSfOl/708SLp0V/T7o4IT/DHlJfoTO7L1PvVO
KDaHdBH6FEMznJ2KEnXnLkRHRUn+iv5xG6d/uEdy41sBasGRY/A3ysBvGaDL8eOuuo+Q1HHzSK9L
sFZuTSBP15rAp3eo6h5FZyuYZ4olL3FZ/DYJf/GvVcHN4ZWS8BHwOHHEsNuGWxINOwpeyTPb1iRd
G4YSzRRuIufc1MjfYGekrSP7EA7arcueWN5sZanP34LlljqqKVcnrCyFHcnMzFaazBilcAPGUpYZ
YSnnDarLUZbNpuXL90tSCFnA4HqJxeMN3vOOi7qhprm6P+rBTKdz6Hseun5apA6h1oOuTGFeaFsG
f6Fxvl/70Xmu0NkOUc1qX8XuydYjR213KML1ToyijOZUklgjS8HPC/7IrtuDN5EmLqfwA/5vb4rV
pGjBrbwCCD0zJ/QUAT3WfbpSK1DDYjvM/T4c/JE/ORg7Z57+VYo/MV8pDFMlfi+BuWBCzB8xkiY4
1g3CalUGF+vyjeJ6vlfiFJKwx4VRK3B7uyKJs1+Qx8MUscPwvDBDdY5D8TLElgNxRBm3It2c+TEb
rhJkHOy1ca2iIEWD12ygLeDQyhVp4tK0gOJ+ZVdGo71NZPC99vFCyCoXbznrHClzK53EVy8qKV+T
2NN4HtMadyyO4+bw8AEXxJB4aZlXNqySqjgOv9k9LNVQMOpCwWLycdAoShX+TkWqpeJp4BMpZ2xh
ozJCLGJGc9nBjTRqZmUWkIzB+noe9RZmwAqSByoNVxAJAARekYQ80Adaf9rFsTNVhOj8SCtyz/Y6
fuEOEuXP0qfdjAzAa4PqdVeVhUHYZb1mXU7/lHCjOG42VOXIJlcjcqfpIJkxVKJWLOPvF0RaWiV0
8SHoGNXh1D7bd9jhlQ2Vjx3nyGaMaHyl/4LiF4F/0OB7S4aC96ox3URWkjOtcIYPicbdm7/6+/mK
u1QyG8GC72jC3iYgI5f6JJzYp1Y2OmOJCWUgskoTwKoQfD1TePN+3fjW2J02IpITwFm645l0IKpo
SzsOKWB/qv/Wx6SeNYi7sqI23CLyeqJiD5h0ronwrCDuXbkjHCLIIoOg0m3Ja2sRE3HnD8r5wsTE
Mt2f2zxSoHNZLBpNnEBTkkFKbXiRurZGwYKMpCbfIWvk3VuIObNq+hCO0Yp9xL/kgGw/zAEknPuY
F66JU2mO2SmtyjurjcZpNvYR+x7LYMT/uD4gva2vpN3hyYZBaAxl6yQz6SEOozuwAS9Yb8vz9rsY
t86uZxS8bOswHzBgloNKMYDl/FmPmbKuDmTmArk+mXEAy+B9ET4MvsUoCAb9ztCbasZwoOhJZX9Q
vpMLxSYWXPOfdn1LodLwSdNflHHisnS28i150WdeHozBWzW372NbE8Bk3MenpNuXK+k67DIrbyxU
4zcF4pGf8VQpnSp/wuT3/uq+d2OHwn7LGpUC1kR5XCXbs0+WfgAtrAYebAt61/D9kBuX/PTN2ocU
ThAFDlJRT90lDoweyIH4n8Lvzta4oGchUPnEDhqaz/wfb6Er3gWo7C3KSK/E1gfcNs9WgW3q+IDo
8j/CMkI9kTj7W7veL/XdprbjDqDCWnx8YBLRWjSrHd10//FgMNcm4xuhDSaFz1D/JkvCNzkdZq+B
bKMKZHpNT4skh61nijeoyBUIjxO6uqtRFNcVj9l5RLkGrr4NBCj9ECWM6gITLjGcpUM6m8fZlqHv
OhXmQdM0IUlsM76YutN/0e+78uhm9OL2dTGb8NX1IMCaslbs3n/pwSMHI78aIjJ27g9vV6wNma/E
wwBreS8Y7ojAaNRRQCsQuerOkJDKwBBr0XFncdW4vuAvFbmEjEEI2HQqSDpcl/lDcVVHuHt8ABWe
v75kHc0wJBd+IJ5fAJcqUboniq6zYJeNpImSmqwFOjfkKEdnur0kwSJevb9x2ngpb+mEuL1XvUfs
IZ8rw6IJideX+8gU2KiW9LytLqs/CUOkdM1zQonoeqXQ6oJi0whEpdovi9t3vNAmkGxoz0+uJhen
ISSo1p8VSB4fvUr4dJKtK2765AMN8qmWG+tW/hsyjwipSZK1uLD347HB350uaUPoScy9TYmnrt8f
AkiKtRD8CCSZyE2Y7tNgpJ6MsSB+0SofQXY6S8bZUICJSKoldLWK/WZbnTCUrFUc2oWvP9ZUgx28
en7PC24LlP65xp03PiR803/bPP//Z8j4TZ3DhfhfczkRzfqX3ZMx7mUHtx6rPZRYX+Dc3PkUEmcE
j6heLQpX5wymi0UOqQaTRasVvDFyAaVIqKkE6rsTkodLna+xi3URkpTbF2XJqMZkUgU6PRdLWo5e
HebgCMeaTR/LQQXYGhUwZ/848Qr8WLBQyGnt95Vei6Z2dofA+vfKUXKKih4nmxMV8I9iRLSHHFOo
Z0yGJIZtL1pHfjjYilXyVQvLkdgDgfh859pd/CdUI92f/H26+JWh/qGD9oux0fxx/UXPk3OWrhu5
LRnGVqpnMsQk5JkzKB+b9qzh6m3wNNq4L/61Qb5ckuwYYTtPQXiSoFs+d0F5BPWCL+f+7doyCwd2
nePyOqi70sVHNRbe+CjzaroXbEqm/3E2fJR40o7vUMB5Kf8GfY0wpvV+waF7Km6BIbEV8IcKcJJG
rzXcAlCjd8fGogLMMaYaQHOyt5j3xOX2T0yK+20HRPbbPEoxKeAurgucMXF5+bdOwCrYGCh3qk+I
knzbFALXk47nsZNZA/P8gopTU8Ag4XjbxU7zkbIw8l2H4KQz4T+pmabcnbcipRUZNVXhDW6j/x3B
puBgV+UbTe1NS31Jeu9x5S8PrUE+FAzi2kJ2jZsyt7sEdOWGK0RwgfumSwx1miYeN/H3OuU4JpzH
c22LEw6s0D6eqffhnLtyWuum/joyRmRyOUpUJGH/93Vd10RPtwZhrLEk2lQd0cfab2Ks9NFGrq1Q
k3t01LM89jARQ19nAkYAqfFdX6MjbzXbXI7CnmrUfIQ6FLklAKLdkZRTWviWkF/wr5nqQPOxj7zi
TUF82ZkqpizQKnXcTMvy5A1kHkUKOTByRbDnxvnMwc+CjuKTreV60hFZcLvRXWQ6uh4vcew6KfBS
5JmZJCe3hBNO9UhbvnQBUk7xUJJgUA/Ri3SK++gQVYtv8oiSYp4BNyTSY0rVqeDUuXaWx6esboEX
QUK9dfW9foIt75wUxuqu7TdA6/hE4mVlZ7Y8L2jRkmqxZ/fi2CRzHnBEYAf3z5YKHdpMw0+i3FFC
GFgW0hliUF1WjXxnMcaf1NjPb32rwwShV7nLvv/4OKb/jIEZPUjqeiNCgeCSXXJVsy9UeRv7RSsF
h3LLn7xMeR7kvmyf9UmsCiHZbRBj90Er0lcCcA8s7kgDtvxkBYxLeDnrlt5slqXmBFoqpkEljeW/
IOaJyat3Q1CamenfTtUKZyg5dYqlR09WKRePhi95jyvJUTnCEKtdqGEMt+RbuUWJdb1YWZKqBPY4
af2C5iusTN4k8IHfFOxHtfnGjn2YABav7+nllp3G7+TY0Ab3AQgBBvMfIghF3mfGeBwkj6NbyD9/
NwyRGiN3Sls7S9QvOgSa0CyXJopNQ0hU2ISIA1dNOFYOFYfhNrdIXfLcwiva339Fg07doRWnicfE
gxyYD5M2FToWYO0J43FAj1ZiJg1Kh68lWfOvrsOBIUDQfcFtL2dv06z7vDBuGgsCvn2DvOMJ4MXm
GSvJgKgFqH9yj8w5uhSOMDFtNFwVUd9x796y2gIqi6B18syNX3g2RpKPJHyZY1FjP0d1f56xCK2e
Jh7x06+5jZ+51MOL8VVJDL2WwE/U6U/QeuG1quGQIcyY815o5fTCt7mapv8zAkny5bxOL6JZNFLh
U448URftEzHANbiewAlK11S6G85eyBXwNoQym0YCJPz0BjG2hi9iKLkjDUgE6GMTCDAjrqlbPcGp
oKjB2fXvKEiPcN9cV/4pXMiyiYlyyBDESAiE57VlPepKiuZ3yKlbBb6A6a4ifRhEc79L+IxY2ofI
4SomLz3Pyso/Ijuo5ZYqfGzENO17HtfPSsSOPz6nztnY+WWOVH1QYR1ltAbUxrg27nehYCDqPMHz
B4poxHTjEoU02fgti5ScRGpeKu8Vt9SrV93PxnTX/p1nqR4WbWqcg2bhlNG/b2gvGMZDS5ycffy7
HPXCz1gP16/LpymRkURXxgzdZPHU8rnGy2+mPPTsL99vhMxWAkzujk2BA5PYETG6PverL2SIsu0J
lt4caPeruBJXwJhA3JscHqoty4wfrCcpcncybQYWjYZvy6z9drlujiWjz55BXUSmnB/cIVJTrLe1
eX6GrGwCIbMWwtc1JnvGTWB2HnUKBUkitpbay3USnzOXe+/02LVdh54tEaNUyXhodhfSj1oR2KPc
GYAAoS8+xX+oKgMBZs2yfC4Fib/CVfqwHBNlDovf1s8oOuT5CzQ42Lve0kIs8cz3PdHmBhrBPtW+
aZAMiI0jaPe0Xh5z6nRNX52HlsFkr061+tOob55OOUcM6/wzwawntxSAWSLMbj0EzEA+TbCvP/xt
JQy0KApFmi5YTQVwjd3tB0ukx9laiL2euCoLgkEdcIvVZBF7lTXTZgdWMlmhPHePeGM1taOIp0rs
gzLF3Qolfq14AeWfn8mQnbUMAS1OnIUUt/f8PGtLG4Gwg4PuKeDUOLIJ2KfhhQjyha8pTuDvkj7n
kET867JSlu1azG9WcPxIAPD/wBbwfokK5VTYsNaR1sTkBAagZxYvO3JreU6pRXSal4BuIFjPcRq2
w5nbBxvw1uHaX7Zxc1FLbobfXPRpMniIbwXVDqDXK8ANNNoc3uskX+1hAW1UDKyhEqJw2In7FQ6C
4FMzsU5lJjtv44FLYjp5gC3KzAIRRxGYrgCnUOZwQTwXnrkVMG3LRPwaSviayjiXZR2A8P1LzmO3
ZVM4As+5Cfw4s/DmMIzShs+9U1fTLyFM3WPyVV8znbnZSv2AC7zCMc4ip1+bl1f0l96yEHlDLsrd
k7YfU7EN6wp+Pz7798rK/MF8Swnzei1M3V/c9sPP0ht3K6u875h2YHkRXZ84QackGq//3vIheReI
L3d7nwuTOpE+bmWsu6SIJwR10YTSwcZiwp9iqEOvKsC17tq66aFzHei/1UsLKXCFGcOgzLLryvBg
bh0gXjRENtF3eybl7oI9wRO9oPCYvCAm7QguY3zwTikVSsWIk5w4d7WrJI1UA5bOWCcX9bzfJptM
x2h5N/1tXgfGt06DBRJ/ox0ZrqTNB0peeNQi4IyVvlsj/uM7i2inIZSbcIvxuOFpYYhdK9nv7F1d
daRN4iz9jdYyDSHzshWrefj1h3fVR5bVgQag/0Fnx39OBs5HsrfIUl2ZhmS7LS5qgQ/uHuR+O5DQ
HDPKkVvAy7f61jj6eKRc3SWwBwkcDyx4wS1h7PQjAxlBKJpApdhkiLZv/MxrcGd4icAG7cRZ7i/9
rGWHfvuBMcDdccoJF1E4mBOb0rllWwNvr8y3zFCg/EZ3VK9aK0MGN2ogBelhn2iPCb4BB4Tf43rH
Z4V9i3kXq6DBC5fR8mpLZJJJN1B6XYTjv74f27YvmTWWSthlnEwz+BqIH1b3OFKAimB/GE9x5Doo
xHeD9v7Inwq+1vp7+18W3FE2DzKnTfOMb8vPf7jk8YiStA+L44H0CIS61r/8a8GJGgvuEF2LbI1y
KlIPdco4PVNK/px1X4ojL/NVKlbFPOFfyJlzotlhvS7vN/7ZXe2ASx4dxlDu0S7lj9K76i+lxjkz
5wSbf6jijiXDDsMG0Av4RR4d/5UMyWsENUOYJwzLYvlJZtVo6a1ZzscL4evxicQWKx1QoBwr0fxK
qzaXoewfkqdfBiM5PNjeF7o8y5UVq14NgEKQ1vESI5oKCannfWCvcGGq1niXgvhT/wQk4j3tPthQ
ucRBd/fqWpj0HN+9KlTgfD+Dg2m5efNDIWYduY0zkDTshNcCKmThD54Be0j/rarCJU4msA+H2DOZ
EakIBSeP+i6/rRSKpid4+aMBfaoPMcKEMEYxW5h+/2JsMfbJ5s2wHUW6DlzrF5EaoxjHRVSGpa7+
6GkiFGucgVlTjyjIeS0hdrj02yV+zv0k57vCZHS1vOhS+6GdLSBGwF6Y2EFjbUQDL+AYg1RCkYKT
4tYRYhA6bScTWbPM6l2fFx0L+KHC6rM4f6KYRUDckcpLesEEx+RGdeA1HcFmlp7F+v5nHz6mk4UY
CxAebqtaQh799lf4Axe9PN4FOr2+ofDD5Vyxjr7uHQJI1mAsXzB1QRbz+bXYxclZUwTH1R6yTBn0
l6V0Lsnnjd8TvXuM5mLFenSlW/AEnwE3lzfKgCWwQ6zO6AMkcyQnQD5Pz2SlidNEorJ2TldZCvLi
wKvf+E3ZQQSDbiy0/t6gpL/gNiT/YWITkx5IVw3ACsQf4KzJ0bmuafGzuN/7yfKV/EvAEPPL3Pia
Qi/H911dh8UEGxiVVdwFOfQIlr0ur9uP6kDoMYm10hxKt27pzH62KEgxHFR0Zwgx4t6j5WGrzn3b
jGuOfBtlxOuO9ODAe818067WrZhd+LO09Gm3d5YW9rdVhDE+rX3aWxeSJcvh3u3r0ZyB0X24iZgO
zDkNLlKn9Tg5QPjAkgGOuT1+1iRYvhAVxf0ijYxGU4HPjo22ffpNxZlD/3YJntz+fMLbxaQfoEr6
M9YDZcQLSusZhL5+fq9k+BAOB2btSETZLBK5SQwgThlMUiZ7J1QQijTRkfR/+WuQQTKM15iIFqDw
cOdBYbkMhrmOD7Qi8NYPLfyH+QvVL2ediiYPdoJpdcx1avmW/tCNG2RAD1n9M5EsjS27vV1yOQyQ
GL+ZwlmohG+i9aNzWDvre7behTG336yipltwpAzVKq+EisYeJk/SzMoWvSshAyTJU2O0hQRxfi1c
pTRej927MtcwUcSGkFt5kcObtelXSBBzn2feAFJLxSsxxj/5vQK4BhNYXkGAeo8igodd+1+RxB0O
xcEFBdyHHjeSaIKxKijaqIO1VldK3/KHAJUkst35FYU5DUPOWltatKZqCdfAr1q4TurQDWeFGVmR
up7DSfLhM/l0f4H/zJzHEsVLJ1iF7qLo/s8GrN04CTnuA/CVKjrBhXGFdwM1oqR/p0DZN7ZOZgpd
ODUFZETD7aDFeEy5wouh3rQm8Yj1/YL2gKWrl82RInXsh1ioxAQW228hGvkB2t4R+YG128mIko2+
SyEkJ2xgdWmEZ4LbmkQYAH3Fn2VuQjLJbLpiJhX7xTOcYP6xGpTg4H1KJdJUf7vjqzuaUr9aAMil
mn8bksTgfJXSSSkxtJVKdlX8WBjr03/u42VACrLv6c/eMF1BEXplHmwevnllHUqKd1IcRpTnQ0jg
LimqcmUwn+aHhXhIlmnfNqZkyiEh34EpkY4jeYxM/Oag5do9conBh+o79Io0qItlFdmol39grOFq
HlqL+/9sJbMKUJ2Gq/CycXYLZv3VgcwuhsLS6kRX5XYrdZnGiLqLVSDY3C/39SsqBYLNhKZfu8GJ
uqqL+YoeAqbItFEha6k9uNnWr9okCq9Nl4V5X9Tc08dz5Ndlz/yiF3MgIZi67ZHzFCmVsD9r9/vV
HaiOZlUQVloP7ufru+hMN94Y1bWomzrbShfbKTQejECvxsXWOsQK/5S1/mdSpBw1ctaU75nHVxk+
bgCQzaZNNMuvp0OmiZujh1yfHc5355ZU38myRUS+tp5xAcaViwokEe4xpYxGYeilx8Kz4z9RMi5z
LstmBwQUc4f0foXBKjjtH+v4PQMbaob5XJEvprwHqvOm5kjAtRycXMje/ni4P3ZgbNrnwyNfokyQ
sQNxKXrZnODGE6KkhxSjJjmsPUXgWNF3U/OYQc6pCGE3s9VJ+A/A1xX15CKsx2RXgTYnaRRPME/V
V7YOn5fit3bSPBTaWkUurWQRshPfBfNjSuR9GwQ0ZY9ApiF3dCi7R0ADtKpUUHTUzVGmMJ1olqNS
js//DKl4WmEkxTpvkWUVAfMRxD68g6n8P7XLv9Jyptx58EDNx2KQt5rFX4WZLl53nGWTNZpfDqn6
ehUvaN5IfwzlzP7DFhQtIbgOSy2KhbOZsOoUfXQfv+wW0yhWHo8H3BADnWUL4M0l9Z40NhnVNl4g
wYj3oNpDucA/t8pTw51ThRz9UyqaBB2zOQZApF+aazOfyOmT5xYq5fVd4ELYUbZtjdaKEv2nyLbd
qtrTGbpBb+XsfwlI1OqKAv/YrsBT0S8H7jR82w7xfFBoBi0CelGbfSIbf9eQku2q+D+yDVbopYBC
u0FmEVtYQNdY17nw4XrUyoX4DdhmtdHJaD9e02ldchWA+n/l5igVk9xyoWEiJZS9UzI/d/q/aUK/
EtsANWAm6j3P7Ps9VPCM+V+hm6dswJnmiT3M5G9YdKpUtVfMfCh9oFnojoW+EFc4+50yDmYyQ95B
8DgCB3B0r5SmEdnfhWkmyKhS9tFcFoVZvtGF1sBAdwGG+8vbGg/HTdl+s63NvKaJJMC7LXa/geiH
siREDkpChEjLOG2JtE9Xpvw4HeuG3DAHya9m7y3jEjZ2LYpUwx4HvbmMKyUTqZIANbQ2gsII2jZ9
zFtJRtQ89I+SRZ+ZIbDfZFGBVcKbpfG92R9oBuuUrsyH0nS8qG1574BLENnbWazJ/3UvzA1mx4+F
oVS9TYnxHaZlYOZGG6VtShwZv50UwGePNpQM0YT+/41WRD74sB3UAv5+fQIf4D3ROPDKt1wO8jB8
/AvJXd1jOq/XNbqnlV/vv7lI5pFRAP7o4boGg7X9jiIky/F4KwzUnqUc1W4HBfpuc4eZ+iLM7yNm
jcnAZ21ZcZicFiQZZiMdDgXzb8DdvTxreidYA6q63Stdz8X055mN+AZ6tKQTdlQt9TXusFxpDgyz
uubEFb6bzVGpbHaMstlPH0UwxVIrxdVGJQPxC/sfRPxhlXl4MS2PowBYXq039WCXBJ71ZSZNauK2
rO2nvzUyKW/MedzTqqvVVd1dqMDpOCKOxfCk+Nb0hXJqlP92xUHmjmUaHA55ZWWZ8bZQ5SXV+aMT
UtaVKWiHCFkCzy5IPU6RKIGzrxB5TDCBsFHYW05/BX09A79AJb6IwPJQfhHja3/XPG5Iq47hTEY6
Htilgdk2/GsuGyHsxDjeERs2+W/yuQ46Hg8WCEf8pbm1pixxADxS8hSR0/B2gITH+004VtW59QM4
RgoHZxacf9WpRVk2N2HOCInpVTPPawnhavTVhzgGoPn6LeN52w+MDE/4W9eH1JDMZ/B4i/CgoPTd
uP4R+oMB3/6xBmUUGCGts6DthIzN7+O5F8Iud21StZIQbncjyBTEAkbiwziKhKlvEKwtCFLSr5K0
eUbEkF9CJfpfAhOliY8sJJfSg6RBtsZ4DvV4zF0jQ8wgZ3btqV0DRJw01iLZ6vxOmeQh9Tti7RYd
L/CDgc7VzXKAMDiKgcwdYLo1hD6kPkBg+fFfiVvLIPBoN8B4aX6IhFk4q31HtPTd/RxZhUDIxLFe
aTDjBZnGFwdL+O+qhO3gdCSg4blwsFjZQYYUhDgduQiCrt6UaaNmacnBhjyoq++wel/+ArcdExKg
S04ecE/tgZ7EZvwqQRKFi/iX2s/FwmVHKHCvUfGZ/zvt8x+qdwXaPSmKCLtv+FAR9ibd2TNcIX//
2jGFEJojvIsaR2PXamo6OlQxVEZEGRmtkAWRX2d7OFg656ihxQMrd/n2nCVq9fH/aswUGUUbsOwg
EapK6gg652/pYcYoC50uAhM0rHdnoCRykt5dzqyOkkk/+ZDvrvoooZMz6sO8630wGld9RDbnv+Qc
9xIf+CgvzmdMoNuzvN21wo2JUydrall/2ykNu+AWs+JYUCLa1EpQ9IFrNEMaC5g7wI0HfczFMMc0
9B5/ITMLGclu3hYvkkxIv6YZUC/c5ndg6aNwqApEc28THGgtzSSNynl/FFlhhJisXu3sZwn1/T+r
DgdegQX+RVZYO9lBqBjfRqQuZZOK+cj8m/GzzwuR/1KZR0ZjZVB1eOLJIity/zbHL9c4SycfLetl
YPKq2Y2HZYR8xGlukZDoZpwbT7zUwC+OcE0ABwDLMttSwlpWzKUMUglwZgxwNpKbULLISolWULQj
GyGdukCIUjLPijjPtqawcO0N3O8URP8t3/MhFk6P+Q8pToUJ1GFjDvpJhw1XMgEuZTxcT/TxC+ne
eji5geSyzNWTUn+KCjpdUSX3+ZDAF/r7MXTW02Ki6pTHWUf3mdrFzt8jDAgXTTBl6m/a0FeIbACC
TbA21zte68uvtvVwBcWJuB3HsvcEZvkCXWNXoMwltlKENps1mc8whaV2BjIko5pBpAhHoWC8fmRI
7wX2hq6YZAQwqJcFEJcRPUYL9zdWEXf4sstNnYMb6NE/rgfUWEDvcktleIEFhdURnDZQZsjWKaLw
maplqIqqtEiVNYjjzoYq4B25p5cON8UC/QM/w2+OIysK5RYJ+86hBnpMrd7/iIJcVYMHzoDsDFFt
qPGnc3k4EoVgZZ9uGQ4/AAOHSKmZ/ms9glCuJT4Rh8OtjFvuOOAV6ot4ni7x60cHLd6SD13hIihS
ZZfpkCBCEVT78afpE2VvddL/kQvBIGLvles8rsAUykvqcvOxfKncnFLIj6U/eaXWzmLowXOvGewa
8vDh/IJgd1PJGe5MXOZ4+OUB0Zf1y7rVe9wwhjYR0uvIWaRehZqJqB0agoIoNUYObh9AteOo7oIx
tX42Nngo1dHQo0bx936UJut2dMfHM8LwpRtDiC4hpqHbrQnp7nmX2y9Cmnr4lavsKA22Lc+FXxqG
1ilxFZGkduq6JHYEqG+7vpuZLifbU9NTnjeFR27hyXI60pSsj/52pt7/z5P0QG4jGN4RzAhNQKSp
NdQwAHY1CnW3FtOc3S+5uRowtgm9+1DEUAk9FZEhdl6mSmFUZFpbDCh0gEBGJvfe8GoGupE4BxoP
TklTexlsDxKlGhN3sxH+DXJpPa8rrxvRpGwlN14wHxN13fgPAcBhVptKZ/hTXIxpDFhHN0gt1Q8u
9/j1izFzW984gOx+MTJWrogy6/60VNG1+BUcaT+EKDxBmAut9W3bAon2Wxe/BrIwh5zeTNdQ9TAy
AbQSmdQa4EFXbI5cY1rGi7NOieEXLsBauBD3+g9PCVJm65BQWjL6HrxuYFJAFoVH+ZwkTO6+7ci3
/hlh0kCWV7ehdgLDXqxrtPnLmLOkCKbQZR8OfI25IWeNi31g3ZdyJJ3y3T4kGeJFDOWAjcQwwwvX
eUKP8nc2dHwwA29+ptGAIXNTNT3jxJNhP97qHBVE1tJmgtEWwCAWaghl75D+u2Cqc4JpNIHLqGMN
kN/+uDs6Cgh155RP6TmW1J9ME0mbGVvxgM5Yhfvx5p0p884VfZCcd9jjG82/tbqsgmY2ECl0Atfx
F1IBcuw/tV46XRoPux0muZwWQVbCfBovuKJ6oyEnCT0zf/P5B5OCSuoH8plcpPVBHUgayTM+FnQc
FPi5IyT8bU51yMO6TfLfEHpbqiE+UM7cQT4/G11YHP1GQXSLq9/F1f6+KuXBUM+bg+XuThrnwKcu
HJBXP+l7JlILad+CuKqfKTb+8Bd7skYkEUk+riuikBmbWAyaVglxWgEhwUzoqF2plqkjtil1aTvk
8FOf0zOF161OCK6qc2Ek72VqtvbWwpTPY1BjD3vONJBEWd55pHnDIv7aEfv38w1wtS6pswle7I94
lkOzqVODAKiScCkFNMHnAs55UIUU1WRNU6/3dRZIXn34SwZc3hhDUJx9hUVf4WmYYZmLdFaTJp2+
7sTBkohRB0ZLy8hn6l/AKhQJKE6D8z56cCNQad8YcqFyEvUfbvgNyRKONHruEygSH89hG+Jy3odr
pTCGQZY189RHYCoFCm2y+dzVcKjKmbLaJpIri4w2asENDor4zL29rDQ7ktT8AYUhpyCxhOrg1Kae
SL7EmnM5da375xL6blHOX1MnlXDx6aBzmIoNkQO1uY+83+5s3GZJ4/rTNW+r332ys1mZRjElqMNU
X6qijElUUNpylz4Pgy39dtaC8Rge13UqC54s6O3jIjRgHnNFmuUyYv1waCuRP7FL+7bfSn9T8WCT
cX6BH6gwa/8DRdY09bHRyov9/UubQ/j2z6YWCEvBW4tTaqc/JpLQ6JT2aWnmwwZ8rIkySsqr6+nj
Xyw0l/UsF01tXUJLWUG0NPiQEOAdMonmwoQLe+K0FC6Epzsw8nFxWyUB15QgbQbEvBZpJ9ru9O8y
/6ZC04H5QPx/uHTl1405Yerghtl8U7HzKdBiVxfmwKQhxEtMb67CtMxlxm+y2dE9zCbW7gqk0Q1T
2MwF4L6GkdDOsIo2O9gFSz1yUUQuvkCqBHbcbSnesbr//dYuJgrMgQhf2ORGQGsZFtcS3AXyxcJJ
EDpILltGNNwur+kPOreWZ2QfGWGInxdTeTDMyO6MUsL1r/6puW2pBd/xTrehxGK4+0SUQ6czhFm8
bcMLv9ZDAlREcfMCwQjsVv7mYhQsE+ofrO8Z3OERPZ3V9AHriY9syzSaVt6/GXZClEK5bVf1tZk1
4sF2O+qhL9FIJsTOBHBj2uN0vWRPOudGpOjBfmPnnVScf3kYT5Ky9nLRu/cnsmS6ICbfdOoL2gTD
kps8gtbznOXV155TNop3MPIzSvEYwKbuCrIqZnzMXQ/PqyYdXIcZW+rO3bKV9kI+CAqH7EH6r5hd
dYA3AX8p+DPW9hmzycZFmn2qnFbBgjowkIHdsADCrbL1dpIynbOnBg/RoBNN/HjFp2I3porx4LPS
4dj9BggWxJlykNKIks7/fOQVF3kZuxcl5LtWUgVHgHJaNlJ24jzm+e797nJVP7pSOoOXaPIxr134
0rwr7eNwK2xwdi5+b+lS97goAd/06NrLIW+ebZ4wBYVi4iwe+poBXhjRVlePszT+qxQG2JBtS2u+
sVP8A/L+yB0x5Gol1QYednA7EeAQygT3mrRhlO9kNusicV4VAunoqREaeXxUB6IMoRV6vbNZqb2V
ZkOZ2zo2Wl/5hYVyvsHxj9q91Qx5LemJOAhCg7MU9Jb6YApNNvhYt2CMReSr5vjYicAu0k3sC4On
vnTZLkOWgJGc2+z6hHYFFfkKNJOI3J0GsaM+UBQYwb3+evImreEcgZGLCL6IM9PrLSPgZwn7xyqh
b5Pg31MtgMe08CZ9qSBdRe0ZqrLI1PMZnTYG7NyWnbnPpbbdANSI2fGI24j5NrhWmMa1VmN6MTSY
iQTDTOTazWZ1zrAWa31YvfZi4kkmIakEKZ5Iyaxm6GrzHAv5xxgt0q62IMI+2B3I0DgDpBJdKMWQ
42ann0ydn1t6oI2HyZiYmWRaAQxsCISwA/bvMlyDF6OquluK8YXOsJGaukzOOK5VtCUZcVj6zfaC
mtkv2FHBkBn/vNezC/6cA3zg3XkSVBbT7y45m/IIuvOYsE50rzao+gqT+GlaYfYwEzsZrxV+qauZ
WvCiXFjSRB5inA8X1D2j0GIUhMNf7A2K5ulDBFpfoejHgsK4UgnWr3FiHZo5cTExQkABAuzazOaK
1JZRxICHImhedg3cDIoDZ8rxj2TDFfhzs0itPfNsx4LYUQm1mFpW5TVlNTqVhASGP6UBo2wns3N1
/PSqZvHo6poxtCviSq+MeHU8uqtNauPEUsw8/mFgNxbWVYvHS30qtY00KaymuBn/po67icIHrBC+
RnQGmQD2eOQDnC8oOkkzYt+14TTlYK3xVt3BHPalNEh7tVDG2zja+V8veuGhSFe8dFYe70r0XDQ8
AO5SeU4LsTcRWtwp2bEHpkqNEBMknwK00X1Q0IAkt7Yv9FVb+kd3+7K4AnnJfSfio3Z2nDhxRinp
Tg50PMV6QmDz88Dp7zQDLZmzqJKfU6/FSx81YnFgFDCfdv8W6A1LUv0t3cbjfclQNPGKVtlZ0cPc
JPs9fDjmJJqGiIbtCDJQiHbAO1Ez+nTrtwNeoosdsTcH8tPkGvwCsU5qONmHYbLNoskPJ1iVicPm
yrDXcZgQFxIN9G3UxsbXrY21aA2obovc3gFzW8moVk+qbzYY6eIHtNsPfNFYUJ8OKmEbSDLXDjKl
VbPJM2I+OuQESetyGyg1QootLHuqhA4V/TOeSJ0algwvdez3O8FSUUM+TrGV65nJUhmp1zxIy3jZ
FsHwFLMrw2LhPODuuF2WTmjqugTjkHgHPZJj3ImLHr4Ml253ICIq4MkdmN6wboZe6kFlDPfC+ZCb
FW/cmr/xOafvlx+yf3qMaLnMj3+LWhDJCwYfjFwgu4QCwDuhTPGiFljZV1hKn3T8+oTTSl2UbPJo
muAsy6LyJAfOo8C5ZL41+k5QkSTkemsSEMqjn5ifKyT1PVZPny3kuTnCjHWGRYnQROlRdzsa0lE+
lORrP37QXF55xdDYWmlG9oSR/Axu1CAd0SYl7hTOxbarpX36BpnpJplP3pSXgUag+jWhN/IsQ9Zk
otv8QC5ydEBIMG+/VvDyun+8FY90UftEnDnM3z3Uay9cSoMbR8PD5I9inrPGv8EZYgmzw4grQ+VY
FdoaAG1pg4tB3GgzpuKYUU1qwvcWm1Lqf4fJUM7fhk7SeIbweJ+DWGkJnc+5ZSArCmByWqfMv4eK
WcQqbcgYX8o/6QUuKOPAusVz6FrVJVG/Qi683Kj5OjrbZKgoLHNunSvNOqP+7TwSOMOUKQsB3o5o
wTtqoHtX0hzY6qjVUjcCLX33NCry6598euiGDAytvgJI4m7rIs0Z9KNu/nVh7UqHEFHSbn51neVt
t3F3ng2/oanpfCPrphXT7Vej4tmDUk04xq19pvI8VplHOtKRoojWHh14hCMrLh0y15ym7+4bz2Fy
JD/qxvJcW4kKn7kNAakBpE729mPNT4G1FhZnBRLxS+rPthpNmwJ5/UKoBnG28yjSj5vkcnl0Z/oB
N89Rl1JjJ+CEso1k1KWQD7+cthep7QGYfye97J9Mo6w2sBNVUwYNJ5WCa46a2ubRvANPCMrSG8a9
uFXb7jfxd2pOzoQqM4d8MHlExdugDukXlbR7+BYFbs2drxIf8IrnwZKcnnWrSDjzlM18D606treY
iDJBnOG5SaubP0DjrC/WwhZKkF+xlFUUVQWUw0ZKMkKGUZGA2DtyYmvdHvI6+RhV0xaVtPkGT8Su
wyreG9HyfF4mQ30OGVP2WPfBsSRd6r4zw0IEKgVIRwBQChEQeH9UJME+XcsWmDFQH5/GxxFEpLqC
n/676exZSGUMpTpdhsbV1yVHgfbTXa0nmkeAs4LEqP7ENZFWaNBsgTeSCCWTHXypLaNK4+QX5kyh
Yomt3sh1WlTvlWVfkc45v13dQ0kJpR2XFeT3ZX9r+eYtAVonvB9vAoKX8qo5czCVhbDM7TBxZ9rg
dvNjt+w2cWRQF+YlUDi7Jf5eTdLjmJ77Q7/BJk1iW9LsJINfRlhIzwPe61KNkFUpS5jKTKxJq0Xb
88NMuRFGmS2us4T6TbeGBPFFBe0ctiFtlCSI2b/CdqkdtrIXVI7JvwVz2niPKW11+A3qasixLc7T
MocEggaQp45QG6KaWZvk3qkA52HFGno7d130LTeLoByoEkT+3aCTW0DGEHNCxk3qXrhi+y8IzDJV
USf4D1RH5n5Sd+ibGgKuQuq726eQVfqIY/qUn78lF02hLk2DPItia7kPQ6znKYg/4u4LjhnsccDe
nZwzwI79mfuduXDm5h93PBtqjyXVIMALTyASKn1XiVyt8AuO30ItZwAytDZ/gVg/heJhgmN0f8rA
7iAjafE/Y4hw4jpz1WoIydRLQmHYRD2moRaruY6v0vIdpqjVGbp2qb2CKkHZJlBl9O3F6Hmz3+XO
UpGNjFptctuyOwhFLMxemWMdKu3L3mCfVnsXgRqY5QR2t+hsHVI6QaQjGYAI+brS/jGEOHfXvW8w
gZFLI0Lwqhr7DzvHi8qMLrE7zB/QNWnIGETXs9VJyibLhFvt3ve3xcbZ8WRiWDjB4B2irHbWqMWX
EubofsYeVLvRg9cyzVkAxOussWCedQfpd5+NSBRisgaxK+VvXX6+ESh651d+LulZUQqoiOkY7gsy
QFGsH9PgqvXAzunZ34Zz3VM7iEEeCHhGbMtLHz5j1cXbwA26+35aeKDjyJ8j0n4/TWGW+1VK4P68
IKwvz5H2LKvx3w1lcHdGv4GVEhXdg8NdkRTpwfOAMegKpamyfc0wS86YO7Z4U59uQ2apFPoqB23Z
Vpg8Ek4j6SvwC1jUs6vIxv75Ot7xqaLpQClsIrcKiJXx+ogtTAA0y4y7ADhcN5DwpYsEOjq1LqXY
LEbUJKFY6FI6cATbHJY3UHFM8Bj+jUXkiA5U9ajLk0eBTGo/K+eT2D0bLFB9B10/+Bp2p2qqQmP3
Aj8PFIj5GNn4/bm4qZNNjA8s3ajoNRFnsRoL4923jZatV98VhyyT9lAfp24IOi/49p0TaA9XIBYF
hCRuyfaQkjllxZboVxyUp2zCLrFlKbLxzwcoV/w5uBISNKbvRDCCZJd/8jeQ/VrW0GmZty0dZt0Y
5pIgif4d6ULACwQVViQC6Y7Tuxnb8lZrNEI8azhUvIEz2VwPIOpnrF4CNhNoQsM2C3JzpMof/gOo
BwLi9Uw+H2PC0zSFoQKiqAW1SuhzuYo5B7hpUSneXx5XXiY3jvnQDECnRUC57VqTB9J4rTqy0q/6
FrmV5HZiXsST4msaTYrZhgbAZouH3qvBZVDMjMiO8f5nwW0JpKjKUt6b0pTL7Qe2HVSl7HBdrzrC
jztenCkg9pCXclFjSFJNuacOdiABBAYHr/fTBnuqeh9Fo7CxLC/D49JMTWUxCCU9I0/CtzJ5jqKz
YzdnPTow46x4W676yT+sJCw7XtRWJAnZTRAnDl+AoAcV9zwwNqbfwL/EsJSbZESg1VF0Ai7PNeje
iZ5hjiA8Cc6cOneXLwkjHos4nLLSj8gJazKcrzY08q/juVPS2tzg3ncMY1OHZ78NpXZYAQtRAQkL
fWJ/AtgEgRQJSSfgyCThIORyHfANkGCRA+1zh0riHVkmGI5YULoHSIpP0hUI7M2Xo6WnOLEj4HSo
ARgZ11cd5ixA7mgSsKS8OAaCDUXzcgIX2jtjbjpHSs5Z+nSLiOmRmdBsJXCa+SL+Snpt6DmhpUZA
JuKi3+1TVKBU9ESbkZa1ghSUGfplkV3GB4Z5+Miw+cUC7D6XwRINsktepkbufHudv33FB2frEbSD
eaADLPnpK83j7f3pUj0HCBgKjisy8fangKfhe4u6Ifu/wLQPddPQhlYaSTwYck7okomUtlysqMXL
Vg5mcnFJuxXspQvupemF8UFwyCCWvsvqFInRmngI1f667JBTHAbNkSc22dojvG0nyXw5a/F59yzM
MmYzFQpltpVaFRnlaqewIHXh9+0kZTgD7i35jHV6lEncSwaINrAO7gYsS6+lDI6zt9y/EjHVua/h
AYWk+5YZTr3kwkioE9Sn5TEOQklmjtLGmEVJ4XsN6gtuWBgzH+yZyx090JrvvC/sUGL/cXN/YmUk
fBox1np8TKjBXzMKXH2EzZtENkuqsYDTJC105Du5/cP9Z+ml5suB0Y1L+isFlxr6rPYGKnqIWgp4
6J3K69s6tvRfs4s3UXQMHjb9AsDDpLZ4vmXTY4YToSAnF73JAwIXFyYXRukTaKIK4RwEu76xb6zp
3It1tPlwpaNwPbq68TtQagdPH5Zc8MMuFhSD6CENNxyKK4KIW/f6FKRR7kCy1Kn103e/O+f2gNjJ
Ey1ER752fa4GymEO8ZNEez8XUfXBIStyTeK2eV7H2QOgkAPe1zoBFMOQT8h+ZnJPgeB2x4xbchq/
y3vsNO52FzdPzLzTtFdGTDa6PWg17sXdYSfKV7nuRm+FczE8Lv5kp88RCNY2W2hPHVY2xgzi9RzO
EoC9Me/PvlOkVLz8miWZd/ScBAAGmKcT8prYoQ6X1a5sbmv+skOaDTgRyagGTsiF1zpKwGAwjF18
WuW76H8Ihz5w5DXFww7QJOzW2mocdaVMMXNyCEnKYbk8pVLPd+DHohZ7vDUfmU/YBqZRgWL7w4GM
0S6veTVLLITS2MMyu6Nr+ocSrJZJ5N52vxxHPAmDIIgPZIA2bcmWdaExClEg4ppxvphEkKLZy9FT
Ga3SjhnY306A4621zpaBEqehEHe0DiM+Sv0zb/pG7J8qIRxxd80F54UabDeanm8BoJDqf6KllJmn
NR5GpQbrrkFo6pTUzFcRJXfVcNebsVPng208tCQEfD/8RKthsjDV2hfFGymK2ImgSmi6RslQRM/P
LwNgeX8MuLijfs8nRl2P7YMjKyEAkGGRf7gA/wWo5TphHg/tjQFPebB9I465QYPU2lCAyoDp6Hgb
kaPJFWOWawjYfUQ5RXR/RmPO1G8kp1OKErp6BJwXn1ezu3PUa8AtLDwf5dWxrNegfy06n8AfcUO4
KeKInr3yYHoZJrNUmuQc7SNjTUJt0GNJ1CP9YA8GLaZ7c1PuBxskKndkDVH91gdtXKWf5nH7TOzm
N/XeaKi+cAlXh34tIXnZTdmn0jVVWbowdC6r9r2QjOthHE8pq8AsfyFKibiZohVNNPgspueE/8ZB
RwiO8sRXPe0dTIb+ZX7qwXJ4vXjKA4mWs43a04hsHI1CraErX2orMB2fXlU31YDdgZmOudDnHNf6
fcbb4MEiQTSMY8k/ES4JCTcESwvu6PgvA/JCyt6q7tD1ysXL4o7IOnQEC0+wkuu7K80djKqZUEOl
EI5vbkZ8HlMziAZdN0T1KTHMLb5f8qT6NjlrSP40FwUHNUVrNraA2T0XQIhBTK/dfmdCF4g8d/LX
7jbvLnsDp89vKvfA4BlbvhL4yaIgq+Oqnw+CvomfwG34QWIdj9GHytbtXaIzp/xfoCTO1h8faZrQ
huFHJGuUNwQdVamVFUTSu1iLdNCiSiSwGm6cW7VwLbeFxW7cgKKbnW77ZUH59AFYn42zrgNClk1t
YQoSL90tg5MsDOyfOfFsRzgKue4AwsrI89Xq6sPz6uAu4tZTgKnsreembII+SxvRidFChAWT+F/6
F1m9em/7a2c+1MPx0IjGvqIFXP/JRu+oP0y5WuNsZq/5CUcpvzm738M6LA6kPnko2uFcgegZAxGY
6S+EGVoy/5evqYyZnzQLZzY0xblh1Z6NnuDqp/E3ZFsAlPGM0x/EE7ra9VwDd3DXaaVTbpdvIPFx
LEQ3I49J/L7im4oL9KF9h5eTsAM7C9FNMiWig90YgA0ESTNQMreFVpDX6R/qkfKgIJpo28L6L+mq
jPVT5bMdEMwvCFDUFrrthnlcw8Fvn0c8AIqgnyGyQjtmpxZAe0hzcGNPC02MWrhJCwmVPT0EH/oU
OMFN5AJC7JNkf8wns3dXUtUzk6qJr2tdW8QqnFvOq4IYpMF/8COpuWp/5dO+a5fWiXk/iLu+KYWV
eeZeQ1janIS5Nt//dEzpwYV6DTJGVFpfGcTqVoaXzway6NtyAhZAo2HWavjBgahNMkJ4x2nBw6un
mWHVUqvXH+NA0CF5hZ5ZqhKDGJiA3dzIo4SSV83DK5KT8BJ2jztNdCMMDitR//ZKvzf/2xFffN2h
sjym5mh9IG4blNCXfPXPKHCrua2J9vwhidExb/vw6lvxJodkMszvhocc4wEa/ciDdFajUB6yDcsq
2b7iTkcr8ABjQt5MbZhNZEHsotdjZBH/+WV2KtmyIXgCkgZFKFDPMHBcGAvgYGcSxMVd9IcaiiBW
6Xjw940BKChMeEmGCf/03rLIcU5Rw+QaPv1MkQhi5DR3gtO2QTUNZfyPHpT1LAgbGOFMPQizCag9
hY+tyOC0+zOSzW2qATZT8E/ENs7w+BIPPnehXj+o3P74IbAqMUEvXS00kH3v6PevY9xGDRYzw6vX
4TKEbIZbnbXgU6ciB5f8qsWVJwGZm02sCpZ6MEOWGXLB+jEXLwBludbAx9NU/nEAbTvtxxtN2XJZ
sCTGF89TTgz9eA7xKhkra6LAU91C34tiSrVAPQnoZt12e9O8IClW8hVNe45zuLNhogj0sQLdHK5F
y3BtFwYyB3Ce51tlhiV5XAvT/E+Ntj8wEcdhTj6zhxU0mKrW49FRZtHGwnJv7geM2MnMazKJ3yvz
Ve9o5bMtUdDqqF7T5aD32elseQTTwwmYTXvkVhCyxiA4XgA6GGTJhms3PXftrXFTtbD60D57eslT
uN0slgVb7bKDqUuGQjxbdBk4JJwQQVSiTp8RjS+Apb4mcF2hmVQT/73Wr5jKsO9fz+fBWpKBRBRM
c5fEGLl2K0BVuXNuH8HlsL6iyYJ89YamvW8pDM7Irisg0nnqp9p73J8+hdxim1ogT7n55NEcSnFs
8YW+9daUqNkxG7wAYGoMHe0lMhCNcgkT7xf3/QfuUSbgLbc6vS6nqwO7cyymsDUDdNMJlMkx9jJV
FUeSn8N7oxHtv23/6/8qVuww9FUr1w126JP0cxD4ZCLhfwkyTs2EBFnB4vS6kSdq7p7yroSz9+EO
UOmQ4IksWJNioZUHDwn5fq6VR5CBFzHeRMCQTpor1/xWHjhtzeWJEprUQUhwKGMko1qJXyJABrKY
8oAYDuLwTmuQuGV1GRa15UA/jevsESVU5eJPYOR7gN3dOMo3QXSq2+CgXJC9w1WmnAJA7RvS5h99
AdpABWab3u+IkEyDdSmtBZ9jGKbzTsOdibGl6xRRAaXNmO0tYOU8ky6uU8jWTKspj5bewMrCcBWT
uIcnLmgVgvf2CKHf4RSqYK0kGRi7+Q3yM2cfgcfyCh6J7RP5m664scmqFeorZl307V0ATMb1EHAR
Cn+XDPbcVuCzJp27WMRLzmLTct8LRdJY3h+qhP/1mvMOVU/VmbGt7OjQ6bWdsVBMZLYHbVvoLxPa
weAAvbjcju/TLBYQR/7WkYNkhCkshZnjaUFKH7xNE6Ya7iNn6f0uIlYdqBo4opgf0N3+/OoTSQI/
9ORyEcCjR5gt1uehJnmVGWN7uB70GuvBD5H3NgZfnA4q27LxpzzXjph6Zh4Tvt0kLocsYHX0YtDC
UKyXR1fgeW5gqxYsMe2D3GvLKxhd15eV/E7hdSYVpOrQ3GhqVx0IgDgc8kzHvNGSG+ovlI5oUl2N
4oyWXXoLTzM9qEXP75XX+BsacyktZIeZvCR8dKdUoMRYPDWJN+POvcw4GCO3GJqpNJ2h6dbiSuRR
k2mCzyVPpKFI8MIEmnqliZWYFUTGBRrtANQ8408mEveJzMmfpPBBe19K52yhplcOxL3TearJ7egK
mnMYLRH0K1TzwKkH/qC/4vDICJa/YghmUAAfxaARebREjhRytiVhAw5f6sybHkjR0gS9cmVKl8oO
cggh3DSiUW0bRV//AcnLtM4jEKb8WqcTieGOUSPT4eirHpdDTDarvf+Yhyb0G8fbzqhQcMADdRk0
gnIWVjtqUPo2d+BWksqcqR1q86mixnu9nNn01yB7j9fmjnOpvd9634xp5xi2FVDalE3O/pxtApT5
cOsEmv5WztHPHh7o6tPcCrq/E9TkLe72ydHq+oRXwKrkmt7R7jFRin9lNRatW0i2turV8uDJlM6j
D/QyYJd4ifizzjbTnJUPYKMFCCCsXL2rNjw6L9OZ+9b8riEAFo82ud97k5wwlLf2hwB5GtwZ+S7j
eMrdzpnLE2Xp10cBCJ8deov4kiZ6imKvK5B5TBADwUb3Nel7lRY/8Tbm9h6yrt4Z0SqexdGpOjGZ
BLFcYcbghImdu0QiNayjCr3PBQn6rSxPP8pWz7PSIYQA47H3O0R8xtqSYaUZAWl4DvDPbIK0r1ft
z6DXccrCXYvCZ+mJ1JM4IzR8GTSIFR3MF+dkDFCJQtWqhHReQb75GYPOdZiXwk9Km2EjPhg4lXLr
OLhEInKGjKzP+P5ST0R1nMIX/FQGH+HGIGsH2/GZoSpUYZ/dwA1n1d5NjOuytpp3vSoXdu9M8taX
9cW7s3JUx3h54g9AiC1/dlx88PUVCnYKo6uPoeK/A5nzNIrw3S8tARsj/0mdupyJoAU+7wU2I3uf
Z2qcZd3ATWgGqxfwGItBU6pN0KdEd6CESVxFAHmLDSJd5N5GgEHElCvMX2iX7KXC2t+L73MoaK5e
Jo1553jmjdT+iaCynTGu5b6GMtIauHNjfUdRr8Zvp/ecxBap0IyR0CiQedwr+kdH/Z7tyWz4AyX1
iDFJJIZAo4/4YIK55ittT3fgtci54Ov35lEKDQURPl9pK403iFMa6msKLdHCGqzHG9AxGVWRqp+o
2a/t3GF4KXvIdZBlICcv9YSsCT/7MYjbeeReJTwQAOcSEVvX18YrMRof4CIdu26uejYoz5qXRRff
+uKMX39+EgAsvV8du7tGy0OdAkVf3k7tOdBDaPLyDhM1fijRDzorB0EBdaNsoMXMWlF4Jr6PxpdF
bp74CE6qYafJpT4Wn9hxbz4Z2UkKQKpv2hZfx+c5n/8httfAQ5TABElQRSkpDMPvvcstCUSHpoNe
JfI++tRoyk6C0XB1HkYaBxh19sTMiMyrO/Nd15q43nSXYFv3raI7VHwnqZ37Kvw9nZa1v2YDKXdt
HGI9Gxat1J5TihC39vpUtPNhU2tfGPMWl8kpuPaWx7qBrfC2GuD5T9sF9zFOgbH5PyL+kKdnJ3xS
W77RHIcOmx3M482CpumIZiWcXii3HKiYY2ggNrBYBiqyqdjBh1B6jdBOi8p4evWjc7tC71M3Xx4Y
Dzurj0f01PjJlB4f1UNdiFxmABnOHJq2mBA55RxXPv9/mnjKtQX537t9D/kNQnvQEP79x/MYLdaN
SXHJTWO71+cKOtVS/SXxVse4rNN0TydjkpUmq37n67r/bphUcPoI9vq6F7uGsHpec2SvZ7ne7IBK
WiznXQVuZumi77922rze0XOI4IImrL2nztY3tLEuByprwE5WslDSrYW2IrJrbIU9t0uowmJXm6DJ
7zxCio6frnOqXhf9DVI2uKv4FEpAg5dp/LKPVA3cwqXKPVfQrJKgzCADHjzuFu4KoBiFYUHiWk8R
fQmBghj+WNu2Gn2nHdvrUOq/Cn2yMcbarq+kmlw3UzbTwzwI4Wnj8NnkTs126W75I/KDIkKQp2GX
1cRTynvs1EheDyPXY/TXiYC+1z83AdCNayIyDSrK/lLCK+h8VPX6vDuuwvt0pjUAo2Z/sU7KPJOa
KeSglcbHzl7pbvVmPC17xHQIFGQICn0qFv8oQ9PYqP+wPGa0b3E4AjRbibdZ2EA9KjSV0OQX/l8E
B7svB/j2Ly2uIpVDiQIYc4fCQDYrGgBQjMcmxp/RNBosb0UexFodRdYfbSvKkgk+/Jzt/ep3Av5c
y7uEC1Hcwq3zx3DBuzK433HFKJ/9qrzoJuHfbyUe35cQzQqZf/KWExrTNsbZVATmfzst2DJnntj6
4Qnf7wcy3C14x2SRgZz9YgwdhGLrXbBwEI4zjCxqPoSY6JgFczTsSikvt8B/qJmekL7e3m/Wvr4S
MOkuX8K/QW5dSQy1DRwMPUTO9I1UavbzbWzIb03Y9jvYR9LKRl1WAkRnAvC69ifhLmEclePGOr7t
BfdFBT/jR+HsWw8l8gPiL7ecH92KSknklF7hl8ZyEv6QnX+ZsdKXEXxiVdTuAh3HkUxJ8QjY5deV
ufpmwd7jerIqLsYlOW2LCe9JXavmmfu/zFIbzNgMgik0CiDvmtHQPZrVj4T+MN27NGicQsRTOojO
QclYgdIi7KcLgLQ96qZPcVIimLWCESbs17PKQPxOO1Orv0w6cXYzAj1hFZZ0ZdYDOmjHO6VsaOOZ
QdWyvL3RsyMEmm0o/xdT1JEAklZXskIyli3PynKbRFWJE+S7AvLYkg+lrPn/yz5E9Wrd3dshV7C0
Hb2jTvky8yLWWpw/ij9RsrG23hO2rcFESxanpn8mLqcZr3C/ky5b/1rQMGNVTz4cuq+5EWwYgrWj
Eiz6Vj5JaLn+w0wZS/QXX3toIjh2ChbsljrMF/DNgWCXn1zsm4+FIU9G5Iwr18rOwrGVmXnUa6Jt
jFFLYhsSJTzCBjecegLBHsmCDTjjjG2KjR8X612mJ1Zi1NVpHotxMwwYGhkk8M4ztz4MpuadMKxW
9yT4ygW6b5BT6TMRII2GphU4EPQtUJbC2EObXSuox4/92WuH4HCAtlUCl93G2rGDypu5msAy8YmL
r3S34UJk4hb1i5TjZ8K46MqjknxYH9FzncxlQXWJzx5ee4otDoCBhtKkjhIa03acBvTqrBUeEoyc
Mc52nbB3df+PBwheAyHlA3DO4fqOVa+rUJ/Ru7v02hpqg6ziZPH3marnhQYCvaTZi28sqqDj/Yq9
3zVE9MCn8PXcxUD57Pg65xE/p57R8ljFAvMVO+Jd5UWoezE5HXb98bKQ5E3OWah8yrqxeQr7ZKrK
Sugv41J56yMZakX5yGfIpTP3sVxB6iFY6N3yL6iHeUtUXbxygzeruszqwC08DGBKi0Dn1ZFcmalY
pp1BGedmKkOcKd5GlW3hcM+iU8bnVsLCWujlhkpQLvPVOHr3zfTvNoCN9Jgt73CbQsS4dX4YEIUX
uNe0ovcvnVVB1MICkVXBUr1I+nbGc92MRjXNk1R3y+XT8K4DCEnwNa8hbDiJ+P1tD7dTib4OcIdo
a7WOvmo3STPWI/v9Sl1ShoFo0fXjqvmvAoEL6bL3aAi3VrjoOZnGoHNGoDbN71jVu4S66uon3xiA
jSyfYwC7AObpvMK5Zp/ABDHXn4svewEXDAun4XVdAEFXU0+gPnBXsbjPlcK9DOgIJZgTtuapU8g0
dgiYJZi8PlDPzi0hFln581Rn2Ku8XsJTMt/5JNQ6v2Ne+q15JAlpmPzo4YYDbSiwtYBNl0LaDS6h
rAfg1VK0tAtwpX7E7hKQSZQuEfXC3jUxiVzzUrkYjZnoHJ5FCS7X+7+PMRmM/nZsp3txShzt1Ac6
MoEMOQhT9Ip/vX2SX9UOUz7QmCUTD0GPHrGSQCgGIGb6+TCxR8KFVTzcn/X2hNZS17xvD0LzpmvE
syAQxftjsLQ5iCAFwtVG6e6YZ4MON9msFBK1g6SAMTn0zamaOKID6Al9XKr7e90vaN3SK3T3xU4O
vTJ29zT8KVShEZxR/sOLZDMQkuXVej8CBYzcpSStJ6svVebgtYPRnEI7ILtbscNdtO2Oi7B06ZMF
GI/iUVBVzh9RTyaxH5D1MHUnIAY4LA8SoZr2QqXwD7Im9f1o/hr0Fiqhh0nmLOas2JxL+40KbW+m
DoFon8uJPqcXaVLgYr39gUP4hmeAsTs8gOYfo9xPiVE3bhXnDZ3PQKab7x2JHzbXrI49S9SZENzy
GPNwbn9KjG0QEt+nUks3LJ3y59/Jbz6kr6coGyNWoteeZ5aeQ4tpa4DUhSzyZppBELycv0TTMHnZ
ahOLmmu5e8w4x9tXJv112q9sSIXCASID590v8J/DsWAO2wtZ4BGFY33bkcKWtPCWDupYFEew+qiG
sSy7pQ4QLcqvZvMi0U3Eay74dwr6jlGvn6iYpEMUO0zYzlZ9j/LM76/KUEU8C4phAW9d/vZo8hP9
VQi0G9sGzurSXAPihXdDr/Wx/hc+YM87jATFm+N0/Bg8PT0I+1zrmm+z/FFRW50wurpuSv0P/h0A
USyJOeXZ0bYGHXtLJUeh30wABwadYBdqEDvxDWsD30MKYWwgdTkjKRMAWtcwZvfd7FYzFNFcp66q
db4ygxwwXa9H0v6MnzX8A1GflTqg/UF9UgffrBGpKeiaK0S+oE21H2iRU3FPvUNK91woLCBhJNdd
+v/F+7IMjGLqpM1txIXEAizqbOpRBgjcGRtdWBdxVHBCjbiT6+7Ck5gr/yDgLZy//0v+A0fEt78O
N74/bTFfQYdu5XavJeKAFdT+wTSEuwnB2CyJha0aV1JK6lppWogbWxuJI9b8xUOJa1Y8dLqAMEbQ
J0ZYi4RZg+orxqXIBgjKXJUV3ER7+O0qt3mbZglFsiX6Qou2a57Npv66wMwyC+WsPuynLXaOaKLM
KqaLL8vuOS/et+8SGhyJKMOxujdybokSdvR6q2UrlRPLsBjLh9xiReFMXuRKgwaHqIWgeZj8OsUc
wiMACvZu1x+YF61VPs/iI7500TodqaerxiJgiG3iWSu6mD2yc/SRnQUfJEhBfIgGo0moblqiTiU2
qIZb2Mlp3LZWFNnviMlMi/3ccuOk0LSL7Q3T1XSq09tDwZPPN7g5jszXjqh2Yh3AipazQXvMg/Km
Be1rxPYFFXWKQeuLBSGRB2q80FrrlpOnxuUdGf8VirrPSEZupL3QzXzM9LTFYuiU2a7f9xHklm8q
RxJ6gxqagAaU0RKcSAuEfhrMNquiMLZlQRHg3iCbXXUcl5ERLV/cqMeho8lOI9pelB2p90aeMVVF
Fwi4VyhRtiMSaXaoC5aWDFCTKz2hegjvI2EvcasA2LeWQI5WWPoAlSwIxoE+r+/OCD5Lm+P3KOzb
DSZkV5C5SdlkM4jdu8E429OqkhmsmoS3VoA3RFWB96h4tiaXWpPFyrNPhVX6dyaW8l0t0sva/0eE
isl12Q5369EkvImQZAPGwbnibDdqDcJjeHmBEsfuu2lYncBacOgwrFHnw3XiJabiIamY0iV7X0zH
76p96eGcCxflYaVL8617OM2s2pO/ka/CysJ2a7u8raBxKI+lSJh2n4VERoYeFtX+ecwmWupckixU
eF8pCKZ0jFj8W8SV8MiwFp4Ci4OGDpi8i9qq6stDcT9puu2DZbsyU3Yj2/wH3Xdb7Nt1MJ+UVnWT
dxF2jQTzmFz+gT/N/ZMRkXZyzoHjUZHM34VIZG3+RvL1zs/aJvMV2+rLObwT70T9BtcqTV7Zj09R
xKw+gb94RHM4tTO+2DgX3wq4gKqc2B1T74XLtIR77MPt/BuBWZf+HKpmLWWvfnNA6Nog2n0OQ8Mj
vEZSsLvAyPxNAcJQYmFyN9ep4oa8F9pwas5RZ+ovo2Dbj+sPKwDOf/SDDhoNsH1OAm8lycATIluO
hKsiwycCvYwXE1FMdRbGTtr+o2ke//ukN407/kWYOxdcBSqpkQV7ij5TS3z1KA6I4WbYj6svXPvd
uMFFKD5TeWqFoyOFD3Q86I5FaI2Wju/46RJflX7MesvCR8eqGjub7grpPEEsXxTcSQpNC0b+nI+M
+tdbgtzKJV44ZuFKTp6X9crOZXS2MT+kMOlpxvj18aLXwVIFb3e3cR+/JRTtgYvzO8q+WFVfeY1h
YrkyZCyN7oL3G4+lr1jQWG1anZVTr53f8zjH8g720sR1xGfXdGuqXv4b3vmPAm9tovMsEXb2RsHt
g+PURev5w0jX5riJtOv7/qrYiQjNhGLPq3f90FpP6GzWxcHR2hwTgjC6A4FMteDTZS/qu4dIZboo
84kZaTdGcp/7dj7UGowWCrK4L6qm85dLmbql9yLOn46zVwrdsNe7fylbJlcagroWy4fuJ+EKk2DP
Ym3FcRXfZbRFG0ZBkwxLA8PFQusftOUy/eWOCuRHrm8iMlsKnGbYNe5J16yhOwgJf18JeyDhO96Z
tB1tGfIXx75HlRc4zziiWpNCFwWnCG3jpLlXMJdUSRYWv0oU5p/ik6ZkCsJs8NpMtKYAN+WO53PR
uZA+qHVehXpqsdMJvOzVlSTr2gumW/zA8gREzwSaB4I/EnVAa+VVLC9IL4IPxpHfVGL7yUxkswjz
O0BhPCKb0y8PFvsYSxpPLcXmWxL/rZO4feaKpoFwpvq6/HY8tprBDdJDaUTylCQVoymb+U/EBMuw
0YX32dcxTee0K5Q2vKxXhdkpnqGft8AsijNBobvTpAx+jXji4F7TApA58XGnrxwbDOHtHBsi5PXF
IVmec4QKAmb2/vIMZILfWN+4eSvIMwFaUYcrUjjJtj0YA1Xzpl2B2gNKyxgCyPfWRqS3qeXf8HhY
Xl5fhGRRftVAuHl2VD4bQJ5hv+D907QbBHFqGzpL1kIyA5LbPdykHVe5XaR+cXCNjRm2ukS22fDG
KE4Ds0JfXOtLUP7fWx+sE+eMB43OuFcXhoQK5F88s7eoRW546r1q3i2LoApYApBlx5x99FrAeeJA
wp8oIYkV/6evwZDTU2C+4mzCByg0Lirl58gybzEbFC+B75l/8L21mKt0YzRRO3O4CR7Mz5HzCqvN
PBSJTlqIhUDpmkftR+vAyGJQzB5erUPNdRXB9+kmlSeXc+TRGw3clpcVWAQJSJGX8VvX8LlFjoLV
a4wXU2SdKb+vvarh1/KgoK1zXCpDtQhDFWNehvV9WqTbMOrpLUPdvWVYDqETO+6+Eaqnd2Hp2AHp
Z0phDd5ZZCcqZ85jdgVYesnVG7zp64TsR/NGNIJ+89tkVRWlEFKkDien/1tognRKqGKHp2V4G9ak
h4/GwVQwzeRj1pyZhQ2YFowJZtIjQwXNaO3kHnOuOtlaJxsikgJ5gkaPgh/KDo2QInNlq9t26GZF
UbhnhKoU+FS83Nk2OSkPkGcjL6hAqTVHiI6rThWmsrw5e52FUKhmQYyUoYjj1yxhKyNgIU8ionTA
Jc7OKsrWxdG0wgpjXmpOdiQLvCXByOtyS7taWEfWzeIea7B52HvSrtD50ODoSlpLvLfNEg3HZ2yJ
5T3YtX7esDU8kk1ZBU1EEvB0F/D0bSOfXvRqAf6Ga0aE+Y0Rk5UCkLXgLxmkFWcZ36Zt4FmNQs25
b44ohphSV2g0QLrGw/RUKgHJzoRkjX4nCEtJsO195Jz3tUXkDWeUGaIiRja1CoX6m5BzK08R91uC
2nbzF1TXCAXsqzXlGIxUH4sGLtiovNHYYG7neTihypv0oxyR0WeRnbfpMR5uxfjee4Pv6pgBoiOs
M8V+i5OQ/qyGlViEs9tzEmyqhKfW9AwH5cQp89GIX80Dq8zB3zdgf1xh22c8nJpVpcQfBQ/jc//y
o/bbq0habrhFoLar7iH7tfpvVeLzUY2wcIze6RFoGIgfLLCwdYGp5Td0t1PvIGQgKUaRVp6wFRHV
ocXWHR1tBJdqsYaRqTnDkDwA9hl9ZI3uOPVnr99AByazp3wF6OFrnMy9TizqDHcSmUX8Xneql7PB
F368Ut+IcIE4FEiFHYHBAX2x/MyFzNO4sLIm/wN31IxlyJf+ReYCh80n9UCO/zT3FOj4ceLF9W+8
WCNk6NYXPnhbNMhENmWpRjCrBrCaO5buyjFxevVQ+Y3K8jYKTBgor2oVlfHex+TPdjJlO3yzrBBL
4io1dNc9Bfj0PFnlmRZlkv2h8zz3AvttTKTqcS0iii8A4etabu5BqnnHu8RBdTS9DZKmrMMA1Dqy
xO+dNnoZ1XihhN+X2xCnPEkE5VCa2vZmFjxKR5f3i7oNtQ6azrdln5iLcKt/PlqkHhhDTYaeJa5t
bEpvGyAXRpq0d2iKqQ2+3pePFIrrVLa53+2mkZ/GA/AUDpjtN4anXYgyO2jyDm1FiejI6UIFq2kj
OBkJKaa1Wittk/RykTUaWClQamzq2DfGBU5OJlYhVXFgZnRrw2MGjj/uTcDtaNbR9y3eFOb0/Ixm
18GhC9sgWVej7bA938l/mZjN71A/4H0Oy0cL1Kj4qs6N8z/kd6ro2ulZ22zzK+WLwARwzI4e8JgV
5CgG8hG6cGmqxI+e++QgYCkIAIYvueX3NwCjbxtyln6VfN+bRB9cYEmeH/NZ/JRBH+pzvSrkOA6u
gq+rb72h8Gg3O8v5PrKqn7bO5JZao8H2udeazRX119hD2SzdGRm3g848J2GPAKhFTV9Bl3JRmbRm
7kG1WCF4RdVf3Bw/WgCmFZQqHUhZI305dp1FH1YSHP2Cv7K9ddPzy/gfT4hfjEbRjoquZVIG+Es3
rAK0vpk7UOMtrq76VrInYC1usROPlJsps3j7FFWjEFa5irigIpZ+CvmhYRIhmqXgOLsQeGPnzxWk
zIMC1+BlsGfhO04c7OPIoQiT3VIfjKh4hp2qIOx2j/8Y0Ci9Lf7Kd+OygL51cdaK+Zfpbb8HzO/k
1LwP1DmggTINmejzeF3TI25vBKhrwprcv7U8+7NUlwI0ngWIiDCXnuYob4yMzRGAemPWq00feVU+
+C7tlaPoxSQ+XpMxwEZvibzkhTbj76DUVutUnh1dTC7rHdUA4DF1HLXmnYLfvNXJ8J7BV9gjUKue
z3gL6htua5ObtLPZPQBsvLvCq9kcTQT8GHksjnMHJTE7DSAWS45y7rUtYFaB9J/PMsaNwgLHamvc
JPujPFkiHtfA0SmE17ATqg3gjaSA1QUz5o3JELHY59IOZTcnSskATjN5YOQUThOm2czxr2M9TQxa
tCsWz+Bo2nO3otoEZv/9BdYN6K149qiffv2Xlopw9n10pKpgR/7JrqViPhI0lmSwnUaiaFDURY7k
qsnq9hTcgUVTQaBRf08hgbax46qrdteLLvb1kQG2nQNihQ/U6ql1pmgnTrGaARzorz8M++JvLBPw
vKP10mJEyxdqol+fk60uEu/KevlDgHTdYfNqh+bByzxmdMuX5Ifo2YsxTs2PO8U0EMZkflITa+8f
Zu8P6apAQqDp/Vepmo9hDmEd6ERjfFj1ymRBrFL5c0g4A6VwRIfKlu5x0NLyfnvjp28VANTPHI/a
ip7SaqqAxb03n0j0VyNjW/Ftqj7Q4Bv7bxq9pO8CaRfluk7EUHw1xO/uc5uZQhsNXVVzKeN6lkuD
s3lch3Qb/7h7FZPw/z90bJn4MeQ/ojXjc8FhLvaP6wfF5l/KQBGNse6fYgORqK2qh2mi98+Xac38
+O+vxb5Xwkk3lyMh2Xv8lSMakx8DymH2xl7reGvl5B3r/8WhoK444RK4zswkUZjvT0IIpkStvsMt
oyNLIwN4iQr0q7hbB06GTgFSjWli3izV1i7VuuIGiyvc2fPUQIatNTHhbvbrTJx5XQV840dg3Mxa
eGY/TmEMg4LCEuS2BnnGAUYktqD7tgDp23lenMEgWjKugas1VRG3Frchb0k4jm9H3NN4u0QbQR5G
3m+Qq+i+C18FOZc/Rzzu3IVQeU4GL6dSk9u9sACTJKpvlGhLqUgow7TcPL+MGIDBy2Ium2LB8zRe
lSQjV6BFax9RC4ipX0q9NWyBxFodJUR9mlun0gv0kYXxOocmvkWEnjD3g0san73nG0UP6S5jEwbY
2Hx5KjWPjn3X6i2w8paJpruoegcHD7fKiFtclKmBKXyHifeEtHbTI9lb5Ofagt7B+injqa+yC7Uk
/i71MZ+ptUV7FypOv4wZ7d17X0KxqbHBKKU/t7ykIW5hEpBZy9XM6FDIMQOzWbCFE+zEJHcx2HIk
qjiR+WbFlxt3DIHziGLhYcN0nlI3X7b8hd5vYgQK1KSgCiR7e7mu1h361P795OmLcc73S/FO9oSb
J6AsmGMEAu9R8hQqWMZURfBuyoD68Nas17t3KUEpoyGdavqlQ0+m6hqbX6p9CZ9+bY1zFzLRjXma
v3diJ5o15DHgO7TW9FWVcD+Ml8tG/YGsE5u1lYdajOq9Mk47pI7kzT17vHl0RfkW35wu7/pQKk8/
4TjkVrvJ1SCyRE7Pcg2oDnf0jY+Xs6xhXQooaGqk9bgicudjYCbp1sefSUUWVk4B4dCObuQnqBLn
kCLqc4ve65kYMegPWXfgRt6/a0v1f5BofEr3LG01irhe3mjmRFK0wIGOd5pcg2EZUK/6PgTWptw4
3VontIHiXIEKsPIBZ6dcA+L6CM5lqvPOvBTXT+GEEiybGYjC7X44m6py1dWs9dRc2RjUiFX/p9jW
aRKzwHehZrdNW8RNKtRvG0G+MGabTqcytoQR69TAN/WyIJaX/zRTV8ap9AahVF8SCKGI8wjk/2QI
bcz3kUdGvmxC8shIU0N0ycmGr5tBFXd0OhfCJi3/MtFlcRlNewc2LUXefOgFNLKxZ0KniN+lzBGj
Kmfeuyzm5kExvr7cy4bn6ZaMuDvfRPGKLjefMk7hVa8OSzsTXJTNRoKXkhaCNQfHGHBjrOd5EE8n
JBy9Lm4XNVHeGjwY/kWMHWIEcm6SpyKD10VG8TcMU9ptpB2G92Egdy40zqSbFLpEzmKsDuNT9BE8
Ba00iYhrdPQbUipB7Mr/B/mqmr/OXZRyd6C+DPxHLp+g/6rqEHudm4Xx0avGQEb07685fu3GDKUz
hgmTxoDeQNWGRzg0hBSFHUsCWr2B3fTPf3qSuahC9kHp6CDDQFdL6WsXk/qH+phgNBAY0QgqfhzL
fuJwss7AX74aWvYEVQbao4IqhAAnO3xwahiwWg6F647s063waRx/iFYWZOFcxDuo108ssnwF6w1c
yO5JD5suZsMNEBO87hx88k2nvLBYzhQdpFI//rHsWCzLM9b0q9Offfqwj/dHfEiul0yO/5h12mNe
VVHk0EJO2qtVBBI+F0X7LwSi68R0WCstS4KajK0Mo/q2gJTdJTuZn6zVYk+5l6MIZO5CcWCfhLAz
23AsMD6nWF07BzqBC2xcMR5wa4hFaU6EMCGcRs4QX0U6WEcwZuHPFbKh4tSALEv3EMMCbPkgud6m
wUCrG2DQEldPlHQFXsbi/LYCc8KOZJUEWjrJxpdYoZOYaY13rjND8LGvud14mt9/u9RxmvvlU81P
BoavcEPEuK6Hy9NdQnOfhjoyQOLOZjii78h3srkbePG6hkwkVY2/DpVvCrZ/jf436ySb4igRgPz9
HxC9JXr7VAXpRYmd/7BwUFBp3xpVxNDC9br+QVgWW6Z/FDN7g1mAEoxWF4+/Em/1Hb0uq7nHFQzA
SgGdQRVMMfTkwC4rU7UefaT3WZffv+Ezilln3jruW1Wig+uN5W3yQZnbykwVy+kTSlVKkTe2FIil
7+hMYGnMOT+mq2iqpLA+wOIltEj+rgviY7CygNlRrk/sk7ECFF8I7iMVg20Tcpqh3r/MmrfDgwBc
GTh2zKVB+nba+GgOSnJx/HVinwBnUUgbN+i5urTDWHsr1iIDPiRuMb+lvzl4itxVyV+E5donVVvW
MxnpvaZMR84E61ZXyDIHDw9RrtziQaYnbvvzfFhQnKr5t38xKqXbI/aAaf5lMfmVNZfDliFTIjLz
miEwlav0A9liOCydypM8aqDGvcX8cpz21Okl/WIguk01VJeqr+6V1JQjZT8piUwCT4/cfx0LSBUo
e1CXQ51yKOZo23qKV1C8v/5YhNulOZoft9lGbqgVuck3z8QP0QOb10pyvoveb+As5bWkcabJ8zYO
D70zEGRgWsTUahicHSQKHcT2OWhhFaZwkwPqJrH4wnjAF0Xr12HTKo1yJd8Eqw2hyWIG/RrLOsKh
pDknFulcHzCXqbgEjbfB+Ng8RJesiBl2oXWpnMYTHDBumsiFad7y2DcsbKNQvdjBZESiVZEmcqM2
+Y4D65ZeKg4d4ZpOAccfEg5RGUn5YKhWWWGEc1rcLrGUHJqz3s7holMM2RbwDQpLFROOnYFI+m+6
1SbrltbHRrQG55Zlt85WvsoFKa7yCtLVhxVYgNJuCoSxhYvykas80mAFhJLsDy5rm6GFTDIxs5Yn
jEVgmBzfQBcfU4db6eq+jypUJrnWgZH/mMP3ybdN0fHhL6u7kztcDonARbZBwnn13NiXvymxE3wB
/N8EJATC32kLKtLlcfl25Wvqa09grZIRxm5RKkxC0s78qboVmJ24OmPd3sstTtkTeniCiJC2Q9dc
wr6PhyL9GX+zdvAkaAcgHmbS/NCMHRV9FI0jRXVNezMzl+tLu8JVs9QHDTUrsOwzUJU0v0kS1/IV
nDBaIriyLr05dgTna1ZlggJytt4kALHDWHwTek3gOVLKGCKoaYk8ROreXyUletXmNvypEL9dAvOs
32ajEBatzpJxe5hTT8QSDyT906EUZTUwn7lrFfkvsBmgbdNRP4tC12S5P1aOqYh3/U+hRUF3N0aL
KzbMwROFTrLCdZqj7Qu5ROspHcOJcVQrPSyrNYwwhjH6le2lHjTFmcu2PoRUg3XC3pcgSXnxEZ2I
F8uNRtzgSrS7ivYYAulHAtwJTNWHbQNOGrgSj1/CFA2QENLGQm7zoBnCYbAzkkz3XNFf1FTfNggv
wJkpuCh4s7u+8cpZ/qh7JPoC3dO1shF7yEUuCX/x7Z9Zq42Bwi4dJMJx+hALA9nyE2D8AFsrTj7Y
kovHeSZ8PpmqIIuxxUpTRcHesu+HSA4VI0EIOGlnL3eZJSx9T5T6gswX9h9spw8pfWeAS9KgZaeL
wCKFR88eRj5cv5YPgec/nMm9Dq7psEocd8C7AoWO3tdu45M/d5GAHmkYW6+6I8cXJTE0CdHna9rb
HX/qQJ5iBtBFehwiXvPOvPt7z7m6gMsYySnIQ1yEz5wsQryX32uLwktFDnydEd1KOdMJN3feb0KX
lOUN3vi22KUfAX1BHdlXL+pqRV+MlV/c4PXrzIRhKOLkDK5m42o7wnL3M4yXQnUvHDvDXzwQISFp
bGkqvZga5QNAUTHMoqxqvBAmhGB3NjXZJaLERhxA39d4F55scJUraqDoGoA10rmZVr8W3Ed7FYFt
19tVy/g9hgdUd5QoFz8TT3vNHJFmALOmS10kx2zK2xqLEFEr9RmD5p0ZXwZ9ceZWyiC3v8V4C7jm
HLBM6xTzaWfZPq2MgRp3fMJszDBADDuurGXufs2KotjD/L3StI4A6Fj8rzi21y3WiWwMWCJXVbTR
1s2teuLDl24XtE0aLuWGTwD6cpHsSAOdhVQ7gcZXEWK367/wUAGB1mcpmFL4qENVdF/S71raBFan
0ECiDdYUmEUjtFcn8clpeHoeZMskBjK51fZdDNgvWN0uhllNTvtF1Tbsjc8LGeDstMrrPjZz4RIq
uAyJw8E9y6cio53i0BHD4GIOvGc4alc+oROsrUrT9s3R3uexXsLSFJTroxX2vgOyP3GaPFe4w1dS
MGLkypbaEHJUQCjPHziSvpl7DtZeIA0MQoyiaLnjvllYwS/WtAzE5670q8cGigG0R+MSqNJwbtK9
up2zdw0lQJ3e1xyVTAiwSP1its/4Ltn9YxzbtyjJhFbKchoz9SALj3DoVShSeuKU4AKGOjw/KybL
zKls97suhpXZEJxCYz9tC6Yqefa4WZ9LN9JGs8sZSY0kZyVEkrPVeHwlp6knnBZfbANKwwA+YGHE
l6MVWbqpSbNrcinmZb/LC8IN3ulwEok3aEwSofKaC6B9mvXRaCbygICx08b70lrIQMqNUSXUXqza
MR/0d/KJce1EVA1i8cUY+eVHkrt/1WxsZxegtl0gwcxJf3iJD1SsIipZbSn/sBPOn6p6gJc8FgKq
SuJCxfqpUQkHK+ehDyC5HKhZzebCO3N3FanWGmzRJNz+wAxXK7r6c8nDZejj7xx6xVYc95G74WiM
x2lrCCKPNqHDMdIw4I4vzxf+lrL+xRVf+5mlUqGd47E2vXFRaSWAmYr8bDhMlVeeu0A3ncV2YILm
+MlAMSIkqEJyH9rSHH3UaXhT6d9Ly6dOPssqHJSaVjpG71niyRpNGkEq3ATdghNSl+N+5jLAfy91
+4NuOPG+A6uBoS2mISKOyOjgvjGCQNTtXJ9OwXYGqYHkcUq5z5VtO0V3sXLM3vUh3e7RybPxSU7a
yFmc3zOtPyzccZCUmzEBMRIBXHCF6EIKYlsoWuszs656o8W8cDd90j4fWni0KbzU7MTMMDNZGvmH
dCKxIpAgfqWFsgT5yWnHVJOP4ysUIOSl+vtp8wlCS7mLiRD1dOgJZqYHDGK3Mnd9vQfO4rLC0bJe
qCI/Bh6KxhAKObz4igm9YlqR4iO58J6l2R+BiwOCmII2MyPvKbpJxmx+gaJy2MHru8XPQb3oINnz
UkfiBgkiZBOSJTTKTSmbjeePx/RA29X+0xJWgeKozft4TLGIPkuyBZU3xFFzdHczVVPWDbquOrat
ieAaVDGQ7qGve4ftvXkgTCFpp2BR0wQIVg2TqsYMZwpRD4afDWHuONkTVVWvdt6FaGQdKIew49ya
M+L5FQJSgpzRamJVlNDttDFYEb1+zA8eTBH1Nby4NRN4MxrH+WB+Tk2511v9ZpTa6jDcPpgloigk
USyNmwqQOiS/GiJmfzm8OGEdhMKc0Wn85dhHp7pXE9907TO4gn6QARs0dVBSwVrC6ZBErA3ZlTAv
rB6XXhMancI9mLA3/PgPMVCwaH9FJksa4CRve+KnXtniHzxH7BIQOQfNNSwOTAo04zRxgGRSggh/
tywubXusryCJcEsWuRMlJzMfPB2F46iKoCfiCAd/avhkqL+jZZc29aLQz+J70rAh4dKMu2NT5ScI
EHv4IDNpD2j6pB+rddC0BBP4scjOXA1ZhCSCyOXD+Ly8MSUcOh2vHg4tZ2TXvJA/ibMtEErzX2iJ
0OphMqslLlQKgneeXKDbZuP5IuIxVu1uJoge7MYrQ54+NwMu84MBAPyzBWekr+xWcxL/mrNSKsPf
AtHS423bUy1i/NfIHVaIxMZ10DQjfdX+WIXmVIzleUwAyX1GmWmyYO2MryfX6ZmzmFd676N3EhYd
f+xsUCJ19C9Eaq7ca15+YJE8zQL0QbgExUPmjaqnhc9nckHsLS2L9mneT5xuzaEHXovaQeQxMUzg
cWygV/V0r/fnW+HZdJk/PY/F9bQRu6yLrn/VTcQCHBliklWZD5xFbIPRg7HUrrYttXc+REs6IO0J
GAebEYBo9ePNj23BG9GDJSxEqz2Ll8sE8JT2TDSrCtzJA8fOToorU6lLYGfcoJTdtfpWz2A6I/B+
hjv8A1Osj0viQs6EU2dBB9A5uwyU5wxA+GW3cnS7hOGp5mmJjY6EkHuHLIEf06N8VEb0VsJI4kKy
s4MWefNlScbWh4F2faVhSXWtGRgyoV5HXZey2yf3EnA7kY/oAogXSeNkQM+m61LwJZUIxt1fhmH1
1xTddXqVBPeE+j4X36dKkrIIWX4NNac48KR13XNxc1tJVlJ7SaBqy7XhigIuN52qk6vrTUWHF1EK
83w6hDy3tIh4FkBOHzUYhbrIRS4u6lw7WREOMB+GLW1qIOdUaGjX89A3o4DY8z+f/bnxF1YIzPFe
fExdnC1Q03qKR//ZsyPQjVkVYmxvlUhSy3bOVHhiJNpeqwO70ax+pSpt4o9WDnz5jKAcXJecFh70
/xXMfu+1XElvDrbn6pTtn0M5x6idzlw6jf+GEZNZOw2SRYVRyCNQOUPFhtk32d2VI3E4LaGZqvyk
USgqarsPEfBtbT0ybHdZj7KhC8kNxu95L2W57SJkLPryFWRGZVdNImHaHR8lGXwgrKKr5w31+TLR
+neQSYcysj7rQI+CJSs6YGKMX7x8HC02iXdFohNQ1ggJf1xiFyJXVCfp1B/zgrnn/vXEtfIYiFrV
J1fC+D2oAWuigRajzIxflNjCLmXJed2OlW0gu49Vol8rvnrD9K7ti2e7pQihZ+Ue+a9CFu6optNU
fgOFyPWRQbgfGyGbMz+GjhoKiJLDH/WMZojnOOQAQP4MwyVMY2c7tKmQtWZ4xjPbPqWcXQc1JYn4
s2MPwE84ePsFe3bal8w4bJKuSEEGgJvPisSs8pfB91uFACl86Snl3c4UGCuEmMcvxk0OZNywFC4B
n18gE65AZnmgLZ9lAyqiMMCxwVdGaNpRGgRKeN2u4bDzKs7RRkIEsz9m8pm6GOE3Lk8gpOfu+jvZ
OxUUFE8SWPldyTni+g51XKybgA4r3NJKKgK3gfaKw6FydbuRcA7m7Mm+wMVCcrvFptXkz2Ts4PO5
wP+5TbL0rY3S0bUJ0TFpyl4q9DpQTxytBf8obGI/N72f4IBw/nwSXQmz1GojY7/4AK0dEvg4kaSn
5yJQMpK33s7zlSRZgEkQ+CODSD4pSZnb/qnVRQsWHLXtXEZ8JYjyh3IiTLJQ43yLdlliuOmMP2+2
8BDCxEkyDtU/ukfZSlAp9Us/epYhvQsgiQEUnAr/7YN9pJ7L2JxIBy2hx8VAh85WdZxKpNKzxZtO
PPvFcbRVmkTAQKxLmltS+hKdn8LiJZ3FzdkXaImibfkz5JWOL5g97s73nuJomoW5QdMow7jWCY4i
435v1U0cVWV2D399ZRPELzLGzvCF+nUkgZNFp9NS7bLecm30wP7Ebcmt1pEmC0HFnDL22hq7sv8t
TXx7eUUGYWFsxcDr/epZ4mnyAfJZJDuzC/SfWdsAs+Nx0xaA6ZVdBuEzsSXVaPfHUbwsXZb/7tT2
jVrGbmQ7eJcbajcNqjPzKBcWWyiGomXkqR129xmJSjW0FwN4+BUthk0NN+KS/PowujWNJMrM8l3G
2oLP0ViRb5rChOxwpKoE2qCW+p8OWw20SdJm2Pf5ujNagp5nOYA4rOJ9I+9cZmn357zkmLYJQeC8
LGrAltv+NElqhoxD7RDx4z5QYd33rnP1rzFR/Zn2LRmWl2rYku87zisV8pSmC+wBOBZp+I8iqmX8
c/tJUWpp4gQk3ZwJZBvWbrsYzW6vCSWBx1Mmbw7+VOBAsXkiY+f1zRpMGpWqLG1ykVljYgwJ197O
HfxZLtR5cc3Ntzu4GN/cI/IWI54x/5qIwo5qhft2RTSpfyLtQ+47nYxV10Kz7EC3oG32lZnr45Pq
+YrESyrhG3hGAVmxod92GJil8h5khWB2wRPNDHNy2RVMKG7QTYi0hCgQ3kBOcQwp4ZjCQN46YYXG
dgIrWn4Ma2TqAX7d4k7veRDous5CRmMCA/YAIHeqqrSz38+1lslKrnnLDfMjUlG91ukmNC5F71dN
3PIz9PIRM9UYMWrBn8KlkRlxZeGS/gyx1AkP8IAzFOgsaUenf9lkt1GmLZsCW6f9iiLoYgsVoDfo
mTU7oks+li2HpbGFNBRig4/k7O5kQpPcvJEvP1Ccq2ZJr/obj1i7NTiudAOYqMAkqUWDCrNiz42L
5aFiFNXNvypbwpDwYNZT3a/J7NYNSDokO1DW26jXwIaCMSL2amYMTpNTQVJCO16STAM2ruY/wOQk
hj6tBIqnM5I51LUtea5uvy6fOFGA9qFxnPole7MKYxfq9QlPl0WZvqOtas+pSwGshVOO00grMmKj
jCiny6VRDF5BdUFN15WvtVwdtf9e9YmtwtVVmsUWN3hh2/Nz0JBN185rhAfxEB4rqbaZVP5xkB1q
Guqsb5ZEUxXjgo4feTSkS/tLSM2RY+I10AHjccbr52ZUTeE/X5LJtutW5JSnLLrYLkG/EibVXMaY
orBXtYNhIrSPUvkT3C6k6fmxnY0AA/z8trB0wAXfTAMql9GEyuGqlpp6CqFBby7fK/qaJ7xmbXNW
WhIwKnlqmq4rBonXb1jVKMrr2F7qFT98hOCsriw96Wz7heFXiDsNoLzAHna5RTGc7D6ZlGCtAODi
i6NNUsy05DXSowviwDA745nNo+u7V501nkIEScCGwAY8MFJ3TybKZ22cdy8Rh+pa6Y9iSXoXyk1R
eONHpW/z/bhYe/55CtRq+zENbFse62kTtV6SO9SdOlH5h0ldq1AS9kDl8O2pavsIn1crJ2UJtuX/
mkkodRrstneLfGfo3inTtwafkQDySjVC9eeC7N0mTVCFBAtJ8cDoHDgEs98K+RA4+kdcZnBvr/BJ
cDVUEGs4DxjnP8TQOzHNc6d++VZtc46+lNa4wNInAHoUxC562ikeZynciuGjc5de5iuvTs0vyjpk
qX6p8aOseeLHtWGkxwqCaWz0V5dX050mbhlnq6b/ZY13hOdBimhys+R8s3EQJXiApANcLKKrPdsP
DpaYBG/xIk+/WZAAiVx34qeONdUpI2lB+qmUnO5cxt65LTVtMS0AvhnXtdKYUA3BTs8UuUoln2PC
aO1QuGxhypuZIEc7HHsfTnTRNuiQf4rCNHnwymhBkj7q7QykEZQ9LCZEzZ8lzkVTs90ysKm588U4
UfFb7p3uwLdxpMIrSrJ05wjmqTSYbVQI4BuTqUMOqUJ2IvPFrBKJfSFHY8GD7BXrCw81sMAsf22Y
+TmsLfxQpoY3rIUE9RZsghltryAjnzwpuP3dpaCAax2M25SAAbN0JtMQrn2Mc4P0po+i4s6Vgq6s
jUGZjYiZx2uY3Z9XlPlfEZKkiHTD+BcohK0/eaBu9O9Rbj+ERXcrnSkBRz4S1ZDr2n/8whO78t92
fkRVsZyg/IxXaJ5WnAUQni799zJFLkfAA+ebVHV6pX8klgAdXfzwKzGLg2j8fwXW7R22hk+j3unJ
YuSeC6YuH1tJLPAnx/x93T1aavAG2tKdN78w3F9RaqBFgHsM/PbSdpn4VA0cunnY+SLlsL6Ha/Sb
zUWcMF7coSddyjs93mFkW5K4tYLaTk3YaRkHFZIY1rvGnEOwh8h506EDN6khnkC1U44hK3iUeBS4
dUC3Jcv6lixK1iraBT3Femr74PCZYv/cdJTtNYDTXhyUJsso1s1th5/MbE43T351E48U6CiPE8R6
Uhocd6p4ey8ZXDXL6FnidPKl3K9a21iuo9BwTajVh9+CImTnpAB8LMIS6nXMrTfjowWgh7hCdSC7
FBbnbq7ipdsEOXEh2TmpxF6DPswitLs8klKB9DxvHBFxFZJGWVYeLdqB9cxv6TA56fb2w1STMDWM
xPatIQyP2ltDvpueVQzoXA3NOEo+X8rYlotObIQLEeTPQPvytw8I0dnjwijj6dqNzz+Quayh8um3
6Vw6OiraURxzLMij8whK325DtA7A8pu7dr31fbQN9/LOOAxgY6DUGWYo0D2OV5ee7ym06s9h2hJ6
ycE0JB67/5d7w8+oTUB6txAofek9FMKFvK+E3/H2BqVrOvBXY1VnAkwGgjHiWQ3chUll1b3ByZQp
F8R6h1rbKQQzjA68DwBK1mEi2RirniH6yWFt3Pc3YVYZLrFpl2rfnEqQ1/J00MTH9QNh7L0GGMYf
Lq/LeQ6cQpY0WsQm/g8tgNlvhXmevrfyU//Du+/fYyqwOwFafyfhBhehzJ352QoLw6DPenuNSaMM
6wpw5F9YuDJ6PekNtAFDjFWhe9KiwtBIAr9OhFenXiR5IBdckiv8PST6+gEnt2yQBtDxiCiYHUcl
5KjimHD7UtlNEzP3hUdbI89PdapG8uItXmLEID/WkIK+TVGbSt/S2Uywb/XDf0CPrKI82uHHSLIr
0Hz0tT9CIsZeozS8H5QoWbOqpssccPLpgb8uY6+8Dqo9nh+4tUTNXjhmJdFq6qHqfyZYFHhBKyG6
ZqFVp7r0rySv3xKG14fmbfcWZerYV0dG47U/4PNTTo4ZqUwy5f9AUeibdIjWOpEehYtvXJy6VQGF
AgOd8rQt212nvrotk33ovSc7B1LOLO7h6aBRrOyOeCBkLA4sPts6n6zX5lZF2c9GsS+6n6fXMUH9
Yk3MSLmJgjC/yj8bGYYPqTa9owPuI56ID9aE8FU7iRsxiHT4OniQPrsaaqaRX3LhGzeMHduB9kV3
/64U0rq57jx8ln9idrDOj+fm9v9Eu92C7RSid3NOLqQbVoyBhDOoXuLh2YyWpH3CCaUPMjx0ii9P
4hvcL39moeeifX3YdWA0TBAeG3Foohi4kulr1JDKqbynHSrPpj9L3tgRf4ml0zg8za2WvsJZ9l1O
PPAYGnsDLQrl7GR6lP1cijsgb3Le69+w2UYQWhkLUBAZQ89ur9LOHgtA/eIXToXsqqHJeQEwKNdr
W/L38JMTQRvAFKrB8e6XKjHBI8BuP15RiOEriJAvuHFMk/+hvJTxSG05tQGm70qbuHIH9RMarEUi
RTUCK7kubmPpdltDLEUcLyACFXfIA1zSuf2fIjk518VOWdGVZxmfSf19kS2OpMZMXehN/06fjzLu
nW8TN2/v2d9O14e0hhBW9tD/L2R9LyMjQU13fWCTMmj4MsFXWY00hzIUD/OyNTRwlmY1cYmMyXTP
/90HHTYaxeY0tIHfZhZF6t6M//c/fFCM7jAyrw5A5gDHVl2gKh2JLTOLX0Hzoq4r/WL469fbmQb8
Ue+5XAeKdjeeD8KoG24uiS/0BWBSfpMt+CscFcOZk05tiLAJHKP7u4+wREavlRqoIn6XJziEjfFY
nIMeoaZ4KYy4uECCJQpJcdGNLoFSqlyFjvIIvYKhA31ixENyU1qO+SzARMIYGZj3MExfJIsfAsdm
LbcDjZRK3UhgdHoYHaYfO51b5JL8xqDLLlean1GSGCTBKC3IxqFSi2h1zmFUgW93QqF1K0fCLdXR
o6vt7xjOyerMhbMOjFFLz2h5ms5YEoxjHQcMEPHnBDOu9hCsaKe+01NoF9EyosKWT/9lBGN+CL0l
8Uz7Ddy+a0JghMwPiq1ThS2M4bGfnOeBPH7Yn/KK+HQ8LgujVtztTumj0aXGFfQg5gK9N2iAhq9C
mg4qhZ61bTyjwCaxegrnDunUPMU8qHfQ0UvRyaKjAZjtInVrXSTZDwdpAHGXOj7kwve/vb81nJVF
EKDx1rcTG/sOuTEe90A69sqwo4ybKmryO16ZNX3BLgLnOqWmA+XdaoYVmZK4JENpn9jU0HMbBZ2+
jKRuhkWaEmDh70260NAQjxjR3hJ06VdD2ObIKD0DY3o6CkyTUBh1+6H7ER4Dnjoc7wtFkthU3JNh
5r7+odcTkdRukaNvcjNrQwHajpUQGtJAgSt+RW4t7oChFcNAOD0nkvtoUTMT9unGHxa32C6VxkYb
INHc54dwXgQu30hoEWPRrVjksHzvUNtfRF/70pz7iT7HHnXi5Oy1SSzqVa7OZtpaJ/HXRuA/gu0t
w2j+0+xpI9e7/XlbSFtxStfDefSDZwmGnbgHol7e+oQKqOOwPlFT7uYJ1uD9S941WCOLXAxqkNlS
dik0i8ZyQis822Fa8bZdeSK/L9YM15BVQIxW2BsYARvkNKJki/VBsHXzWnT2rnbfNdMsN/43aauC
PER2MKcV1aJnDLmb8JhS2MNE9Wa/4OTOBQrpCl+q8H43HezaytEkJdzvJciT0mdahtjJtDq1vEpN
iHpXhoIG1/St6LzihJFpV4aUnTKFrIb6KLztTwagXLX6KeBXJIhBUVho+tleHgE+JheDmnYZr3bD
arlNGzMXBmaxYCJVW7NxdzXKhjeGzfThAwYPjA6WBwWFOHHZqYEsJi26NsGIiQ6Zn65eP+bjvJDO
i9pd3nDDce3YwFl/QCjjeHv7cqJ6AfvU/AZA7+TdQL3XGHphHWAlofw5EyCYAy4PwXd074E94qYk
sl13/9mbEw3MgFYl+6Y5u+Fcv3z7fuIOWZNaGT+a445oVhvBHIcEzGexpqfu/PVN+JEdzXlvo105
Nkrm+H2qN4FPj3pVBsFau/u0b+NKBREKEsCweNRWE0ORlc1/33GTah4FGNYn89swx0tKQE62JyNc
7fa3JZNT799FuxxusIbD9BWiqIPTIxtM82UNMJqsTmEooU8beec1Ep3SclswNh9fe2cTwfSV/lqP
hlSib9cUMXSX1lRuur4dO3979uW49rPDhY+dXECnBhSe+0u+JmndZXDt4NZx8ePd+7bBdSAGQU1o
A/SnVr6t/U/tnMnNe/lUYHGX5icXPi8/9pzzdSa7V/ojxjyBb6gBpdo5EjRW0HuwyGlL8u4HAm75
8/YkCFPCtA+/tydUw27WpYKaw/6/AmbdlXa+mguhIO98g2pecu6c5tgV/Q+rgoKtWZk78a6HXs29
tKpBuTmtAp9aYlL1noasG+Ro7pjMOnZLU1UsJqOd6s/9p82KWn2xBsEp5yrfzczDFlN8LSQdk6Bf
UX91mSuRtRmVPDe+x+TFek3LlnelvCY6T8i9DUiEvt067o803H4W7zSAJKcaZoedFIzfzD1wrZaO
PMROurAq7V6Ul4JIZMVtowpjs/qEzYtmY1EtLV8LzJ8f8/+GXmuCWdsw1eqeBWEwMVLfx5FDyqTU
dUv6v1GfNydPANPWLnSOVV2Q65IEkfIVQaSStYicHU/NBSJreagcXD8cRYbM1CjpX/zxducnBAxt
Bn8X6mAq40M0BhBFiflIOj1ewPIdDF2/x6uPjmOBxecLp2Ifzd9DINJOs+GIn/+mqQKj+gDr3fBf
jzQbFMnE0JMdi8+VG7z6+eQjCq84eCj2DQeGC8WvnCvGL1lbzeXh9ND5tvfRtiNdwRJBRt+HvJgK
J8yzkIx1aFGlBJmD7+lxYemqo4+uOi+Ew+TQW5+AJMZjtfDV2gduzQOto013/3iDV1RffbIUHnc8
TKgfSKvSdN5ZWU1WFebO2sKIj3noImC9ZrmJtksnu76qY+a2tjll4cTKw5OdUYA7mSV/GajD1lij
ZqJIAjnnzZE5qB3uerJYX17WCVP8dkrooM/N7/rkDPyqs8cdqHv6OmwjOEqEUN+n9FF9EdDb4FbC
xKzOIAw5B8QTJ8x5eQbg3iCUCeMT0bTQIdDwcs5oO3KCyw40GcMpXomwjgqDrCbrR2nj33qjHRpI
CIJE12OEayfWKJKoPq0VSstB3IYx3A/yNZsz292BSG/JHvvNBOanLvOtlvgDMXwF4uvOlqeS0eHy
7kVVcARKWQ0I+PZ4eZ0vFRGvtq9Yj/Dsx/LH/GfMr/A+JQVKBajSu9O2H42mNd1OxSSvesY4XCaG
ls22IoYzi94g1wdaIPcqyxr06Ji5LFyPVjlofa9Ivkk9HnWcHaBlfNjIkfIzBjtjT0vXQ2AyLI9n
/oubGvZEeghywhp2H23nAq4WQj3WiuVz6MhH+5fv+9DB7VfsN+a2wil3b14kMhA/uAiUeP4yvGNo
1M8GErD1VU1eFS7WUbJP4BvwkYRlsQ4L2xUzyq6YPq5RnDjd0re0VrG1xCuYtv7rZemy5HLRnrLV
B3/DOgO4NCF9DlFcH4Nu2tsRzbB0Bu+iflwEYp35W8g+N4MrnnGmCgHMRoEChnYgcY3G5CzwGJ+0
QpA5TVAMzZWf9c3plZfqfixiNPN8NM6SagQdxVDqoogRGD6/YZNND4Q7yKvS9VRzdQf1kiT/IpBN
tsHYfqHaWjDndp32abp54qTQmgzO5ECGVGdh64XSGMW66cVXRVUHISlRO6v5MS3cenTSPjRIgS4W
+iFAoBKzuCdFvxFjdI6Fa+78oEy+sTx8tB93wxH9dncg3QOEqsd63kYquCo+IBMJPWAKqEOZRiwx
q1s47FMVAnOT2C8KRXRk6nFhP6qFya2wZmrF9vuyug6aQ1Wk7yz8zqUtLa/DO+lV3imHS0hXSu3+
oRzDYA8N98zl0Y68e5R1NE8tRBlkLqes0WydMOObGJUQjSAi+2aCNvJK+wanS/kAXW37nlzxZXFR
E1Xa2WtiHYqUWjhY2Dzs/RmcoJcc4lu4dXCHyYfh0my/l5HtG70i6jx8Eilek+CQm3/Kh6SjKHc4
YzigN3C008ZLFLe4M/EXpz28093BcEYBobLAxYS5G2JSwRIfPlJWJnRraRajEK9fJSw2MvC8SUpF
9VYIYALc32Foqevv7gYjHhpEQxnCzhU3ohhA/F+mnoV5xhds4RMgh/yUVStGpgu881J5F1vQXncJ
bki02yprfATdOVf7vaidFPyNxJSCFlgT3bcL/Mwm2UT/gfrmSMe6w+JYZeljJtse+m2qjN37B/+G
KPraqVD8s+bxlTWozI1zI3DCMwRKzU4XT+HdhUA/mS7WSXFi6RmsZ/DO0UJ+FTvDe4WSUfxVWDsp
bNNSL6sPEPzcsRYUN0BGgm2m76D/YXqU2Emte32MojjLlwMUOLSm2ZbwZ9QL/yLLFkN1/0x+U91K
p1rlvRNoYI0OZxbltjJijhYSIwABN0JJrf6+sNqlF/OL1pqVwveY3X/0wcWqZD4dhhCsveVch3PL
uUgQ7eHSqh17Yv7ny3cZKOu7mZEo2YyvBRsysvL4K2XRl6Gdg7dBnl/Q4MXt3Iqqx8nd5yrAzAeF
HVDzG5c6HMCUhzUUOV6LJ21H+ITO+0QAizLdGsWZZc2RIL6H4JC63tD7Bqk0HGIwXTqu/vYK1Tq5
m37cTTJq1uy0sa0DsMr1rHeiIubOffbcSSHbgGKCluKZnZIjD4N1k81SB/cAvdtPDHTNwMhaB2Ez
cCdMIHnBrjyirdMByPYR45hYk8tfT2PxYavBlzHjUaprZsBoLcRjIvPwoOMe/h4N24Ceu/qrnHbf
hyFTphUr9xzh757JLExFB/oL3p9CwMjlWhzCyL3d8mBPHlr2LAFvjdAFESf1vsXq34FlzhlXTK9d
DcAL73ibanD9tO4WnUjJf2MOkyFPM7cbIQ/b9sG+yi13qsmm9sK3RF/Nccv8HI3weHCEtWTKbQ/B
qDTRbaO5SpOGoFsqm6sU2KSeSYWfwAYOVArYLgybVdBXAM938iGNpAHposN2gUFS2pUNwMcQdK3S
cSFA+tpNCWM6WThtVGhPPz5ANhJNeOeOqxEw149DjcvmtmNUUcJVvFyuDR124+cMjrsjeH5FF9Jp
uBq3/+iKu+2BUApB01XOwSLi+pBPMqSvYdx0mPP45ORjDSPZtbheDqedZJ3DxBKuXKKKrYV20R9s
8EGfwNNIdXxQwowxLbXHD1yV3+wDUQugGOpNR09SQa14co130lmCE0tqGDmVwmEhoXR9bH0Ewahl
H0cpzhfwvEHyEIZLdl0E8L3p/eUA9wQYDfCd7p4O8wrYKZLYDi4pjgAQNGOvZL9K2RjmzeXWzf1I
wuGO1rAG7uclwEGdfE3GL8PQO7CKF4DiQDHrXzebKlL2rdxEygbSh6sC32Xpi5Ko4GufwCtgbmWv
grmbP8NPUGM26dhB7k3TdR1WCd35pnc8Xlb7AA9Er7VqfsuTRf37CQ11rt78gE1E6zfI7sp5xwVN
5mLy24hMdoBYPmY/Z5lvClZJnZZmqtffvGPahRYEa8jH7/TXcYWMmWVr+O6/IIEzZDjO8MAgSEzp
ZD4bSIkemkxXI2Y0FxhQnU8Jb2ZTsr0FaiSBWJvS7CGMDYLqX1fte1JMKGLJ7FugEuGI7PA+oTOe
+2qbIqCYtfCt/JUa/g04ARxuoqNVrUNI6MBiUmMrFqQ1WdS+rkkTlYR3MTuVwtolO4Q3FqeND44p
qOqD3TBmwPfR4Rqg5C0Kh96WkrUiM/nBntdIrvChAqoqkiPD1g2/YqUpWwyKSOuI/OKxYc/e1YNQ
q7ZXhu39qGTeIbzjBYiOoMYiyUdO4/23hbTACdRreR7Fc4bfQf/0zZiCj4SPzuZdqhjkAkllo017
ywDdoFnXWyui17JWTamyJCZenaN3uFem4z18t/Yk40yM5B4gGV5Dhu1TtRnyicHXSgg89ed6XSws
Kh7GUpjomlrn+eyvlgocdL15ZTJSexXVNhdsohM9kxv0T94P3C9mzWT9xD1oUJuyBcudXg/Q4X+o
BCP5K1oN29r2L8qLs68coyzgkjBZBqiHj4eIy8PeDM/9P+KMuYDlPqBpvpEf0qbFetPLa+FgKJPQ
kwfXaUL4gxKu21zkIhXUNRGWhVXiNMUnnSjweDJ4/dBIkj6Bgnfl+HOMNDxREA3D2wpSiZhhsb/h
ETZstI2pRaWFaqRQ4hzI7eaEmeb+0EBci4Ovv3O/InhJjwrc3oEGkJxpRX2541fMDkVSunDG3H+x
v8WwbK9iGVbPZurjWBxX55X5zZrVtbRGkB6Em6JqyxyCQt7XJHbST9dJrXxIhjvMQbPho+EvaQMY
F+ezm1fTcQwfRP04Q0xTfiuE8H6SjR3e0t6eCg16sxgUZyXlIu1Mx91NtRCLQ74s0E1QCW6P2rNI
qbNQfhenftogVtu8l52yGV2zuausIudEbiRkYEO/ZR3G0Drcc1fwtNyXzbUAc+RN++J6+wuXHMzU
3ER37mMxq9zzpjf8Sog2sF177VTk4I2EJ3i2gGMT9vZ6XUSkqTS6OMZLLHEtVAU2pWC2h+nggwit
bY3S76LAWUXkE9cit7tJGvQHrE4ntYr9Bri2lzO/A/ihwx1Z7uxm5WeVgnjooaxt6oWvlvzai9Bn
7300fbpUfKe2laksOxfv+2T+jFUGrJogDVVPbyx2N+OStBe5klq56a2e+stV8fbmgC5N6Odfqx/Z
H/bqBh/zVI11J2+thL3suntVDEaR4MeqI3herS8ROKa4cRiSnXLT97Iz/feh+vc8JLhENWgBWLqg
sL/DJxkgvQW6Ld5Zn/OwgYAtWUTOIpIwpCeJAZrj8P0ebAx0KRSLrzpjODbU6AS1GKJ72R+DREyc
Qg/JaWOiM3xKtVsTP6/FpqBJ1P61C3fCsmWClPhFY2+wnsqfCB5oj5A3i3Bt6wNxGnkPfOP/B4+t
9TlFT1gcxFltbqAVfOWyj/aZYf9fodr44EvlyghrrVDv6QFjrxIYtCvCnmrYVP6rFxURAJIyTFjg
5a48wjpNSTXci1ny4kPks0KKx+E48SVap/jT3MbA/DNxAofUodsh0l+D/ASZ2b/5DRNtqyOELp8H
AhgdkT/EKOt/ickciWVKvWp4WQ9keKlCSV31grb5ytalTxK/xFsSzhQj4HwJKCC0GQazwql13XhB
NmyXgXxwbBVcjaw0sCgzeH9vwbr+1JXX5cvaTVAU0Hk9XfRupvMghxH3jr7fIH3enTokAyHE/XBq
A0ugCHyQWnGhYgIhBD7loGobPIuzHVjNtkQoPFWssCi2RTf/w7Hzbx5csFkNcWpyHxpm88vU7H9+
AHahMHHeemHwM+PeDIwS57X1KxTaLAW1mqqt+9BrZ1ml137PC04rmKoDhj/QkQ04nbwJEVT71tLv
xyWDg0EkXyD5IRT9+G2ebK+V5fOY2smEA9CIeWlRemj+n3cq8jqP9VqCsI6gHsrnfpnF5r95i2cJ
BspWNJoYRzuLdLGh85xIX5+3o4FcKeFECq7+v/qu9LOBS0O7IL71/4V2VuzebLXQc0W6QXA3gj4N
n0MZnSQkdecBdCy1s05ykm5UJQA3ThAS7N22e2f/aANhjqzylKnKvO4Mj08o7x9D4WbBE9Ky0fuZ
klAxQyuYZ7FuQGMkZmAvtYCaSBcBa1vnrbSoEctCza4C0omkCxVbZ1uLQs1jDIoZ6s12jJXhvmWM
X60q18F5leaCZ6XWpJa12s+6fU3zo9PlqTW/HNhGe/aNDPlzmqtSG+BkX0XKpnOgiTrzKMdfHDKd
TEYbRj8W2o70FSFNw+lXKGU8PMBkPH/51wcxF0jIpNoGGeBTZ7W/AvpB+81VIfrE/p5ZHDRhWP77
3Zkm3DCe9X9EYJvR0veSvG53KY5x9E30xAIKUXi9H57XDFdsFoh1cmK4+Cei6LWhkoenTXeJiuAM
Aj13PKa0eFFfUjzvWB85klTtBT8ou4uBSyVb4Wq+VxH1IdAORyKPI+t4aEsjqC+p0gn9U6GTp+zn
yxwLockZDj73Z+S8ou1+Fm1OLJorL8LZ4j24pgY8F/bxJR4yP45PT0k2b0QjqN6Lk7f+MI1LKWxB
Ar5Wnue/C5InGHptV8i3WfNxADM6TDd6bgvCKttemqo/HIUPbB4VQXD0F6KUvw7ub37amFaets5s
P5kFav0gTy8t9GSni2QK/YGMnch98ck+2Vm8k63E+JoTuwcVOFOnr9dr4DeTYhobmh/9DznikSul
PWOj6jPveBaAS+fmBV0CV/diPWpz20vL9lQRnwyKMIXq+4lcEmUqpSCGpUU2l6RInUsFwDttMBV5
XXn1ZjJwwJserTzn5zd1qANp0SQSYgReU+iuuU/S607msoKrLZc2it3uNNI5g686c5Ok89Dj5kXV
HGkgKPy3ARJpbUKxXlmZCHvu9TPQ0XQaL8tGC9IescxDEECN5JQ7iuQSVWtKonbeg4e1CC934u85
5y7cJ8ku6h/uE5cy9Q0I488L1d0oHq0ZXpCUs1I15lux9UC9FzhOSnq7FaZJw046fpeynike+xqf
gBau8UmwsYwwgawmqN1HkmH24tAlXJwm87tvlY5i5QknQdl3B4+S9UT7+j9EjC1XYwZ1xLjRdQQW
P9dhl11GKdXD5xk+f1HYzV6ndYeMhj2geNvGZRSe2iQCwuCe50JObXkwj3yeGOrnbTgYXKKBn+54
ebjuwYOF5tRrAaVObxIsh6K/vsrNTlzrAyvMLXyvNaMhck/K2tuzdaw53EPHYuc2HoNZWeGJFA6a
arRPowPIFm7/2vlai7gRTCK5ATbxudzcogv7z6RDRWu4yfFFxGiCbEHcuQpt842QmDobpP48H2Gq
8V8J+rceKNbmqgRRWMykLAlnM1V2cl3tN9YkN2tUNxLjO6y60MswR/X0ERlGMLuhUrfcF9HvZyd+
Dylpq6TCQOd7L4URyxgg0Z8nUA+Sigubb02QpVq5TgAN/u5m9BePD2CByG0bOn71wwnjQ++81WcZ
5Iv9dXdlsF7jvzuz+RnN4I0FXAiSg+tADzYzwm6OLn0tLZ5MfC71bZ8s91gbCFEcOGdHRJrxmrgi
gRsYhVsfyulWsobVpVouZUdnhWQhRH4k8NaxAn30S41kRYtIJ7sCDh/ZCyMxug5ezcqhqGYWV57B
xzKjs6EgHK72WCrYbBLwCqoc52zczpMH3J6NVSgmPvGLFvDJJ3fF8diDbM0E0NXyBradQnmjJrMY
nqDyjm0QUlUduwsNc8iatFsKix6f9L8l+31bgXmpxsQoL1qYAcz30Q9S2jwcipdhqg4/aQVtTShB
zArTex69S6IW0cSTn04fX7zNKLZEJEvpEWSoa94rcIEQTfJp/T32yKv0MRmPCqUBs1kjZzhdSGmA
fB3WbUNR/FVCFghLSj9Z0y2o3GpS5pWVfdhjw+k/0gAA0XPjGbM3mFV9eoi27ivwpzdQ7+tUlokC
kWljjkAJt+jIbcJoJgUs+mMoFzDzV+ZCHFvRKI9NVhCe5j9wr6yOvcd+qBuXrFjFg7AiSVVub0CS
XbRQ3kXzRZP/wS6cgsfyp2g4TkaO3NOZPpAWRCGe9MpRP/JaWLkZpIcdY84OV/78Q+Ook+d1+l6V
nSsveQFhQRf2YKV4CPteZtLc1i2HecMJRHYPLTAkEQWJ5m2di6/1yvH6EWVc7/nYDlYY3Od5Rrx1
Z7H+kSDA1pTxnIc016MjFXBkk5F9owgGUVZ5D8jvDLrBgpK1Oajs9HW21zLfTr8uk9s3wY9jlD9Y
QbIcQdItFs+07FEnZcLAQtNYtAzaB86G1YsMQpGIRZrtm7R6RQ7XX3lYAgSWiWQEA1ioAG8iWSMR
ZAToeOCgyFl6eWbbukH8W6oUxZm39j0FeHNerq/tM++nYLiIhtBTr1jXvMprME+Jy7ukeOF5S2IG
yNs8CskvBoovbod7y3uvhYeUfnDj4RuIjn7P4cYJwze4jkHb/u0frU10yDpiv3YInv5JKqQqPnKF
TiN5sMGneCMBiYndWhtUfj/fcVOSbINZvfCwE+bAEKm+FuKPwh82wKwqUxchv+NaHxAiMLXE1XyO
1t7BHZicgbtgitUrDWxKY41dKei8PhY4v4rGfXwYpUpCHgMUBhqgA7YYBasknYPSoqAcVbMPMzTg
FK/EJgmafaWQwXTnaR+3Zz2JC3En8AlNGLMx5ruqcgxcQjGAp8dKTlPQZIQAHbZszZknAt//pR+G
DoFcUgGF25zNErzWI9s+Tf61WaT8ufY9+UdyYAGKm0Euz/gkGE3lzWPR7/50u5+6YYzBfTKi/B9k
hQNEkuVhR1TyIKXhc3RuGlffIC0L5NTOdRkHQrIKB7oxLFBXhAOQpnttXwZwOUrHXfOkup6hIedH
2q02AdiycrmjU9POgKgs/wbE4lsao+NnvPqNMWC2+cYmlYiT0K0E5VWzmUp6vAe293LafpABneS5
zSwxKpSw+O7AAUb3LltMnbIExY9jFW4zhuc9xMegtGIbnCwhRInPE6lObitzwWzWe0Qse1Z4X94W
UgJGcyz7iKSzcwVSTWXnP/pstEb5UEKEg017RwL4XywztjzEUZP5rhed/TxeFyukT/VXkOwdWzYQ
qUwE8A2UOrhQZbFXuLPWFXZB1MW5bZIMcDSEmOT+KpCndJY5TooXasTBeZKAJOSfhkLRJSNZuWTm
w65BW7hCn0Z/mBYJxqeLdz4Xt2iOFyqrQQC1cQVyBxGIGdJRxbfheWrRT3ESp4gUhiBL+WgRijCG
6hSGbLWt/7xNdxqzyqJ/FXuzE4a3/RAIsXHkPp2mZNKNYikU21MqHFokmLOFRKNHzF7ysoE66uKf
H93YNK1b6dpdSX/yNcn3vWSphfve3NEuc5BhUNh4MPnDueo4nDxRx+QvOpoc6Ci9Q4VLKYR6AJ1v
r2mr+VKgu1VduI2ZMZn0iaLc9Zf9GWgByW8xfg8EUaF3XWZoHEnRpTapyRKUQrvD0SENMitcdbBw
38hKxfCNWwm5TZ1M7mebmaqwpg9nw+Uhx/xjr0eNt9QeggVnM6Qn9kxkxJQFYTemsAJpx4r9ykMm
j8KYwZHjD/Fnjr3xOZ9NURtmWA6dopaTN71nfJFCLh84q7GbVFf+qqaJf2gzi5Knoibfxv6nrL7s
CA/O6CxCfwGhMWtwxnMT6lLeKez/XsM3eFG972uAoLXH7FfnDz8Md/GaAHnlOFOTsWD63bxH+Fc+
lw1CD/DJUCVJFNkHMTNusbVdgFIa9bjugRHTTy9KabzAnsefzh1kvD+pnhyYLagCY5xi7JRbGRzW
3/fjDATm+GxXQ2oPjPNYZRQ5Us1J62YfLcdeSW1PheMTmJ6XDPKBZMOvrDsjzcgmN/qgsG1Pc86/
bZVFgiw+C+s3dlsAtstUuOxmbvUc57tJ4E6mWv3Xrk9dGPeTXXGtqg4zrjCjjPPKNxPomgp1AI3f
VJycpAT7GhhkzYPTZ1Nar4R9lqLvJogv0IoLxHX+BDN7Y7vp8RLsxTzXS9yG2SCZhEYEdZDOSQA3
QyYK48qiaFqKrlq4lS+rQ+CvA+O1H9hHAH5XsDMQtLScsneoXDL7VbzInYctuQQFC3RXX1hH8wMm
r8uPjB9TOJT61b0WUWLKR+4mIqLEHukNaStUvPOh15y9E7LtBPMrzDA1HC/suOIZvx74S3VQYKUU
X2GtEU/O2fvkaMbSjfhAzZEB/OzzMhTonVD8TW7L/z0/ll9Oyd6SHvYxMiRYGDUD56YNNgKNph+w
vNvOc8RnPDErQrRwPogox9/xTpeTw6WSR9I34IMHtD1kM2t4J1OPmJ89Cv6gPsH39yT/FHaJ8zqs
QR6mA/X61Z3B7/qTiKM9hxhXhye+sWqoSAwUJpbNSq3QU5M+275FcIz8sUMfYsWUXAzMzEMR/RMv
uF1FczG0cqYtQmQZdwI6+RKDIhdn7rOSRgXkaPOUDizQn2ykQpMGGRrEiLTlFpVjBVzOPN3I1+QJ
93zlST2aaKunvPdai36sTM448DYZiJZNXUSku2X83dx4P1TRWpwVEy6rUaQPgrmuOZR9UXmDf90J
KwNVjpnBDEMCxF4v1nb+8CRSy3c2rLKYQHGd97UlL2D3A6hvzSLc6PkI+ZFtGu1m8SQ9S4WkTL0e
ynSfDQdC0GPdyxEf2PEw65zB1y8JrJgFbjfeI69dRVHPtpaqE/hjmqs1Pp4OzyxZOvmGFc2+C86M
IzIO5fQrs72E9LkQdVEz1ycLFYzv+cbMyDsGwiebuZDiUHS0Tae4le+cFGumkUS0v0Yjlcj1akET
rBrhrsJXXkD1iWS5VHOWa1iRPTIpqJ+OEAcj4WnCRe4aBKtXGxfmwwSsqXqI5C9NQEWWfPKF8kdd
yqvOjxIHL/hm6Ap7O5NigMvfPkA94nXCMm47iIxQT7e0BBJ6Hv4oG6YGVmSqU6k987WA5dhr9OIk
sKL8jRtc5je1K+FwoXI7m5lhqp8LbW4IojUjFP2sA0libPuOAFk4Wc8a6MDXTh66q0+uLSLEMyeK
lMjdMkhMYsXJwxW3IqTteh2o6HYaM52lB8wOhWmyx7HBeDuavzSHuY2k1lgD5yofFA4CSSCtG3m5
fOrWQNvzbibNTEAhouj3tFX/pRWcz8s7lhbjCFBZjr1PItW4jGqxtRUsgv6KAz5IK/UcEZ2+I9TF
WmlfoeNpN2q6OJpSOMV4qPJSSuaZFLPajYy/nN9p1ttaffxZ2GCan0lcnJrMCD5Jf1Cpk7pBnI0h
gP4eB8YkUxlijN4MgTOhug5spx3lMy65pFNI95ZIrCvWHm8GbT7oVtuSh3RSLiYZSefb0XIru7QZ
TgJKV3ynVmWCS1PrTwWf1zaO33leosg7zAtT00zMW1o8mUo+yJ+jcjQRztTS8DFXafmjR9X0tvdt
YDYAgxZ2EHHft2dkiXwkkR+0SFWdjTMtj5OHojwhp7m1yardSQS6i9lmrqcHfSmAUJHsCCzhbU5f
CTFiTpmfJTTOYt5vvpp+Kt5VmckOwvalWAy5pl7tB8v+BOMwJr1GPL5+BiUIGFX65XYV4fN4Ya1v
Ohbua4ChiiWwW44g1VPZFvLgv7oPnjG4jW/fIKfbHrutlmHAZj2Ql7eOrV1/ZhzSgKvnIGIZmuas
80sUCnjiATDeBl/1EjYZtl5hTeQWZig9AdgfegCNT5YQaYOX25rD218GV4z4oNWUJPgDyqXc0Wd6
iCqLgSWPrbWPbW5uN0pCSrIfBnv4qX95YX7m3ZOhY3TOl69mU/ox/IwX2NAgThmAtijgMtX5otDG
EiRhM8JguwqCdD59ucuhKrww2yfI/CsDukTDlfw9y12g4ol1L9SaLYxbh2TrmA/GP7SRwoktwjRO
AR/fzRHNJdFXihUF80YxfXk/gsZNBk9Meju4qou2V6FfUvTkE7Du6X8/TJJJ6MqwEB34f1wO0Ef9
dvOSJpMj/lUReorkxB56T8JwYaPi+geBcRzZtDP9ktDyuLiT/Wf5ggJ+TetaEIMcLsBg4oIhlgaq
oZlwh+KcpdlrPmOvgPMmPuPdE4JEABKXlb9otxe9ZQFjjrktOhbCoBtg8KVJIB1K4sNN4d9+G2A6
WrGGsDqvB2fPsX5nabFJadqAu6y0Hg4NQhYmXkAa2cB6KLHlbTa04EPe56Py4+sezEfWEPKnCImu
I96n4gHOt0g2FZjEiS9IijzZ7ZjQSa4BeEDwU2+HaXGzIwXfUpwI6mXkR7VXLYGKvQxhTPEwb4Fo
vluiFyloliFB1KvgxJWLo7AjsZnF2LJEWsMT0pShvbQCWzNb/Rns2jE4qFjStaG7rWyVv9WibVya
dEmfrjMuSAYww8R4IqL6QcYVIrORxzWU6wzMwjqHZyrpwUWoa+5j/eFBcIGVBV7VWVgqnqBXdNSp
AHJit4o1eZL8Z3HuoPBVFniW17gkFXlJykakQ80TDKMSQeMJ1kRDRaBBVOCiDsBZdI4cLsU2jQK1
PWkIzMX6cqhtC0cB5pDFGplTqxTcVI2QMXQLrDGOKMiSFLXjSI7HyWOvBFriqY82VNWA655ZXsVd
Z68T29NYcWfICQeIOq+8Nit1emcaY0oAeWpLvcsKX9s+NBVclJdPh0v0DH6SBsUKlsSanJdjemLQ
qyf2LTSkrYod8RVF7FwuXBRAW2qgBDUO+R7w7X4DoRStkfUo3kK+GzT+MxLyRRj1jeTwuTjHNpXq
PPjZ52HuOOneKDzSIqKqKeCiFjZq6eXXAM360r4SShFmMGSBs5Y8OfZTqDsJMCJBEkS8vbjnQx2K
u3hiqs0d3YxhU+CM5swFffSGxcpj6FZCt0zvscoi46TOKTAKEJpzeAW3Jl2/CrQec6N+LsJzhfVL
/dABEt8tGxdPzOZPxnKPbo+AO3PpIsA+clwzGDqWbAZsxUt+AqgSksPeQ90Bp77mH8bdGkfcZoHB
Byin+dSP4+6/9FbqfQCcCwwgSRyW8+n+oAuLeecCMEI4quXRW0rZs+lW2QjxkWOps6HcgFhnJmH1
xs+YG5lVBcJoI5DOjpls2+ft2PTQHSNv5rJhlUy/oSuuGBR4GFYPIgAOTbkjuBaw0dcRLzFZ+AaI
ieWzC+5RgVEkpWveydbqTYgge94HiI26dJrD60QNe1na+AOVvM9pe+Lpz4IMzmPLjtTcDwbdyi+J
fCEMJb+aKpo1xlVcR23nhnwUL4UxMF9wJ2Qhz2EdIdh86Mx2GhOdCWTA+Y3ewTWMoOq0wbQm93I8
P03lFAyNcm0ub0Khgxs3eIygflJ254uzn2e8E+GdmIlqpRWN16nk1PzKjn+x4kERVRRctiV89yMQ
FoMUZuyFEJXCtv8LV2N5QFOJu0WRS4DEk486BD72SW3B0/GpgrvbLgeatiDdCwCVbpmypwh4bQcH
AkbvDOptiN+xBMuKZ1urNZrfI3FskKv7tSPs5NqnVqnugCX2i7GMDNzq7U2WNuR9o7tv+Y/PipbR
/iP1E2LR/P+1mugXftG4GEyemA1v3vS86CHo30ZzjffNxZgm3vDGg5bIsstCv0IGZ8WFvKGRll3k
mSIdicbSaIPuakrCKB7iC1aiBruvJjg2bgmMdXOPDLcVoOyqzuq3264mtOmAxiIMC4sBFCt/aw9R
xyC8ZC/JnqmKkQPV63FQ4iqOVBBI0++NVXPbVEPzyJUhsKwfGuTB4TQm7ygo4T1MUX1AKd9ef7k3
kycBWyPBUmPk4NvuRd/NFngLrjfGirjTy95CrvXRHVMoNULPiznbMfLllkQqqd4XYQptE42TUjx5
0j9tzBq8DefPzrPGVOVwPFJk+2VoGZLk1oOedzhCNcJ6HOZv7XMkr/UzQTbhYcUVLxROf8g80oe0
IhvE87iP9aVfzRs2Y1ZvIQxMj7Djh6dCPpwEt0OETL0DUyEWzaO12cVCoIQ134Q3Mii0A8UCM+G3
QsaaLhiGUQ+tIk90HZzW+pgmQrWLagxfWikudt97D4YUEtzUVRERw4E5eN5oAD47a4OZbSzH6zyk
7PECLW71LJpfOUSHIqi+eDxTrC2AC0Yh8JNIoZZyJV783Vh55OVBOGJOM7n0q81hq8x0DAhMEi/d
IpdHwrH9gjzDoaKA0p7NKc2tGDo0Fuu6nNZsnaW5qj1a5Hdae6X+i/bcVDXkbm6bIPRbDmkuoxN4
l1oOQ0x9cs/5Ih5iFrEDxxk1gKURODUollXvPQbcP1sVqZmjAbMHlQbvBzwHOc7qCumIZvHahebM
WGN2ajNm33zpHs2d78JnRxm/0yumaVIOn73wbH599/sER5Px78Vfbf2KNT+XWnmGK3+5ZdGEfsG1
Ge+r68v6gk0UfEMZ+P4RjPDysi62qxCjuAbmIDs0CQLtwtg0xrj50zpieprljjkjFTLGwKOn8zaO
Pe48v8oyqq5TQuh77aUc63etRyFQkJI1m2O3Qjw5zKx0ccolQrJpp3TA71jLky7UIy+2jgMILAtS
1cE4P2D08CUrStGYpznOtAC6AbDU6NqTq5XDzVzmysYGtIMV/brho/SFSW7nvcGLMmlrWz2CBiUQ
SDDp8c8Xh/EeZbnbcxoTOwHkFYcqakh8kk1gk15turtyNHUHNf0bxTYiTL/dIQXNOBQhITlxzK2H
+utx3xHSPSYNNrKF/LQ9vgD53csQCE38Q/WM83GZyeLkNXouiqXbEsDy9q2OY1IvoNQ+SiAIVprw
ewZZ1xqfNNOKiChSFuCSoETVrQsLbbjWaX4sbnJxVsB7qLT3jF/PEFnON57nc/+T/DlP8nIG9IfY
368iY6bjeE8AhceEoSeLOh2w5nd2GeE9WgANVm3vwNDcqgxGRxnC4BJ0+mK75sNMGWiji1c9Zz+/
o4snFqAtUdZGD087/3jyUBbsMM9SbTIYtkpae8eca8h93Dpw+kgnKGSEBxthMzGrQiLhzdRnGDfM
GPeKOVIOansI32FdjA77absYTkCsaEFvL3cy9+KT47cieS3WN75FQDJDncgh4c6OlQVtDslv6F3G
NxYK2S929k8zi3EkV+MhT6Jl5sJJe1QTcEdU46EEoCYribdO1XZitsmPckwR6q/V+DmlRev1UCBI
QfPGu/uzt1iojxAk+pHRqlk64dcxfOqyv11zztJZ/tGS1mTNIBqgIRIY24ZcHtHYnF4gL6QoNvHk
rEICV+98hWnrLMnawAFgHqAw3vhFvfTxqXi4HJbt5oLsFsH97G4a7HOTniQvYFCMwZGbHFW7wybW
WULEw2r2wcFN/YTw5b6oOacvLhjvKJRokAmFu/E7ZUjlKxxbnNzwvooh3w2CG9EmZS+K/FWuLWYm
WkPQn4/Epsqn0OeB48kAGD5a/e4qg65T9xQ53Op2zUoehUFCbVyNiH/M7deQfMaS3J0vlp6UUakp
hbO5iZXCSMK7rZkn8sMTl637UatMoAfGQmCaWBvidm0tNRoW//hHtOVN51fnaz4AEaKIzbFbXpom
ALQ+IfMLABVxnudpIA0T3P7LPfy8y3qe9MWNpLBL1iN0xJP4GrT+Y6U0xMSZrwE2f/RV32rbl3zJ
xajo7BGgHUBg+erHao9o1Iq3Eg3WBE18PrdcsCj6C7jKIXRhrrZPixzeLCiQojgPGPQv/OKTyIZn
Ujr6dXMzcnOkBUtoWj7kJ5KOZWcKbBGD96D0gwuE7rCOwssWs4y4HxPe2sXGvUjCx3SDFWD8sIEh
a478jNp0bvteku2uk2Zoeyd0YVYfRwGDXPQp47bCrYfaRAY+wPHyD0kPCgMRc6xkwg3E6rSN1H4x
AXifQ7fee+Iu1vawSwHDepWFlyog2bIsFs7F5JkUfJdC2nCGAUrGwAcKYa/5BZsR9Cc4OeEllYke
+LUakZCeq5rHfZfg8UCNIj3DWaMROoohNRFzgCjzsUDzh5anb/6JXmLprGVqFRpFQPIbTjqKnQh2
3F7nsi0w9PkWYBwZGQ4o/u6kH9VVNO+j2amW3/DRMJ/B4VsyIis1pa1fsHJa2hL1YzRrl/ko197s
xfZsfUGs5mNmWWV2sXrp0oh2pHCXGr5wXGqbqd/n5Cm9TFpFuUaVyHqQ5TAHIft/ysT8IqgIC+ue
7L8o2xadBu1xMacoti7v9kycZyZgOBFJarCZiYVOzqNnBk7jmIjZcvZkoXXWw9r27179SkBbnLxt
uQZZgX4IezppbkfWQR66GAta4+Gr9Sg6OD5Z+dbX7s6YmmVTPc13Qy3bjjmjEQPuyX2vuc0KmzYO
LfhEbpqFL/Mg54h/i84F7IeSn5sRZPIgkx/GdOIUgpYEhNrRRxpcLY3xKUUQxkckKqPmopOVV3A4
Agevx2eI9U3w993TZk3Si2UqxGviZ0QiCXcWMXo725Wg9EWrZ+8vwKcM+tWkoD1uOJqCZQPUU2+z
h/xHPFahck8/dPJPcJNz7O0qBvzmAhu8MotwXiBMnwSEqzPKcfzF/ImTBxp4Rrjq6KL0WJ4Jn4XT
i2eencrDOG4fa5y1EBxf9FZW3LetItnI4k0mGD2/DwOuJHxYXNzJxacFjiQMdQZY7PEQEGh8KjPp
ha0yiwyf0qsUTj0ptSaMdwdBpGKwLi2EkicdraAkhWIAoKWGm09KAEhhRg0HHeI3TTlRQRhCPo0z
u74Fyk1qABVU+JJD1C+WIzpRdGrTo2CjSyh4Er4eQW0EHK3UXF0bkYBUOAMcBko0WJNKovjQX3al
fFvk1zFkKW4uMvvyt7Ckc+2RVjxWYkwS4jRIs0xS5pKwjP8WvKX7PmZuprx8VmaT0KhJWcXUWcyD
N3LrkuzpCvbuV0/K7OQtmf36MKR8XFtmWC4hyiq+TQ4IFf8CDnFZL1vYY5oan+ea7qFg7+pPms8H
q7sJAOdXg6DbegVMBbKUBk9J4tUPd7KmfZ4GgCddhHSsBYgbSq/RE90AEzT7rm06dGSFTS/tGskW
8J0xJYaeY9mPXL6WXUvN/cRcQmxIiZNhWI3XsAiq/2hodWlfPMVi3omkPoOiOdNWoDLmW6SxYUed
J30sZsO7lUSGdMFJrr/D29XCSFhceSy4HuU9PA/aG42ytv8DPdFP5kIBHC6W/wiDD3xS9JvTxzbp
5gt9jAs78mtoczYFiARFEycBPPOifGFvyKzFwPltk2XawdgJ85eITfe5dKo9V951qx2WBn2hEhn9
1HLPwuDxMxcs1toj488wlSnuDKkSEVazkBMmFw06rZJbzXEKbTsqAJvqmlBTr7ttwg8o6DVTtWe/
5fdK25jr4r/BomykR+wGCtXh9A/z8acESRudrBhnrCGtDtpgfR5C0C+94b7FPNBbkp2Kpr10E/g3
zbcCrC5/AG6lBxrhs6Xe3JXARkV9XNWbppWcHDOOGAnzmrqGEyeDvjg+Xr1qGgFyA57tTtQxs8t/
zdxFBuzZQjsrVfPqZoSlGW+mOYDf5/CPBBPppC1K50yE9hIarU6dhh6SMqPBlLjg08aBBhJcOfE/
/blqi0cCihUXnJJS8sbjP4ql4xaKJFbLO+L/qd9dxj3BeoDek97B82q2Xs9DXx9JeKEIhbexYo54
n3w+XNUqkRt3JQyyEiRSL8EH9H8bys2PSQyMHU3hh/t4z6/94wUrSEPvdYhgmOzvG4YMWTzYyqG0
RrlPx4K/5VXGPBTNFDit4IUnD6OHkFAE74rOgMXjHwmV/CT/ixYglZfGeS/fn/JXwN8gWU94zJ+t
MuyRt7W9hM6/j85NSJu7YURMxm7443LPqoE+eYUYysmxLtLcoQyAt+dBv8gnR6w1VHpNXcDGSTuW
mACfx0SBgPOeeAwWbfXtAQCLkubW8asJ9Yngv5jQApaU99vwDpKay6gr1kbQPO1ZqGVsivjqtlkr
elcO71H9kQ6Fr0vJEK6uoG7MRlP1TeDAOCUsNJq5e8DaY0uQVNSOk+o72DGTW1+MABcQ4GgBx9Me
4KZqLZwDVtZqXlZBerXKFRilIsdlu01F35ss1GzlSft18Yt75qi2dvQvEHMU/tgW/FjrinsvT6p5
oQDvjGD/HclfQmsEG8n6xX7HtO5p+o4FQY7AyQXBJ7/pYp+KBg1E0h7J4jkDtj6Yghvslxq5wfQW
nBEXVEJr8V95ZJ5+SDlsFrnGiQYhwyRzCDvy9Q6TcjaQgUPG9bNiAuM/ERy8Xy6kUCzBR9BQ1sl/
jOm9w/NTy6rKyYchDc7ZzmJglDTk7p1wYQZ4cY3S0eWBStle+bUO3pu5kJTOfrRX7Kfw3nvboSfL
ldZBgEROOldhaB4/K81LP+PqGGUM8M8TcgAVPwNBf51+jQ+Se6XTI8Wjdqa454AmCXiAGUWbv6Fw
t25KxRgsKeHWD53bH4ymLZ3PSQgfnhacnuyAIhAFtpJjol6jZ7kPOdm1XpnaR0pjooYneq5cTQIC
9NhHBRxc/57WKo2LqNbY6j8llZJt1zBwq6N5lN2nncrJwjpLfNRsAcG+B5/CBdh0y3DdE5JSrs5O
/OUe6w4NOnokCmfFoigYY4b6of4DXQ+MODMlDO9IFQGjDmDosApU1Uzittj4vw5q7rUk9Lw/7DQi
2gjtjEE5ozFRQIES+59hNaRde92KWU6EUMwc9bPh78wxyycZWBRa3KJmuT3D1dVSXtZve6WGZztk
eqozO+NA1NPQQoZv2rhNgGgs1w5TFMMrWkHHyMfL35T1hanku3MtQCifhpYwa2Q9uy1ksso/V43Y
M8TxvnRIS3cA91Dzop0Sp6EuvOAfvHV+ZzedmOCAO0avUp6QOeKJigLL1TZV8YOglox/PkHoIXfk
FZCvDIFlLoIplcs39Kp46sl0aRhlbnKHAQRA9zVBXFRv5MHtF0RHT3Ar0lCq1dwKvSuU1Pjj+x2k
ToEn9KfYf0R0nE/xvpa3U7nuC/uDWv0g/oGzwT6VfIG7e082U/IWk5fhQJkzdxZcApLTErHieGLb
JCSYbONyN0XhRE3XAWirFgc9DvESvloORev5Lo0sX22dg4z8M6/Eq7aKOdnADTCT1P27thbdJDSY
9twhlOiDmwp6i+m3CFGTS6aNQsib+EkUiEvv5xco5tx6YQMwcWnx3CbQ0NfsssChV6S1Zkm+noEw
R2HzXjsN7rlxKxQvghHN4UKO2Cutc7TaU51xFQZeS4LZ4h1u4x4Pv6oILB0aeJUUKe53QKlAr0lt
5f3QmZxH2qemusPbDqpAWtKnD6rWqq5KqJcX/2uuYKVTJCIXxmyuRy464J1ZDLV6y0O/tm/VowtT
JuS4fWHs4WZsjp2iCTrMeqfYMaxD3ZMuKXBrSa7Bbg3AE2b9MFL/LSQLHs5SLKEINgiilc+bIRnL
HLLGeaShdxfb39q2oe9G7rm7DxPahgXCaZloj49vquosBXjgGetamZAdIVqHsZQnEdQjT1Epx7QH
iVNYxlqvRgKMXQakQ4h4WR3sNej52RPhtfcdxhsJQk+0w8Hky7jDubJ8MkB2i4WBC17qY4oBLGYB
us22AY3UoMmgISyH90K2KQEhcDl3oOHS4LT19qdZyCuLfbgqGBQjOY+xIDswTYMJJ+yyXjsYwU1A
XDHqV9u/xMXMcmgYVNW0syc84mTWUaYq1sVLSywZFlB/gBgXZVNExqcFnoZ8skpC6CqlwD2+wA7K
d8EEShmmTrMeg8IY9mK/UPni56FEcK1YZKzNHBaIdd+lPP+fU3iFwil1vQIs0tcm8HjVkzrECHSF
wf2zn6sVlWRu/9DHv9OSGdzFdfAZKKwB1/WnAXEonzA1zD2+a5Em9YcWRonLFusYBvq5HJWDyJD/
XkuysrOTopfzIdOyj0w3zLvgy0/2AU+5609pvKDNqrgJVqunu6nY0aF83OM//Oe4fh5s4N9eO+Sp
bhrQOzYD0D9ldl6dEvE3ySbx86sRJ7//2c/e9qPG4VKJlZin1sRbYDGy7ObUcK6RP8ceIyNGnQen
inE5rnZ7+rzvQ5lOCY6a/QGrqvnpWGP122CQCPsugoyEaWAHg03dJfJ8ytdstWW/eokd4lLqcrUI
LMyZdbhI5aaQ0Z9GG2Tc5bL5m9f8tuZ8I3YNyuHugTbH/EgxfUDvx11ofcBVm5BjUod7tdliq844
hJQIIwaTK+kBo4tfblyXmio7zt9E/flKvH8tbaw0/iXMzDEiC9weNZXKzSEq6/UaZBs4toaEJjWV
RxSJmi67bU6uUluz7dKEArmeU3KtZgpqyhJog9mpOmu0T1zX+GpW3rmWIMYCkRgaY90LMPyFHrSG
PEU+i2tSodnUiQvdKzoa6NTqvOJ1FEMkPUpUqXn6u1VtZNmhk15S0u2F07CJzATTuqvd9vVESlHI
vck3uB4pumwFv1Uo83R4ew9ctIHLKjs84A0UHko3hB8TXWOOmgOmjPKV+Xh10Q3czlmc58maii30
Ot0fWIviVdfzlpppVHpzds1jKQPoTv/KALGYd8dLN5kAarH15yCOHX0lXPAMDSvz5jyWGqec8Lf6
AS9qwnEOBDTbG8c8pdjG83EKeg5MB0e9h1KJkxwXknbk6ZipyzlBOCUv76IL1Rm4beaTPSVF2Fkw
MX8fHJCwbcQKhe+lO6PwYLiT8Pw218UQP2XmWc/W16xn69geKs+FpL+h3wAqh9pgGkhKOW5LmhjF
kJdwtCxle620+/aclUYkWoBhAnYCmo6+yytThhHKIrh9qxhDxnHgxSdSrALW7HQ1dvedDi5C8g9p
MYsCCzlg800K6mS8wHy2rXcQ6pY89Dec4XX5kff75z1Lij7sbn7Ca7jqsW1elZ8ShyR/tpeN5XkS
xqMF3GUMY9ttP8px65PasCRQ0bMBSJhgfy8kGbB6LjiuSAsVzNJY+FNBXvSPlSZW3KOubj79MPBV
QhgIiwBQHX03nLsV4lNCj2oLtNSPstlTbU8jAlTe4mdYQIRNQS7f95tWlXaUQL47OlbzLWZbpEAB
QopfwXhoa948u8y1mWjaIObp2GS6hqhrnrWqDMHuyb961/RjspGy+EesB++7SMPRNzxR6QcNqaCD
TbWTmLUWzT4+DfoYPeEg2thIDXQIvIg4LIBaqmE35JvMUnhFonMkesxnqfVWzA5ckGkA5dhZ6xab
bqyB4j2uNC8dPLP+DtsvEX3gclqU+E1P9njLNzqKteFFBACYwVkU79b7jHicQF/IR/rVCkXq1lXV
PHl9Y1Zp18pOcRuHL3iBuis64QcKusOXyLnl4traZy0fdBYyceldTZViIVQbV5g7Qsgp/ozxFfVS
Q3G5VGlP4HKvC2qlTHdOBHOAxXH1RMymV9GPAGdxpPqTcy2ZmLL1LfykR0wG8IrYTPMAfWAM38CA
kFDGhVtKMtYNs/D8oDCIi/ieW3uhYHUhJRYy2Q1HG8jmmA/b+kIvyoegCIfLV/PyJg4d76AmWdIa
RP06dGvpdDAIe2aTnvL/Aa98s6XvZIetw1OeNs1Nd+HcdyxWu3Wngblqr78beK2C4+IinDpzpYzQ
/GW6kE8p8QlZTuceqdtcbAimDtknuRD9fQu9QRDadskk1BZeoF+8rBfadQtAPxPtk39M07P9uMKZ
R8F64Vfo+BlvnNQpgSR8DTKuOuxnK027m5WbE7sCK9DKgIFzYwcSAfV3RLXXcJVyX8GFnof9CSpK
qTwnxzf+ulT0jzqFDhxZ2nb8TN0/rDJMtii0OzE1806pqudvZyXXyNPzMm2lZnL21BMQu9lizbB4
aWUwM++BVgh0dqCuz2pW4yk0k5EyDgqNWhNRHXWj0jB9piyirgihsBrhorQa6clyznQEUAtPITk2
dlanaYeLlleIhFG7udqQ+mxwCbiqwkZTys7Z1Z5WRSB6SRZcAe30dIo73700TdurT8f+VWcohE0x
en3QvDycU/cLmt0hK9WbOPg2cr2lTBVpTfjHJ/0mdErTFez1xRaJZNQoSOjws4tBLPdaMhNMVHCD
gNIt7evqATYTshJ9ygGrhK3eBOZC+RFcIJq+u6zZ9EWiOwKqBYS5WjRLAU+6xuySX5L8QBS8L+97
mKO8wz7FW0ji9Opq2Pn0of3BhfIvKI/e/4eVORy7FvJBdl6aAUTlnbtdUnRmbFpAo+DLS9RENJxr
CiTgYlaEmaiO6kDiTflK6mAciUzgl34r4pgE0OpXAmDvxFHIA4By08XGEJOdEY2+TI6q86Bu0Zu5
FktR0xqfdoOIwdsIpw0JGEjLqEPxIcjmwVRiPrewgkR06f0iAwcJNO3e7FA6L6VgonHsVlgrom/A
fiUdFPhhEm/ty5i7xYA5IT9bUvFxRP/zRByADCLnevgKP7ucJFs2rl4TLTepv4CmLeQFDy+UUZgR
Hn22c/PWvKT/29veUppRYmN0aWjyR/7vAQxNsHMExoWrWLCu2NW/LmcMPLClvjp9zp4K6HU5LYJy
PfaDv0aUrKEdSJ6PC2FDTGjadGCYUdr3v7yfMn5ZuJmgSEEgxryJOwVGU6PMGqI5e8Skds3bbRyt
gIsX0vlqFO1Kerg9Y+SmTT/skniiH17bWj8K+F+l2Nt3fu5Wf51dRgTS0QzyVtqFxEy+1CndOKKV
umvxQnc91EVCouQwHJxXFiq7KqNcLE6wuRIuUxQE2Yk9xinTnCTpRp0BDnQY4cqA9AKLMxvj7t9T
3x1WSTjk6IfKBhWqgz58qJ9vwEOogW0+yJOeGUx7zo0Cu8Cgnl6R4K0mRnZTSkbofJqpCRQyfMC/
nE0FBYT0niX6+XEtz3sJC3JNWR9mXOaxHf1N0ZRZ6+LWDBkZ+LylvxRNHha4vJxZOobv7sq+YYQB
wKoArRq2JfZ1scPWkbqL2Kz1ljCZ6HyelcWZHwz5/6frAF+PRX57ittuo7A+BPQC+VNbDojCGS+y
Z91+qAYtrkWK5EoVg4nl4/RaTlnwCidUT/ylhCBGq5YsUA3va2+4eBgWBYCBqykHDsm8uSs+JaST
YQAzBvdu+HfKasbFc7rwA6sUn1G+bh8w6pUFJ5wdDUWANG2ZkbQbUqCuTcPBKGKXk/uSxpu0LJx+
J8HZbwR86YEqOv+C2HmppeVEKdRXPjsihxKhtWNa3sVjjQNsUx2HNvjalFNJ1UwTEnvx+Z76bYK/
z7Yl974Mqn6gDm2mK+5/lY0mP/c2IoIoWmojO6H4rBjzDoLK2Ggp+rCxR+0JyEW4D7jHSbIuIjzb
m09JfajtD5k9EHbKMwE0Bs8L5gwxn6ANFb+InWkHBfy8NBNHPmRRrvwRfnukCEJkI+nmGcXHFrH5
/NQKTSWNT4ny1PzsHypuMF5lcHUMLJauS9iD3BUuOPm7SASHJodNMLR9XpZeqBo+2sgPACktXe1F
BUJGPil2MueKMDB2aj5DpkWvywbba0RmDo6DMURLISbNowAgLEnoWxpf48fy3y8cwtU59lwbp8Mp
4pPBvZLsIVtj3s2tD2nVrobCaZhMdbGH2u2lf8i1u0xTUEsW4vfcxcbu6M+cMCyWZktr0RC0Zzm6
4w0RmjEYwEZh4OKnH2UUrcYnr1NzK1zv/p3LMOCOeVsOg4hdXboSOXACbL9TqBPJh8jXjI9z9eQE
ySzgYHhSIiF2tF504Q3fAusg6swCPGXhKTzgcV6ctsqrrkxKvCYffz6cSGGSpl2vtqXQYLy8ltvs
FwJWw+TK3DjBqzq/OQq4G+gTAea34wB8QRZfj280JlxwstLzGtNW6j9Ffcqe6vlowDoAwTL5HdTE
V06X4UcGLjUguSavHyI5L7+cC9pWKd1hHeh6HpekhqPXX/pUF2VY5e1TN888SrUowIeyhp3pe271
cyZL6J5oq+xa5W/oMmc/P078LiOpuMRJoDfyTud96nAeJr/GIZtNtAvpw/oXeOAvrQsyl7mCZnTw
6w7Kz13axCTung7geQJjeOeVZhBOWfZhvvHLnYTg1gUEJu9aI7C5VLD5ClQ48so1NcIi1uxwJtZr
akG3tCqyRpBEa1AQigFdrCPNnh+2EMxRySV45u+XpuFWcBfIc/1iY7K/XqbxVUgZE5j/ICxbkQ6q
7KKFPhVpMcnHN7bSvSvfvJ2CgnEjdws9qV8+Sx42P5fw8pmof2VQHh23qjc1JSy3/GR3B3X0IfV5
hNRn0a/N/9Dwxhqvvpyr4xaFU/Mf7Yg1hOL+rCN3/LQ3DUINisFp6mcGTw45mjp7vb+a8AQZkVHh
DkcGZs56U/F4QgreuP7dklIzWjXZNSeJe3YH4RbQU65tOgox3QPjMwa8JK8X2IevhkkCgKEVZqhr
gSqsucgNjYRyINKRJfs0a6WITEnm+27h0naE5dxd71EN5x2Ui47NAGU2ZndHxyOv97b6Z2XI0ca7
HaIdtx7/RyfHs72L2FEHHk5yCWwybQmSIPE3iPIt/OzsFwAkhFtVmiQCluL2ZA+NsdWvLDVsZ4c2
abaWL04yQP0+paBAUhD/MEZTWO9NTRYsyRf1UNrYYq9vQiKeY9CYyG6g2MVZxh6pon6EGN9k43vB
Mm09ZNZj15oKx30cRE3OlIKiHUkYza6c/mfnOkV6HGV8YzdkeoszkcZ84gNwMN69t5miremz04em
f7vU6yrvvO0WM/1aCNYYWNfgC7dkJVYtywONutheEsIBY0g66lORqUT1u/Xan32bfj97HB4CQzOj
y6/usB6jIA+sKpCSQ5XO0R61p1UTDlYjBKadYAcW0Ot4jQz/2BirqJIKPPkChKNoObTwmeTryjtc
F7dsiB0yG+HQSknFgIw3Lpde6XTGG5lzaaVB0c3kh2APjkoU5C6qaQNYlGmfkQG57iloSibu+9iG
M2xlnjV2YY3WufStJupmWiz/J2g64Cw1q3QsukUmhOciG3LthwnljG3DTAUq2ziFVbTnHKBO/Fz6
newHk/BSECwfTHyMMTAeuIuG6eBaZ3/dE3aOQRwxM+t3dvYMYsNbnCR/1rE1ZozJvWREmktYC8Xk
co36ED/G7VLd5nvIlxboSp8xwKIMA53bD+rrgOnrW+WVdmlUJxMtMjYq5QPEcoq5SUk+VhbB6H3N
PGOWKjjgEXWKHk3pOkOCSVwnkOOCgIdzoSWDpFwLk4r4HoKiMs99VsOLOJLOCEXV/BVr6toSU4Iu
+qSSD7Cm8JhFnJZdMcrkCjEIkwKxRUlZ5ia1RnbCEovsQ0q8oxl3u3/d5SzCWWUWIBQElYcRxM4k
UBxO2cXL8hC8XjA/EGtkDvbucnUSsYPrJ3rtrXwRpl43MyoFJ9uhauXw7NzKv/8Z0uZFn0nT1ejb
GYpDBXlqVKzGaHeC4844MsLLMpk39Sn8+GJq7xP0ZcPcwuQwxRuLt0x4S3woeXJcfvavvjCRRVqy
HN9wSOrzZcRkDDJuFeXn6pOeSqpMRC4pv9uf1/xdMI+OwDi9ha9h1x/hZXDSjnhHnXosQSXIz69Z
xlui2NDlUptaNyxZWiry4ByAHjGp2Mg/MMdtj53i1riNfrh49GtJn2mqM6cMRVBZmcDNcuZBsHWy
3DBtZfN0Z5Gg9M2VIghx+CMQ9qY+t8k9TkFjMjmFeZBUj3VErl5kXRD/Ij+LCtNz3vIK2nuUYUQW
Pbgrakg/IxyN8w+eVNlbOOzltfbVKrvO6lubrZQgpcWlU94eI3HgmzN03sqpdH4O0HF9DdXt1f2Z
NrLYFDwZAG+DpmGmE5xHViyv5kYwcYRweuxs2YPLP/LMFwwAY9yuW6Ecl+ELVhnghLofXHhdYmz0
SVMyi5y5HaTRLkH0uxsqNTSH6z/OQqady3/OVED1IhMwgM0Mar5XyKDleGkMyUS14HW04uDFVNl8
2INGyj/3thV9NfYAFivIW35I01KMCFaSY/bWKDGKel76keK+meDd1esca0TuZGnKMhAZmSlPxRcl
5l2q5bez4cIKx5Ywjj5qOoVSczf/HH4NfnKjDwenyVMEFY7wqBq4LHPi+1ht0aZ/nB8t57RGuV88
pESv1xr/51z6KBNqPP+0yyEMBbRyyET3a4jPKahOFoqhIVm2TBcWAUOy0yoAlyl4EgIRyP2sb+72
ZH8J/bPpg33WJ2UMnTnuBXY33SlJ1/55PwuCad6CWprAgSsn+TYFbkFEhCeYC7hY+Sx+/R5PlGFw
Cwi0iw3yjsUumDvjCBhjIIFQgkxYeXCfrafXyzWEAIHnFeH97qIImlNsBJf8XIHUMqoagSjYKld/
yYlP/omBJdv5PSfzP4tHnFIK6QnX6emZiQswb7bfUcpdzqrrP+wT5cWlqARUC0VrciIU+az88La7
hQFJo94S5HXdZmfzZ18wVY/RVEDF/ksX55XMnoL7Is++LrJXS9C/u27v0OAojAfGSLDUs+BXEK0S
PLcKHRVIsFdAAiQLbFjZk4v3XES2f+BCXmAqfLrQcDuz+KJJRjYkoBR2CySPSe75RUqXbJ8AwX4L
hhI0vwD6V+wpOrYq5BPjd16kRaanRZ46ul9o4kE8KsJrdCyl+IkaM6Y1gF3PXZgDxxPV2fag2TVr
j/uaVHu37vaaHXL0sWjDmiU1vpAjl/rPiXQlK2j2tKFXBn2mUxO+8qbpg1TnaV0QYiSPC7mJ0JSg
USQnlJEPM3hIeoJG/ILlIqxfs8fl2Dn3HqJV6ezIODEtgmQz/EpXzlrJAVNnm4HXTfUA0znfV0Ik
BjYaODZoRV4LMSI+lImhEcy68g/XDgna9yIIN0aSZCxQBZKFZPFk7Q7TpspyAve4K+XuU1rmqeCX
NkD4wuEKOifQHI6aDof5kh5cVNIekZ/mEvTPoPJydL6/VC0bpjDzTWpXA+u+oEP3BruMa/mZfjHa
oTAyg6YRLGmjU/9SuHWdNgPZ9BBbekeSCu7IrxED3e8pYsTYFeD1WF4tZdFn+2aI1F1Y3HKxnytE
V2XHlgxj4P/PRylIVSRNIaU13Q4avEXe/f7LD8id/yGt3/4A5vRmt+wJlXoXDkdpV0uOkrYTUmKR
9IuuaHzDBdSqCFB5JT8VVBlZ39BMyMWNUoyJLRqeMZoule2rfNkhSi6IuaOMckVmwWMQauxNvO1z
drSBLodw5m81+RSkVn0qCVyP/eJ1zTVniEkfhiK5zdXAO8Rco+E1Ah2CjMGsw++dfTW0NZ0dvg9N
asdOWTiai0NXZy5+VnYsTh/E3C5l2+K9mMMwP4bplXqJJkyCq3Zi9Obzb4Z6zzqd8du4XiTVcHLk
Ho7fHRH4q3lNE4lWemfc2TgTeIR5Zmm6CyhlNMZDG72qBEjjNKXHt5o0IwuPHwDD0UmmH1huaaWv
sr6SpzkXHlpv/JlhLHvrS6pJCO3/7UJRPPtFzvCHshl/gOHy7U3cexYRWkxFsJQnw7B8QTTfPlyk
+XpclHR4K1x0UvbNr+azfzuo3NsRFPRMfw3CSdiI86CoHARt1/Xh9PA4TR/+jjaIdiCXH4jXKztg
N7o0s7yNNX6rdp6Ctn5paYFXvY4z7JLED8qCDp7ZBK76ycq3F05sxxt6r7BcPbchzks/qa9SwlpL
20EJ9UAVl8XerlIuPl/zG2x0e9wOV0ZpCx+DrMGliMZmXhcpommf7ET5IrehkdXRoKV6+Xf93BW0
0C7va5NFKV3ti0PBfnIk6GfKZLYowr+LEQZGBX+qYoSGnYOUqeHIa+OovyYJ8WMPFhznnUF+B9Ft
ghD9sQG6W5A34WtM7OxnX80wLyIr+sCTUvBOCeu/cjS8vi/fNOvY8hR39KQLb0a8x+SaVscSLsJK
LQMDvduT6X0ZJKZwZhdOwLG1amitO3St1Hbuuu0lTGbEnuciPdLngU5/HZwH/X2sW099Pwu1eOIR
43F98i0VnDTjv1d7F9YUZCYWq61sPinqNypyttFo6GVsaU1Dyd4tw3VWrWWimb8cit+fNuoIAqxE
VDB5D4NKq2Lx/o/LhikFj3SU/4l8tb5VjbxdpCYsAv1FqtRigVtSADx2EztIq1Q+ccp5fMYKeffq
msRP6onH5UOLJp+uSb7WNWVWmkKTYCuja1CP0fWX2KJRxrnClVDstM2NAwfrZCqNHa5IlXginhDS
YXc3UE5aeKKre13eWCUUn6zPSs3eniiwPZ1ohb8pOD2GEsrUr2XAYMXUCRnauncAJmAEmyQKxy0B
V7RDrGVfBr98yHgM/afQxCAmMAWJrfzammqOHQ+s3AZ697OoIF2+wHpEXjwiys3HDv+5UErTzkoX
3xUO6jG1/hSKD25+dYNV7U67HF4/QvRhxM1tBkd4O+YTKMtsGE1P2qeo9gfdaKGJg8CJLO4s6he6
9JP0qHRwfDyBggiGPsoK+mQWuY+xSM7L4gE7GsZBLHa1wyBKI5/SG5SPqmbUcDn/sWrasTjxrBc7
A/uJ7YsKS2W1Mx6SI8lDHDsGgordPUJ/YGVhzhOvUGg162XXXYfUSOwPHICgjb10+Tfa9SG8CK6x
XSdYVOyxDiLG5u8d3uVLGmFUYBKfaOXFSb6fxwNTvHYr1u/bOJsBYfL5Kt+ajp+9TkFPodT5WORO
qxL113Q8+tcg6j/Zy1C9ddySV4DCJllrGZLN+MmzmR2lcBbhbxtSnvlDghEFBKtmLj+sN98+bjs8
UKuJgawbdCDQZGnFRRXZ45vQTVnqcDuTp3Bsnt1K9nlAq65byZjNPVV/EpQ4cd4kv3Q3xTZwGM5H
IOJD5hCJk0S1WXhUkOVry/ou2qxtxOJUIp3z4y6EzToIi8ngQplqjw55stybRefv4IDxkj77xrOF
sO9qXKI7hWZpFCJ3NC7UJaRHwa42BkSWpNK/94EfFPQgikZWhv1OaAmEsPRfKOQpxWb92IKIeE4d
UE2suMuPrEMdsqpOK2EcRGUEzE1xrAxhBYRxEKavOeupjIlel3qI63L1rpU/n0Q+GO3fKBswwpXg
IgVRH3LtPxi0ZP1wLDP+XTChHNWv7HoJp9W4SNOu3PdXt+sC6zgX8/UCmqinqEwk/JR1eSv9S+m7
+JLwM3R+lWXom1Iel8KgHviviKlNoSEhFpW+xNHARKnvhLXooV9vrCkPMybwn4xamw4EzDQRDY4U
ZPHPCfvoMJna6ce+42Dqyk44gLy9VtH9Q72ffQ+HQqyqdBKzq3IVhcJ4jMbNaKbmZsHP8ke3JLvf
+xO3duySQm8yXHwSspIOWlYILeqcF3Mmwgb6xUukAli8Nsx/8TxsLBIu8Ez3JaMXvl/oXoNR0rAA
N6nuNVb0dMNS+ZTK3f3bjrWMEzxUTQmk2fv/wIMo+IyfhOY8/UrEds0h28e/Svl5cd8/ZeEBAru0
Nkb/AUhuXK5mHziVcnxLxcuyz4sFYWVqcbr3Y2pEM+2jqlLFZBYdJHb6u08SRL263m4GGFLZSjcO
t4zPKfFdRfuCbLzRSDqd9eABR6drZfSy7vsDVZv6tto0vFvPaP8k+2T4PiXqqvZtFTk6xPvI6zx+
H0ckbkgq+xMuKYr+vGKcBFXx3EH0sZJVmkulp+BHyEiiprzEfhCzvRblEishmvF3yvTlaM5Wo2tj
7iUJ/a8ODykICwzS5w+HNljxmktXzl3Qp9t8RlWoHfwFu2vK5NCEVxHP8vzlsheYuq1b6GLBQktg
eFGpiqr7nc4KRf1pbaXsOTPKUKQp9cK2pZ5i5Rm0ffsqieVfUS6aoYY2sXi+AygN16NFxmx61Y65
8d9qgr8ruLPJx7EVFFuLzAPxjVhGUTHlHGq3PLFVdzA8xKc3O2BLwLMFkl7WYEsI+qjSE+CzAHGk
cCWGWiYa1rzCL3kBbKO2B7nYkso2ez4Z85V6VDpuov1cwhfrynxC08owIg4atErlq/wqKp0ljswQ
M5grSPw8p6DGON7oAN2YPmQoGIa57pLQd/gGuM3yjDWwsi/hlVM8iFQbW9UVjsz2QsbKCDBJSxMm
6vZstssmm//i9DRBi3xwDXkVSuvDYN7wyKbmxIhIMdf4AiCXDZZYui5xQMrGDvdGQYifnaJiFYKE
5OGZMnCtiiKIjMFr0qHRxPSXtjUEbUlJ+Gqy/Oz3gAJDwkXQ8k+2ygCwgQZiozBlZnkByM39GGQi
eqEL+Kj9fEtwgutUMMmuPJbPsK9LreKeNJ0hkHPM5IUavNZkCXxOCSfM+YA18gTtsFx+gYRGgGiY
W7fkGRmxREvE24udpIiZdVpaHd+GlkdZtqILsqnnz+zKigAGCB+dmvbjz90IVph4PF5d0H4DUyiF
NbA/ERF0iAFs3ubrihX/JykkG2ojG4gSecBHtr3lZyS2GymvJxVSNBQxCWnxTdT2XBLF87dEKOqL
r1hAwFfWrdFEdXyyAa0N0BDsSXLE3XUmn5b2CLCmvMe1AQ4Kw27FVZVloBZIHPW8OGSLEOMs6/oc
/7609Hsdz+UqvX1H8Aqu3DIV14r2Uc7oxuJ/C5Erm0wZv8fcpA3EtDcBWlqTO5E9SrGrkK7SEZ3E
UqjsX6T/1x9H99YUWEX7Ol4jpQKDT+KHRGnM3xfkXYXh3KFYm7d7bxiJwMOBv0ErvtSI7ppzaVhV
LVdkgEyym7a11G/N4jZTDxonUiufCfCrom3Jt3yfeAwCVbXVHbddfzZNGjPdtxQHPRH7z3CJUEha
GnQQwZGCjgbZIHPDO+APTldEZvMuHD5fFrqtMn68V8FukEegvc9GykRmBMLRgAStbnJx/uUdr1mG
TbeWLrClN1ud8pg8obgcveTMEVCK6YNLuTzspOMERAsPytsIfL6jUZUNePH61vDUw9ZDfHn7xkgr
z19FDu83i9eYb/ZDijO3S8sGqaXOkV8Lq9BNGeQiQv0QahK8CdUP0De5+GNlniEZCCR+x60kkWey
bWyVwjmKDJwbdnhDAULId9fjC2B8Q+VpRqxj4Yj6T9ZbtSM0p+Z23LYW3rgt05TK1BEqTxmVAaI5
mWb6KP5g+dmEi22ZYbrkjNWaKH/SM99ad2owlXu91p98/5t0S+I3Cmy3Mkn0Oes4pGxixFm2JstS
UmG9se2V1BDzwi2RsVHSQiC6Nf4LKpTFdzQQXJHO5/tylI2twWHa7RrbaJ6PNF7gmaDwCM46XX3V
2LfBUe9KV2pPlCQg25sOac4zhzQAuLrQ+Clj4/ZJPV3dr8Hgs+S1kCfE7UBHQLEaRHDBrihwQEqH
6wiHo81qNThNFe0brBGwEEC17H4TXPaMYRnz06DLLiJ1UAx2hv2eLcuXAYhF52mzsU1KkUeqs23Z
BEtT3vh9ujqrauYcgTB/V17dTFd0PQtjXmLJUA/Qs1G10kuSb4Oa+21eL0g+hHib1cUpz4aNbv4n
RzxU/YbwuK5IUKpNvDBz1DZnq8WztPn3s7WRB3VWmX1JzOGqAlyUzvTSu8rO66Ihr1KrM/8amJUe
0FVgRbtGeQBx6vjbyuJk8xvj7FMrL/w8slVYWqvA7rowrPOPjEAh8hS1bWaopdYUEHdTxsTcjgkZ
cwq/N+mKs/e9uqIdeO6NrBp3m0q2IuaSuOs9llNDSfO+Q4bNm/eF2pffqln2bwdrj7vpvITGoATk
t0Xdny0GVvyAXppthWYfjNceZAgV0znN4KnojVGrieq8Ilff3oojQjDbvLPbhHN4Lq8/xh1opw6i
kpWX3PhG6V93UcQ/gi8ukd2BEMYlllMGr6li7eTebgI0UMYdyM5n0oEiJinyCHkDgSlncXyc0+es
zrF22s4gTvzpvCnJ4dOYEEYBywYHoBxXNzylUFC2SFGgq3H3MVU1P88VLHoNBHBVmtEVBwVEwKaN
4uj/SOa+s8UNb8lGd50fJpiODiL77u3HsLFzyGqx8UzRjtW+TRKTBEs1VblVjsaHRTajkIHFXVPh
Yk4Jqz10JSS8c6ULDxDzlBo7Aw8xXN3nm1+J4BV9iokmKShrx6d3h6VkvRdQwPzIpIwbFwQO7Qmn
KKUbwNTlF6DpPHcjUkf0czmd2m8AKzD4Ge4Rb3ePMmOQlJSQYN0fABPhOZVs7REvx6Gf+n2CyOIX
lnMtgzSu4dZBreAoSL/k+qe5akSG7/rViym23A60u7LWpRbcu1XDI19Z8jpbsjD90xCYez39AXOT
pxt7/iJGT0YHfiy1yJCwilsSn7LnRPvx5ZS7zhIzVGdKJVm93PuJRG2pl0LsR4QdrY+z25mzeini
GyXczLsQYZRlakeKgElVE/2UmMQCsXY/5zaYusfAITuOa3POa3hDSU9O7RPB5+5wcGeW6do0Xh2o
CM71LlKflty/MucyB5iYnbBoCzw2QLFyMFWeH+mjf6ImIfCtzXdNjw78lxjJisT27/FnFH3fIbMs
hAqYO9Rh7M4Jg886JnU8bpYeOJJNR1fG5h5h+AyKC37gsYLC4Pp41x3c90CcfNAGlSx0rxhSpmss
pBieFiUaLFFsz02RFPm/s4vmQl3xWPSmshIv4DFHblz9RKmTSAk/EtTSu41xMPisPkBX6C0gAqVj
H7y23uI5K12nVWyNaVTSCjmUdL8Rtb/iLCj54ApU/4UKhOZgafzdCVTyO61T2gHrJajppcq8wRKY
RjBTaaJ5JV027W+hbzR6M1z9Scoe9nO08eHq4suQh+yKHdkH6nAAq16ICKXgpfsrSitIm27Nizsp
lutMC+t1+nfG/7+z1gCrYjqjlAH0TJXBnWOFs16agp6CnCqrF3UMA4hFNEngbcv24LJCJcgACaK5
teDb35KZhQuL+6i3rD5VMWUnyOe/u9m7CEAzDHNJES+cSjy8xxaft1HP7RnTB83CFRNqfOvqFOEH
za8S66ps+DRh+KcdNIcSJdlMsuy+j9JStwmeiAgEY+Gvh4yqCXC0oaEU5VgqWgzxu6k6A8xL9ygR
+4gnPicaFGIxtXqKRaEbBa/NmusY2TpkKImPhNIJsVicZstWrLQ7xtQyB2HZFOURrA6dVN5zZxr3
DvhxQWUQHfvetMZ/8Yb1IX4MFHC98q5l959dnOrcQbfMsHwTC9F8MX2gUuB+y+/NzIXFZ2Oouph9
QsicOWwFkEXacIkCIGweItMqyJEcNh2ebO36A8+ziRXIMhatWZ7EnFLgO8WRkBuCA2hb9gUpegJu
5iomLns7487ipNfs4iaxteGK+F0P3fpg2/k5G5uBqqPnEjq1m/P5SUIHM4mo9RmHELChlSW3UJsX
Vwvk+IiLUDnXAeROQ9Sl8I4GbwZcqlUlNon3BtcrhHyKUhZ6r220EevNMWHxGXjQS5Eh3WeUb8hu
FmDCIw/DuS5KUkDMr9AQmHX265Zzj9F8EXPoNDgOcj7ddPRUosrQwxM+CRelrCBYnWiTbQpnqhVo
D6jaeyvK2OY28Q8mILIvsI0PG2SqkiD167gocKzJWQUdKmOJ7jGF5+/0g5IbWj4HE/oSNUpR25g5
WCqi53m9B46wmKAp6+1JTrTQr2ENshTmodcGzEON3NAmH9Cnn0xvWVwb/Ic3f9648INq6ZjIg81K
YxQIGKWhL/LSQALMptn3kerxxaYnXrF2dgRrdsuDaJLKvZTs5+rmlNMHcGgfV5FXGyi8LrKWqqWC
B/GM/WbYnDI/eCnAVXfjwV6rgdUs/4G0HO376kMYOtlwGXj9FikYjuLulUHl2GynBm71HmU6vio+
fe8RPOGtdBU4LnoP6zbzKXIGUXjZUbbI1AGPhlhc1OKmXeEmqiZ0igdIU15M0o0awSO2ZDs8WNHP
gD4GAgrZ/BR1c1Op9gyIrLpkTntHj0drjpqjZeWe4nTiRz4pNh0snlqnhiUeIUOk+X6IA6ItEQpR
0Vwc7/0V/jNlH9mWeLO2KCBEe90iDclypGNHh2TY2rEGbw2QUlepxf0fPnq/yg/MfR5BhYX/3ecA
mBr/UYmqDdvHMNyX0QRkiBctI62LldCYyBs/CpfKPEx61cgmKTlr6TEHnpLkXnk/VwiM3fbn+umZ
h9DgawsZNYAvIVt5jZiy7V7lgIsk1eTHUXtIFqgru5Lyc7i8s/qN4RmcSnFi7ww2KcNjpX9S2EGW
bSnREEttGMjilnpq6MqiDjkVK0zs+l+96to0g7kfM/j3HpKEYT+o96m9deCl9ALsMxe7QOqC77cb
foGjX5YuPDLka1FbZEUAbY8kxvHYMCTowM2hgzw1qVQ5OBkoUSQSd86E2a/he89UNuu6vOYi5lWq
iczF47/pKKzeDu9Q7X2BoJ1xgYb3fmtxpmQNhTTrByf47L9NNJR5uXDGPQZcnwzkvKmk9rWZ63bG
TnZVX1LSEXG2veUxYZ6zI4SUGYCcVSFYoC2jlp37MtoAbFw39Q27bPhsHszEwy3Vgof71I1Lhseu
VB4ENPgq2gpcq5S6gwzzrnsDtPKr88btMik8RkRhNyea5R7JmYyXBS67iS9v1BbvCQQb9F8Aukfv
8QctBvgMg9ORY7OPjXEDsy/h3BQ8zzInwD9CkUiFvD1e9ap/7nfEc/pC5RKdRyYq2FLfOTfosGwP
lw12wJP9ksdTN/MCQFemSdn7L+dtMoWnkiZCWxoIDuACfcsDsTzOvGVIhi+Z2HgWFJx963I+vU59
JSfJlbJqAS53uMb8o6YUQNW8KFRCz2CL2XktDeh2SEe3MsJp57CPyKT7mYvZGZdXJFZvCkjA4mi/
MS+DEICid+a31ymP9I1ZxI1YqVLLwuxqNb9ZYUAQEPqP3fedZJFNoYQhmEP2tseDZNqInKufJwyM
sbeXMWnzxtOzV3U+pXzfbYHcGV9fBgoJbH9hLJHVNAjcMi73m9kR73d+C9SIFeSxK32Jb23UsVuE
aNilBuGyxybQEu6CqGq908aDemtmX6llrfYFro67vGH6LywcBrVqlO8WPBskkJETi18bWeGi/DGd
fRlxu+uQOgDo1oUZA6A6YTTI/+s5IP17mKwPZ8bOsb/iTx2dVLod6LRNMfcdSGL8z0bfkLYCOvXA
pVdtLPClmnivX+H0Yy1a6Fqg7rwLcugfyU0Sjqla92i341uTZ4SsY8UnNjr2hrJTykbfrhC3mqXM
xeNCFdHNul3wf/gy1z6s7hghJTuBdHxRamT+WMa+w1+LkQAjuTPDFgumG3dPsgEy5+zDOBQDc3WZ
1paImOkNHKjFg0F7j/Xl4fMbdJQkRIExjDVK0QVzXw7EIuEL6u96Q4SMbgTf+7QjZ2BWp9OndifJ
c5qW0BszX5Y2vGVcdsditeXkWBVc4g6ycjUJ+WVWj8u11NKQaA8vlou77ktKFvFD9119Gcb/NHsM
a9TUi9neteYl+PwTuFOaeNaYDi4rJzBOui9WY+sxf60338PBb0FEaVRbJlvk/7aWn2Q4Zu06O4mn
Jo+UxLETEazqZImASgm1e0Nntlavg09nJS38UsZ/p1fydCEZMOKM3VILTSTW4ikjR2CL4CWoSZWQ
GII1XtgdNJ02e51oCarxTKBVUPbdOVQmymTJJBsmemdBB0ci2hd5HTl2uZaOTXTRnAkOZcyNIl6t
bwfzI69KTvF678LUuGj7WSlgLPWayiPRXAx7VaF4Tli8AZuFssmhPD76aLF0hbV4oBUbr4/VwdLJ
9xdCw2X7ROt9VS6NOaC14uReD2pb3Imjd+ILXp41uwwrffMi2pFUuwSbd5+N4i8gb8SOo//Qafsv
hHL/p1GNs0eKSKwGxhEjVd/GlbnsCZJGS3WK66GwcBXzAXDqn4G5bYIBH4/MgDhdZTMljZkwWwVE
FjvtdAXcnnkTCpCyG0Srzy7oC0MTXDeTxvAtQz3iMRuozyAhF4QEW0vBBWPe/781qPFcUvAVRyVl
XYVof/ephRP/k4GAOt6cD9c0OCqB4NnE4FVvHtQfLgibSKiw0svQlkDFHpLcqDFbGhNaSK8DBRTA
f5XGBgv9QIRQJpYcsdalFu42cO9vMvvZc1zFsPOKNJTox2Y2ogma+kSYF8exj4cW1R9YRchfVi+v
4LKUlpLGxtB8Vy86U+PX/X3c3oDOT7u8G037vQYbvEezQOKP7MpcEJWbK8qHHvFoneMAD+xtUNvc
TWlg7aMqQRkqdOyYfxqrZFgWavbltjDBNOW57ezJI+8puinmPqMASXJGx7K3E0BI6jeg4eWlhkU2
l8C/vtCnGvDlSLrJvdup0KjbQydz92gyT+HFgnYUXO3ZdCN52/smCXQtqO88s6ugntqPKHhl7Gx1
t5xh1msuV/E53HLv56KyXSRJh6LB2gZGbuTZ4LNVmjMRvzGayc0lVlhhTZ0WsbWnReDlspOivhTE
e/7Bzt9zbikG1qS/bdE54eOZ0Ck4CvOC9aJ6+PhfAtC2YJRG03cmYQhht7IE6gH0laFDjs3CRJc1
lhSo+5i0MZCL35Rjm14Y+Dz8DEmFHpA5lb0zHLmugDFhvKX2MrTIkXRtdfTZBWXaVwdz5sckZys0
jE0kB+6cb/7j8Yq/hVoDEjS+1qlNeRaCbfd8+iX+Ytt0gCV4bfdgOS/Lzpt1O+VOXcea2GqegDf6
EyRAAstajKZhpEDNWaeniPvaIRMawx+QtJ4+g0AhyzsXzXiYisLOj+GyCPst2CmcDzx41PF7rE/c
bknzLCrxcslFGeeEg13uGebpSjoTpztLslcQFegZ0CUFDiMLA5E+FJYGxZ4nHciCBSuEmP/l3wDM
EjgHPBxS8w0LA4T2W6Gg55IEh70PA1ermCBx4TsV/SYZn8PH0sJHeto1bkmWrZUY0HkPkfj71kMi
Wtr7oNGLhKs1FYSJ5Lfh4i7WJPeuxHQ2gUdMzqXp4YRQNXKnxdbYxUozeX43k9tv7bFpZUBNez8j
cxoiEimIANL/nNu+hz1q0m6uH77TCTN9gPdjiV9b5nTNDFIrZGX7E+Lmk0Qxn96enj5AuiHfpdP2
+dqIaUMEMZohGVKTAz0BPeRbsak+Mn446jhXKDeaZYdj6YDxkHEoplAyw5CljwJBr2PtyDU6KEjp
Sk3zikuD+a2WDxY6EbNaxDwcnwwZLo7QhVuSc3tKdtLF1gPHwmgrlglF5UOiyOREcYezWHHFxGEv
q23m1YKWQGHZiS5eg+CXJlw48lxUsXSNi+obOZga3hbNO2krW1VCuW3EbFKfHBT3qVPiRtN2ziUz
INKjH9hB0G3KRSTRjbUG1ybSxlhK+cdi50YF1xbwfnMRCxf+u5hD9eEG5xJcJ+Te4cmWvYmZ2FrA
bI3cNvqVHJL8IUDdSaR3yY5LB6i1Byii2pcwrXPKWYtyYWEgYE+qP3lBXXZYtIbQAHuPAFn7iqAd
ULWW8Q8UPSg9BQnrd7kb5W/TRtrcSf2jnIn7uoIR79U8GSxexoPSyxveeVkilbBXAnlg91CHohqd
Odt5p+OSnG7o0vD5Aoaa+nSh+OdBE4y0t9flbkB090ZwJOM8NEYh6JWpxfog8WQOB3KGcg3ERkAo
qtt7yRCEuXt86rdZHSgIzVKcpYj65aGgknE16YZ3riAry0SJBIllARdBL2S3IBPay2VxJi5M5ODH
XIAnm7QO7jLkMRm998LtrOtc5mdnYU6oWYDHduKp/LBwsnRvtqQ2LiWA/OKUwoQISP1/jsXZ65RC
kkxGQs4hNgNKk8jg2sZDr5QrMHghnfEJWf9yFQFWSmq5q5lDndpwECvyJ3CPh9EYV3xTuyWJ027T
UWpwzPc7KHXojwqSDdZdofB+C0AMeYamKJRqV0dbZwN7sJXkNt0OPZc9Hjuf4sDRfxrfl/OP1YKu
+tNgiwIDssy1P3LBHcPQuZqSllInTXMUlfL0yXz0gPOTbtAq5rIdpf8yUd9OhrhBFBsykR1JR4DJ
jIaNUdlTeA/6r49RMTZYox4rJd4/BZDuobkT5L/tiiknhtPetR8BmWXVmZwuRKLLg9s+AnTNiH51
JB3er/bBsTbDb0YU1OZ70NRumUaA/qmNQzTzTfyO4AX7QbBOfcieIvH/MMdry6FnUgU6+m7qwg14
Q6Z2ssME8Nih/28HHhooS0tFp2joTRSON4blIJooLXkA0sw8q8l59uEU0eoa6oilhaimtNVXn583
JwUSWnkX/QwctWNbCg+4RrMMn2hhNXSa7Ra3c14q8gNqrS6I7frHNoAKoRDK/7vIhQ6oMNMJmMdR
0Q7nH3a7v5gtulOiBBRRaR4x7s2sJRrHcYXRCnzGszaUgT27vTjedIt8p9BQCOXU2pbmBeBqzkVa
FNAjDd4o383kdn3V1q9+jxRr5QBgGX50621MF5m8xlj+W/nqFNn/gZbCBQw00EqPmA3aHf+7469c
LdxZ3t8Zl90Pb4L6H8YiOzlFTwtobhxCbBPcsvwmT0L4w6XGcshJjM1AXvEK11nD/EHwbpaMgeZz
q0H4a1P23v3Gaw6C4yxDFOmSlAA1wuCjwe66RajtLYoOgbuFWfxSjLXsISuMsLuiumHYVZ/UVDDe
EnS/6ueVn7Eo3dSvsbCbfTB/0hddyAgtdhZRBBCWIh34/ICDcsw5h5DDKUgr1oz1PMk0n25th91n
gbaA7Cr5foHvk2i0xVojkF+ZxYRgvqBL41PHCBEGPwgiTaVBZdAnALbsEYjXxxReEb51slUUMb9Z
uP+Y3LkP2ikgXxQHFKWf2/5NMLH2GKs++pP2sBPM7IbzEU8NEuIF0QAHmd0MqCQZfjGmEZ2y+EoC
ctabf0vLV6+QmlZSB2tXZUExsZd+UnOXMHcJQtcqa/5uHJ3rx5YnoJ4qKjuXUub5toKX+SqsgxB/
x2Tk3+OO2Le+58jG236rhA0Tx2frZ6eXzqXk4iZeJA5IPad6xPsWWOlwOBBEArunKDGs4QrmPQTK
ID/oGHx46fDuR++OLX8znZi/VUJnyDi3DQVvhfuGYLBUJRhBFJdkpFpRJrivfMwuE28TUfvPla7v
5gqa4DoDV6dntuB6d07i9EsIWEh5DRdpIAoB5HS0OREx7fMt4mBNaLKQHTSWZHZgwxXiUUS6XZ5m
9F8YzuX6mfTTbP0daf71MiOScyjZHgsvTBZ/4SphP4pErBFWx+QqWNX6aMyP5LwDGKwNVHBBl2Xr
Dr2Y4Dn/Ad8aHO3nUwLIANN3jjrtUE1xGAQp97RpTWwAEE9r7iaoJNjXFnuasR/XyFQlsbhD1hRa
0e2hAlT5dh+8XeNQH/7zOpLQ58mCnd65RVbY0JVIaChIDbyPpQ9nD7J6HTkiGTYmxswUpFODdJ8/
pj+a6BqBrXn9XBQmXWq5LAo6AzRYSIptgfFQkwgtL9p2iR6vFFMrUM9USO+/bXcJkAwQ9GFx7mJ5
uxRIVNn9kCzrM8LygcZ9+exmGbdE5iWcleRMqLHCfrsQ6feWQlR7SpVlWijq2ltqh9Yn7/wc2cMA
StWHgwlWoT+tZagoQAJx009xduITZuekF0dRap8fPBM51yprb2qphKTOJseKAT0bglxbWtt6nYLr
6caeo3jdG4JqEPHxIrIbWDWPyATKdLc5G2w/4PAsWEhYZM6jXsLT8/yFyR+7d4Vk53kkQGLmWMTE
ld+C5G5o/dSnu2jm7Br6aOBpUF06Z6xeAgHq76DcJSSZAyIRWMqvuuSd3UUx+4m472QGSV2y6e/w
UOREQ5WUOypsbcOkfL7T00kU/625WT8fwO2z2p0uMXSFDb4BORD5gNNmpxC0a1xOlliq9ow9zFBB
GqOK24FihC1LZGqKfTdUGJgz6UviPrAws0WjjpeE/fV8qLP7VQFv7/9mIwmIo2eWaTGlCDfIPQcC
l9EsY0V5rn9YFI58zOrjtNxW2Ewl1sEiVy22Ij8B+RIU/wWt0JYrfzDc8PjYCvokeiPXVR856eYH
C/XOFX9QDpvaUXjcLCLZNMofJo9VTYHbSCx0xUwRLKdESYcCbho4BbKv14xGE/0WDIOz9ajxzRce
Tx9OOpa8VW1miK8bGv/BW5BLmmLEbP9MSvLOkNMb2JLeC9qU0qKhY5fXV/CHbTHjAUvFOVkGvP6N
ek4ybUwTtrPX6hcYYYGERoWR6oSxqiDUPv5AXQFtN5lrHxFs0CipvOY/2xsI3rWBvj3VKwjNSS8r
eO+Em3tw534ZSpF9LBEQudB+hMvhs+3f/K6SqZMNBkYv6NmAyR8+g/tI/ikEczyWfEvw0Vjt8iUm
nMpXJGJ87uuX579yyTKAu1uMpPMOF8qYuLvfL5gbAAOVdpnIlBrX4ngmuswjWctRJ2WqDMcQYH5Z
PJ90UoHq6qJenJ0hhRmSXSa7yvIt/NzcYk2MYr2V5l0sNPMQEUprABhOI+gbNuxnGFlZGV0558zi
QoKTdtQs/rjB5PxGib9IdBsuzaC00NCJaDMQTz4/CkFRhLr/rQVycySQTj53Iu+LcvqvxKoallKj
U+dG9rrDFdbbumjRbeYKSeiQ/RqHen7jgHbBRiMVGsaDi/rc/su5ZtUkeTxR72oItn3JOOsLklTb
FpFUam0sn9NJ5WY+QOvOcESA4gZYjNySYg1oMEmVM0WgZfKmLrprqxvr9CCTStat4RanoHf/BefX
9wzwOCgxLEiME4gB8BYhKKLyIgE0CL/S/rH09nJZiLvpwSdqQlQ9P9j4pU3uB+2fdGCpsfuqiS8L
IraSR5F1/4CUuqiiLAvB6ic5OscWhPq/WMijGFXhC9VICxJA7Sqo+yEOcUCW4nzFxAFWopeMDm4X
QpKHGBWsUfW0FV0hnIT6IlZenSuwUlk2e/yUTWGIBsC5poVhRCZ7m04Grq3LbVbDZXP0Qh44Cdr8
YgKPL2G5tPWsFtQDgvSYMJPmNEWWaxn6BuJLdEWHgeDgINKA8f4CGCRzsOpN6njnELBidu+jZOAI
smOLt+O5iW18NwE++4OKRhAons13WrC2mLavhNTOFPODd+ftuxtV6DhrgJsHJAg1JJ2sOzGPlVoK
vHOrf2Env567TUBruZHVlY3ZEhENIWAaozTQr+rSuYztk/0io2YGT+nmIt77HZGjnuaWif8spD34
ZK6Zq7qNf2v0EmWJ9NYHMBmYSJQO6hUr0JNzX6ZEA+ZTB1PTSjGYtEvTEdL2F5aoo4buKIRkt5+s
Qs2CcbFyTMkyhq3ky06oPVIYaax/G24qppUUiv2gniLtnVv0dq0SK3MLHJPXoxKXXCs2kfATwu0X
TH6IC4hpHQcsU3a/cnXq0bM9NX2prMdyIWDHgyJu19K+GMORbA6qH5LZv3eipoBF9wb4MAIbJNoJ
DNM3Lcz5IYzK+tGUGPCRXZvNXI3XDcaqTKk3zKvAOT2pL2jZiwk0PN9O72tqWsr1LrdLX9P+6Lxf
0+3x2jP1hUwXCznd+WlSRY9BhqLTQ3UEGqogCTKIILSIRKdVCairvkh+9+EcqsSRWc+GRV8HuBsZ
OJS9uhbwOZF/HHc8pHKQPEMKN5+2Mfw0NdqONR4Y7A999N6qMFQEO9COm1+adYPDlI/x/IOLBdNu
BrBSGJTqiSihKRTpPWwdWqBNsLxn1HIZ5NdOUboC/NG3yFQcJD8LNVIXT8G26dgy7WFi0aj0nzYi
5vIt70AJOCc7Lvf95TgWUjqpNhSYiczrZ+eRDDIFbC2U+tSrwUBJVLdPyxETMRuHCaO5XCRht7z2
fdsxzn4a49MoaMLLSpoiQO8V7TEZeh1oEKN83oMJQ7vwpgIS77JyQDOejt/0xMnXIWGw6e2gnlDB
DAtDoUme1x2YMRwO/0BQVqdF3flbe1cGMEK3c/3+SwcVijs/dwoFWSTgJv8XvR/nlHFCejSC1HSR
vDUty2H1/bL1ygm36qxySuJDOt0fGf1mu7u3mqq0U3ISnyAB6lVSnQSyWynqpXHuUQ7aKeg3NPsd
svItod/EUlV5O7IDvSas+fcoTVlZddBpKpFneyUvaCqfBrNWVlgjbOZGB4nNEDl1WNbhH4G0GNDF
tixKXTuDs215klDWan9NK1LzSv+eTuqqKAxCmgJaZl8eDpA+BW9rwJARxquLhW9ZQ6Aptrs+4YBL
UIeEhnh8HsL4hS757j8MKA4vpIgfIb0WzacZAbjGvuTAELQ5Tr1cTecIFB3oAR3RHn9O9XsKgNoc
bAsujTQOIavmAvsqCGG+WzPCPWKvcbNaVlvgo85X9hBmk67DwaxNAxfOeYZp/QHt4ieCU10NiBVx
zf2Hxh5Tw/hJ/s6hs20Nro2RgVYYjEIIIriXfqv0nf60EYsOfjBkPtiEfeNcwd/nLTWS0AQs6KLv
p2bG2gpsQK6SKUvpE5m2X72vfJCevW8rZXc8+UAYUlmjjhHCfVd8VIXBBWTfPi8unbDAaKi1g3OC
6wXpnYq7A4ZJFXpVaqdl4oJ2yPZkye2MrfvChQDwWZGHndttwBRFohVN2VDzifWttk2ul4BkzR5i
qjdAwuRNzjkTTYoEKYUhRRmS/28T3NO2EIpF4a9L42IIiLJWefuMuSoncU75GHmIfbDsm4BJEyDt
VkU8JAbwjKyDC4ZGnXu3khuBeLhoJhARb8V/p/0C9MtbCl/6kXddZ2ctNx0KHv7sLdL9cUR16P7r
imddkyhgX26Oxb5eWJvFK3m8vTu+mZfj6bWvZHQcdg560L+YTr/On08fkYJU+Q0yk8zTBVux88kQ
ldurpRz6n0YH0VmkZcUxIR0eq1+FRzr8lugn6JyXiGYJa1lpccEMb5nZIs+uQR3fPe+vIs4sNTRJ
rRhEfnMLvjDPgaFryrYxBjVxXFREu51quWB4jNpQwXrH3Tio6VXoLjb0/UPynBSPS5+UJKd2L7qU
ogq90p2afFv4+7d5NUMi5Xd1hjMrIF6ptrrhPVCC43h7VYYR3ltsUjIJaQ9n9Sq/lv82QVtps/kD
4AtdWVCopl5TW7jkW9hRA2Aj1QU9V6/L5S1ktBX5h3kBwOXpyTT4b8TyCuJm1rGtGLpmtO1DEyCV
dmJ6MiVYf3hSsezgvIFm9t6CC+s5xu6KzHAnSQoKyv4hLeTitmoYbLLZqs7FXKKsEG7E0nFOpyZU
fyu/3NM7Gtt1CRkWsJAhe9wOd+ZyZx1aUEfD7fsd+pgleuE+VijXJn9LJSMrVtZKwbjVFWWiXLBZ
ykIcLby0YPTRcBYDERlCpPo1clE0lcYgtjlXXG3CE6sfhTobndeZ+fbtIqXyo6dHJ2TRJm7VX6XZ
cPbku0dpQON6ZEPSzJZpSaxyCrlBgQog0ylD48x5xKsCwsCY90tnZhRUbX6nCBHUoEwDKg2BAqJ1
B71hiTZrs4hCdMGE905GvXpgNd38gFRjDoQY6iGt4LEBmby48tZxDAe/CqKJKdhznQMBn3psp8Uc
C2W8H9ZZDbrxLY4OvjrCrxLVc6Gt7DG8b4QxmFhQY/pw8B3NyyhL+2HI16tRCOi9RVnf9FuiiH87
V33xgkHe6QifngRnjXcoEKA+kQX4roLk+ar5ghYSwy7P6k2sPgsUK1bjLeppRyu0/st9M2OR+EeF
c4wnpScaXgB+AaqRvxeFJr+o/of+0pCG5KO5vFiqzmBsTo6nxPu7wXLL9xMZThuHk9h/bc1Nru8k
nFA+4WnMkstIWU6MpNUy0Dr2gE5v+laO/kBcqwIjoa7LeH7vb/fa5oOTpBOFRTGxqizmm3u1qbBF
EgM0GXPk6tfu9rCWSnEOOAvQmfPBDWgaU0IAEwTSeBUgUjcVah6Zw1M7rHM5Rfw1bNbrFB9/94Ya
DUZUFF3+mBYFAtxahQdoBeahEyJi5a5ww4Fxk4GE9TEwEnUiLFw3hD7M5MFhbkjzH8e73UVco9M2
m6U9+4YXc42YZZ6evaXkLu3oY+ysOcbiNTEFGf1GAll1bPuWCyVlRLo5JHMpt2ibP4dCSH9K/0sY
pkDDgI+KMQ6jt9umTgoL1ajSWqwyAfLYnbz8elVLk/VZ7vhhXHuDW9KpQDkfiEn9HfOqvsOWVJXw
ujkUQKtv+Wguk5lFHo+1n7Gsd9gWq4e2JVcmkOuyGxAhcKyGWB+rEZkyPR99edWbwvmzSOuqI9Ma
cAdwrURXwxQbU8qB5adAW0qtF1yQNOTU1/0HeUFkkFv5+eK+g7ns+lZucq+F2ZZkJpb/81EHRYuo
Xrmt9EJIsDeSNzV/shN86WX5I8mxgc7qVnPvrXa/9Wbhzo/jV557vM1vgzz7K7/p6DA3d1OWjK70
Su0sZwQHI0NS8twnYeHjvl2ar9TsJPDMY2f19oLFNUxy5rGS8yYJpselrtuyOi6HU4/pqwhiD9J/
t9m0PKYmecd/EoDzOm7pTPbCouzoidK1QM77HSsleBbDbZQij+dzxo3aUeonFb/SkGmt/OyiaFYi
Im3xcPNFsq93xpBpRbMG7mOiy8NFHcchZzhntzfkvDZLFhHxEwmsptXe+OQOX8evoNchNrVVJgoP
j6SAceTwij8r6f/EIs/MN+OE6SG0uMtKNFyxkShDzJZhsWaH6nOZsoPNM96u3J7hV7lk7Mv7vLpg
GHjAOGImAt7QPAJw60lMDqO7f+qTjciuz1BXTS2JsuoL+R0zreHY18x5T5paQq7vOPFTf2ecGNCi
xC/5gdkuM5Pcs/GZ0ldA9NxXg7KcaiAky8p7PrrHAPl8O7Q513QggLnWPutNEqQ86aufP1ueJZox
kSmtAx/rkXQepGbZbJZv9hi+FVlD/G1YHVPrNFfX6NkyIqo4ciBqgd1CTjOfhW8HFcWcuw+lbkTv
XRsMzAZu7VdR91SiLdIZEwq7MvDt4nyURp3j8URORC3MgjWUZV9l5IRntfbzwGxmcUIOkjr6eFoG
kJ6Vwc6hifYLG2V9VY/rE50OJYUC4eXSy8tVyI/w8Xe+T511ui7xrdCcy/Q51XO2+aUKdIee0bMI
dSwunG97VW2/kD4R9gn7YralXWwJ2vXhpXdQrZKnPrUBz7EMKgOvyjxe7UAnxZYtgNCtj+WAqySa
s4Vq3ERFTRqyLjNaHo3OSYS3awfQdWUMdU9+3gozj5dNip2xajAvX4rB3jSbtvar3neSKdea/nmy
pH+Z3ggmh+lRBuQzft33/mcH8TJu3LtXQ5qOUrj5sfuksrAFYooBG3vXo1evleu2WDGl1pZPak3t
GNQ1MgxbpCMCDvAo/n+1xt5SCNs7eurOHh8ZDIASvY+nApZTjnxkhhzR9kStzlIgQYihpKhLwucy
OeR0xgeIfaLRGiMVOwn3bBagz9kbtKlpGaVWgsszqu2ICeDZlgZ2b6/0vC9XsxBrA2Js2WJLdFvp
w43IsLWLw4KGpb3QW3VQGmBuOwzpoSVrbw+MyHk3aJjnKJX4y5eqdiD33SybgvAbPJRUvCHk6CsV
6Wqv81wZzaZWPONesFIveW8WuFQQ2LEcRmemQzzetFn0B+JcSQQ5KTwvUoqw13KNw+EncY7Fo62X
pKUDCR388P+Ea07XfnI+lWxJ0284IZ/ezD/VxBsDomKPuztwQPudcwtO/C9VYI9I50tBcwEW8yGO
Na3ucW6fp1XqX1Mo1yqe3XoHaNna2R9dhJQ3B3KSybaSbt7AUhdxgMCR47L2N17n/MzXRPb5hBka
TV0QGETfix04B80whl/UOAYnmT+YsA7CRfwFwNx+ORo1x49awkC4zdntfmxik99ACY8+AYJ2vQRd
hpKjaFy9NOtwKcgvxT5mTj8/3uL1Kw+cHbpHBCDzxMxJv724o2T8wp5En4wlEn29cY2xaWoel/pw
PfHslOw1pujclRl+2TrMwzRL9AiJ2QKJoXKNa7fsqL5CKgkWv+/N5gliVFprwQFYyuC44mQd5vdY
zEWPAEsf1paB3ZlpUuI0AUb9I53oA1EHlGUBpgjE0DP8o/f9tIqqf/TOPoCyAqg8oKWeR/n0ar5u
/oZHboOTy/18DK1q6vDMgyMN9sq1xtm/uZwrfnDk0/94aHoN+lo9ubZ46ec4OXkPq0Dg2yl4ctAY
Qfknna0wDcioeHDtfxCe6ax4xkclDm9DFKPu1ruLCT9gHwZ0aGDAGjOB0iePQk1z3ChAxTXG+gN+
+pLIz5VbZ6jgpeKa9TjPHlh/Lv0vrSQ1jwhSR0sC/gpOhMsLjpRGgRsZMw5dP7gLMbDrrH8pLyfy
VIKi6d288Gu/jbwEtZvK0lnRjHkOSXZw9CLGjiQjf3L45I4QYPjxR782pC0ckfpqtguv+lNA8M1i
BclzBU9/Cy4qZGkM4mjaxyqA8QZoo2IeEhthkK+8ZuoQrfLn7fVNGuCNyGsJh5h/6oX3UqRHXOmY
CtL7VM2IFwnucwPKZ/mDVz0mpVkegPSRS9FxPzr7UN4hqO276xsg+lNfCTbjxoOXK9x2Of2FxC60
XCOzYlEe+fpZuB8keczTxSwQVeyzpFIzneL2XibGmtLtgeLFvCvO5CSb4a0bcrVT6CMDKhi9pr5v
mnpaE5jEpKM+/73G5kPa1xpgeMSBzexGi9u2YCY3SoFwaLLZwu8+GU1eUZVuAl5KQ3K75xhKPiBo
lLjaA5BIq77RnFg8Hin6doGA9FD/UJn4uWtMUBWFWbDRxjQwGr1rf3LwCXQvriu1PLMCpegMcsnX
Kemysh0XTQ+CYr8ZacwIQiNURmKhLYHNEJj+L1HP8li0UqIscVt1d1NbF1yjsWvre6gp6dokrw+4
DTsC9VrQtkjj0xVZJb4ybzFjIRS17ncyE/BtJa+CcwDUoB+AKi1yb2M2eHltw4qKHhL6dDDVNLqY
g1YQOttqSt4/QIJDADHKb1Cnjn/YidhXhWKJe9CKQ1S+9nbD85lR7vHgXpzgv0oueMaVlKiLmLQD
DcI0Xw8wCqA1h3ZcdwPYYU2uhJOKRiJYMejO+iF1mynOKLUAj/xxXkF3AajqweLsr1aDiBBjrUAS
4TyDej85O+wP1fT21xHFosesd3gYdYYKu0EbMCH4Q0kfIz5qHkrsKmkt9VYLCML173lTYhifnynx
zl7+zfqROz/e6xACS1BV1t65TTu9HCZnfxQAxcZ6O5Y8hiXyr1V6GvTA4ru1bZ9+qI01hjSEdY1G
9fMpOGie46Uz6jJYnMbTfjHSEmDnUbYiJ2YF0StEXTsdeGJooDaJCIZuBRO9svSX7wrZnzn8f/Lc
s4PQ+Jef1Hz3q65i6j2gNAOWXDsk1VQFMa5iyk2MgLNR00SO2VP5IXViJcyCbj+s6b18btRk6pat
UwGL/HQMW+DXQRKmKGbkERLWzLZIaqYhFiyLfVgJMHeX80kLfvwuektifpegjsdScIda2MnGKDBA
BQakhRf0s/dvcykna8iU9WZejA8PY9X7lCCoj5fvhMb+6K2AbQ6NffvDLRRLKDC09u6fc2ao24km
8f0uUMUMRVd2p1CJIhAyiahkKpx+y0/qVYsoBMJndmIM/ozCTX1zACmX4/ECMkfPZIw9f+s40fYO
1ZlalaqknBUjWpDeKfIOCZfLsowHk/+xwsADbXfRX/szYx3yi1ub3LRuD1bwcWt3ztzgqFNCAZpr
TmlTNfXw3J6p4lbwTGqv1CUGLNwXSjKesKmfvxgudKLRSlUUuXoFa2HVVfZzUy+sWpLPFW1rnUIf
igoKg4gbZDAPza5MyRnaXl+CS5wnR2fb57UUyLsg1JN4ug6HNxqhlm2Ojmbc86yOoPfNryn/XwwA
GuQKS6Lks2i9/T//E7bVGwmLpw2/Ss1DGl8VYX4HfiMJv4RVDO3bKPRnzB+mtM7MmcrkhiSFrETg
SAVJzq6RPZwpy8n/nDbgoAhnSdhb8T6jPnpTLisgIpDwDDowXhgvE/RVfjmhQ9ca406XqSrGw400
0s1NrpoykBmtTfKCAnqtf5OZPP//LIFvx0rfSelq5Ag4gjF3dmykgN/6AyqJafA7k9+soYBQBI7V
txT9T8msp0uHVGoG97VA7JwkaZFhq2o8TYV5hMlplDwn0PUzXkbYopW0wbXkZw2cL+NnAH3dg39w
t/B5Jtrbx6VBYb7xT9boo+oQiBaEKFW1gq6MEQefAvBiJwn9asoRwnxUKzoA880Nvn77IuSoluDb
iO3dcs9ZFCQu6ZGyICWj4PUe3n87ocxaowWAmaw9O0d7k2dgRMA/16yZ2QB+qCYG5qmlrV9aDE9x
XTPyS7cGDeCUD36ueYxQQCvy7FqPHGim9z0NjSPpmBSSVp8p/EsfmfYjipsKLz9H0oas02V6KkmY
qe/jIam2cIa3marY9dnKlPtbYojBkuWHcG5ghV4ngUm4zM6oZu9JDGcxt1lgxGiLbBrSyCxgFKXO
nRThjC9sO2wXQwm9SXoMtJX2Km7jGiPZymsLbq00hDzjG+SQlWmFT1dUF567/Ykl4+97800ujaSA
4OHcam8X44kZ6K3+cXQ9DGcT9QgCLAHA1B3PHEsu8zs7+9g0O0RtWARKH9wXidSEm7XdyQBCerKy
BixHwhCPlfM1+9AnCDYAQ39r0TQ2ICIlImNUN4qG6K+nLz13MMRkfQHmb52NmqlBVPzmQpURAoGY
sSV10TXr+tT72+w6jibzL6MdNHypkWVmZelLHFHPHn38+080/AMpp538ZflP2x+b2tIueQ7qzaVZ
9cc2C31PB/TZf5SJQeL7Yxq5VeZkfaZiNJLK7HnVUaL0XSqHOVaOl5M2Y/br+PKrPBs54+2trFzz
fciXdGL6z0C5LJyGm8r/Yl78Mm9tHcoBJBwNlZKLsf92tv/37rGTdzfmp5oRxwgK1Z0x5hhOxsQr
cRJXdT0Eh4VRuk/MyxRt1aUu8N4MIGo+ONMc97dF5G3QJyG7ybCRaGHptmvgeCQxFZ469C6j4V12
kuJlR9/MlqyosWj5WJaTrcFDZBwgUunGsLjLV6HvE8fVqeuA/ZQBUd9ebJvPcpS2CFemx8W6nE6N
hGDWYj4gurQr+Uyq3nmm+7sTnaPEANkUSWYrthCGy4QmabW5FwXpWNMADIdZP7MSZtS6m6Ct7y47
YFPGmGtBvUDzjporXbLVI/WZuy9CN/v+D9HKz9fzkdt8HIDCxA+oYejZnHrmPEep9Cwad9DILfiD
bnKtC0tpW2EK4nR73XWdX3aA2t9OIG5opHPvTK2/fpj1nzaoQ+gLepjgYxXM+2P6sLqB+Yg9j/vD
8IExVotvxvWsN23AUMyG+lvNs0XQ56l+9v8VJ2zkAVR1a1kQSCgNyixqmSVATUTn9gkNKEU19TaA
4Cz70NVvhT07Vmgcj9LbZlsRsEUWws/QpJUvHT8H4scsM1bPGWL4OpSeA8dVIipa38WBzxMfdls9
dyMaXTSAZkDuz3fA7TU/LPXx54yvM3GwGkS5Dc7kvMg1iFkO/b/D1ppRPXtK59U25HmvTLwjdwpR
fOLZfD3fcbOjPCoBznhSn5XeHlqHy2alvXFHdlKnPu3i75ecvxchCiM1nQipS9+CjfsZXQPEL89x
1vcglBpOrO1bcBeaJoH++yBQbEctK+0fv4pTxJ4UZcT6SkgXn3JpUd4nlU3vxnEizEnLHjxMTI5c
3UhHJWtY6RWGGZgslpGoH4lULq0P3zNUDCw5gdJ8X9ITRTQDQJBVyb507c1eQdHLl8GW2i4MnKY6
Zp3xrBGZHlqbULNjo+zOvHWEucn5nk9qexHoezDJSjCW6Epl/FIWqQ9UoxrzpOzcUib2xl0fRtYI
34gS5OFE6qTiBUPbxYljGmqCubtjucNksIlILHcUsCxjMUssBVWSr4pGsx98GTJV5esmCn3lwWfL
BbbkPe1buLx5tdOzrv+fyOiPbXV8Kl9IZ5QWygpw/MmdTtH/XJJhvjAgG3JZW9+mtY0bnKRNFZxE
NVakVXNRFBr5/tV44jgw5u5QoKXJFJdfKzbvtg2goLaIvniqsrcHXxdkLcGSlcmdfxN7/j/uMI07
Npjmpdcb9AuYotvbympSxRsrygZi7OFnTwORmIxtQmugqe+50CjDFHbrwPeWRQbddOVFGr5zmgDd
1VfHOWzzhOnkwiQORZ1DsCD+UXEmzNiLuj8qVDVax4x+k4bkeXM07B+z1OzOYHkNc5OeNXW36e1P
TUsmif7nHkKS5glIWuXmv0DQHJxPr5vJuV8McIUQzrN1eknCIwJKg/pAv/3IUEHVsfxkGPHdBRVq
tG83a83W2cstrShw49PX7TOxLlsWEJi4QQOut7x1/xDgJCjEsQBx3yMgCEkmuHPO3LBSaw6IwVng
R6xL/Lxc0vwOUPiJUf1osUNFDT3BawchSWzmI3hx+M1qoC/ROxEcG9Ax58mH7+hL+06ccvqy9Kyv
sNWkqxOZiRyGE7581X11dPqLIIqI+atymjkF1cLNovLu4i7Xxrq+5hLEyc6tDmQRE/Vio2yMXo2B
ng4BrTz14xM5breNvplcNHSR4wJPLOXUN7XWKIVdA55WHf1G9NHOUaV+/wL02qr06rPPTFWYU1hK
OlNjHtHe4utAj+lG8DBHK4Xd6jfABB0iee0Jc/ZQdmz7YaNlda8U8jMEbDOcIHPe7LzKrsPn4YPQ
7sayzOp94zJDgEQUueyqmjdTle3MW75y7wDwV2U7uW6fbs/ZY13BtQpvATK2rrT3FsLiftm8QsJn
AZUjcN9iMwdh6OZvnOwosLHAbo8EZApQ/gzZVaFc+JERVrCXokxvAp2kcEgUY/pJVddWX59/MLZ1
s5Q3JPNtz62Jutu+iMofvzrM/Ocye7RphmJ2VOStUNHszY0TWtwY9e73XrUBxUM8Je0k9pq1vd+0
d5elQEgalNlGP61MWIwPIYxEMljyD6OQ0bRGZL5ri/S9gO5fruLrb2/CUMayOq65xLXyG8FJN8CK
WesP5L9CiRjr3OUOlJTyBQdiI9/dn+4Me6AAvLCnkUobgIszIvNpQXtz+PLibB6MbzVQ1vEjDUoB
SBCjjCv2gP1J7gEdI4YicHbQVlmkIEnHM+aDzQio2ZEEfvRg22t1mPDqC1LiLp/KtU/Y0i17n8PR
PNB45JLgRWDi8gDO3SqrrkzcKrSurbbisqZ6YIxApTykzAPz32njYctJ2+qaOWv5OBhQ8ww5TgJg
5X2+WKdSlCICmKh4Rt+dXUsdSAfZ7S8RQNqGfQNigoz3sJhWeATLrBB626GdhBrCWMnBNsv5BRhK
u3MXx9pebLifwssp1wq47eVCz4jnpuBBwvV/EMcwj1xgsm0JIpFlOA1olfPvqFgMegCpk2F4YsdI
Bi263HjFq+iU/T+NEXz5LSZCiA2uK5Sm6jM/v5j9WLG0x3z9rFRhKNN+XUoG+A4z5aNdomNojTY0
WA9OBn1j4+/C4AEas551nEWVUb1bMGXPUf/Oei98CYajr+0O1rblWVaWHb2qeOiyo5BerDptGCr7
6fhMiDnvyjyC3x/A71cDinKSy5Ott8V5g6a1NS3j6FnsYlfasI2LVZAUQFKpIPrIMLLl41lVt0XI
Zt4akuBbdeoYJuRzJhgsWWmS0VmKM2OLmJ59+H7AWxqYWWEotFD6emoeYySb+nPsUAk48XIaulnk
eh6oyhLpBRDvuyzYoXCcwjId1bTBsnzNxfn2sDK+JpNNGPWVVMRLAkKegorBoOjc32ddcQCL5DUo
4AvHg53Asq4r75h2wVTlMukQiYf6AsokwlREdeMRIwlCiG3mVoDY6OtIxlz8S2d2ceuhWZCEobop
GasYdw+EoePGOf4gu6lgOT/mcPee+Je33Xd4rARe4vV7O1qiz9NEmrSxbGCqNGDAroNzAdI5QF1H
kbAamom5wrX3AZAVZxw5UepiD5lu1WtFyCwehpCtWm0vywVO1KTtu82lWXzOk22H+8GgtjMZxxIJ
9MOtPcW3HO9mfzaV0riuVGctvH0w5BS8huOBng9B8Acxpnzue35xTRkNOVxrDs2O9prj5b9jSzBv
cOcD2v/i+F3xEUFH3MhEmuiZPM/KY1i0gskRy80dGEIDZx719ci1KgShyxEPdRQ5VX01k++bOFzm
9H7Z3I8zKaxeAGprplXO1Q0WRxlnH/+dzhNfi6794ncWgh4jgRfzQN7Vev9knXzSwJlKi+1BvchG
71XqGNPeGArRfT8ZaAYgSwzS8r+QBcwnk3TyFURKv5ZR7dYO6lTPB6hxve+9JFn70TVUv9UI0JdC
S7G+rMYV1Gzi96YDJfv0s2j+lNPB9w7ip3IlfEOyJD0DfYCzDJHcczQ2h9XppEKjuyxdKJ+3Gj/L
03DqzSOLw8snbOlyU5Uc0jn1Q8z2OztdxiX0gLdwopANd8a0OPmc+46u8oMUZ4ndWDrlLdBx2NHQ
cIgehNoWm0xY0tX6cE5Unun7Fk6lNw4AQr/H5AmYJa9NyIkZMn5TipsI6HBdS7cWqPhP3/3uccOQ
m3tWgzwR0h9CbaSpFATQCPs3rQ8Q8759ILHUxq8qvsHyG5A/PS4sJ1aKKbym79C12pmENo9t63Fo
Pk2stcQDMjcvV5jH8XVroAT9HFOVd9/7sKTJULN/CN9sczybbsKNjZixzDc+iXwQ6yjIrQgIxusM
fo1EV7bOFce/sYG5R3FZG9CR1qI6/t5a2qWizyMES8XqWWxUJM/F2q/7geKBpx2sSq3A4w/aoX94
clufjHFQGgA/RHwxau3qPP93Gn1gVok/1PfOHZ0V5tvrCtLbCDYrVJxkdbAn9wWfFTpbTDXu/2YD
qwwACJdu/Ec+B2j7VqUVe6sG+OE5W2XNGsNqbJUrVBXI8/UoXWSyS8wv3aeuCs0j+7eNfvcBFcNh
B2/mJeKMj0DBftHjwk80hCbAdtqMKTJNmqwOqOgkDtBIhEPiVwRJECKlBTE31qsUaS2ShHbxV+Pt
lXQMnwdEYvYlbAD0ucwxNOYJ6syT01PcCxX3JxFtDTFpMgSX4UUROQNXzHePPNxi1Uv40E7556jq
TUAKw/L6T6L68q7CaAMYyUW2bseys/+qBXGFg0THZi/7+HDQZAzA+zG/cS2yFFGxhapTwXlbHQNb
wYJeA+d2LtBi+PNuz4kIBdE933L1rlFquOW3shm/NXIh75g6+RGGtZXSXXKRM86ACnTtue5DL5dY
FU3r5JqlPjyVuJOdkYHzGm+ZJERzL3IJGrWTk6Ln+MXsbZ6Fc+rRGyDuXyj7msZ3cavgCvwjq3Lf
3YrgPjCBxabBHd9oHaZc7mYntcd/wGyp+Sk0i6PjL4dtLA5yokTp0vjUz6zDP0feIDafGy2oLpaf
LHHEuzDz/BO5dpfdcwYfvs6TpmEKDzQZokuO1RlFEjqs96bpKVUbEliMl2boWmTa7EaV3RxAZzb+
j8E1FLNalhlxvNEvNUvYM6awHuARIyq48PKZ4EAsRLnfG8wyvupuGO2RfDvkgV+HsnXpk9ngQraZ
pWfcwVtZbRyJ++a4drgmJCqUcAxSrTa0mSd/PEC4rdeJffkXFc8eLXLhVR888+o3dOOWzBMOEqCL
a/ybjsd1xFw7WhWnev2PydYZobKqm701CqsPkSKaljwK8SxUuVTLL2Db7ztdMwSBsf9lCbYNnwbD
by7RmU4HspY+VhXwbYJA4lMAqE0V1By3bY8LNAGKMC3imvhE8yCIdDkPbuuWUPOEh5zz8BkqmUAR
lG+Xgv6AbSbYBhln8AW2yogVHJQGBGy9iZIw1FtROlDcgjeWHUVkS3jaBxCCROZ6kumXPgyqXxRo
icqfaPuSGwPcIgkMVb2DNOtLinRGjsj3A328qBDdrWjE004pQnBiuE/k1kaiP9k2pwlKHgB3W1o+
rvX4XRc6yz4tup/cxTm3w1k0vGg/MYpzvg8nfZuISJ9Wmgl2dPw833W5RFViSkzQWm4Oh0usp6Hd
uiYq2rRO+Gqsd+1gqXPbfBBeKlmLmU5QIaV0dZfq/GaHrfv0T36MKCpg61bFMaF8KxmxJafSCIUL
GJJeEIUn9REKYT9nh2Atq7SmLFV4/kEQbpsBtdOHbvxPXR8A2GFWVz/lMoUBVNE2oZsQ6zs+9J3x
tFA4J5h+8Io3/WJD7aDdsAynR5anB08VGdj+JZ/gPVOeq3+1FelwqGoU+hHgNHW2Fu4UwVgUIiiq
uYPWiVNKZ/CYlMlok0xggE4ypribjjMvka0vBJK0DgYkautgXu2dUJuLPqdfnd44ho9qNBZDGB3H
5Iw2iwIW6XGcgBDMA/3jKtJ0Zslx21+/RRCsAjS0C/SLzKxqzddBYjP98AqEhq05gANxwt8U7Mcs
4bo3YPc6F81q8UxGonudMmhVU33GhnTmHs11mCDMXIoq77vbLfhDhBivRWTm5ZkZyOfiVIJam7qV
7WQknQ9BVyLF3zS8iRZ1gZhbDYs1q9i9wqjtFRqknjgFw28dYL67dJMn2fJapABdLTaKsc/5LQVL
udriHSviWJw24GCHbj0VQ7oBmbY4mfghR1X1KyyT2PHwNtJWXNkcM6b5O2U83S+jnX78qt8XtONH
D9NOl+/SptlXZsj65n1U0WP521y/H6OSYmYsee0JWycJcwQgZUj0X9V08RR5OQY5bY+Zxzi615WY
hyV7qedHGycgjmiqnN6qNa9FEyJR0GdsqFQlqZx5HpOQdRDso034CgjfsrUF7krpxldzf8PEi8ZC
cr+59eezos1q1wGTARI7W3zQRVRpg+4svyTjAX20WmhtGgVCvTIyxqp7dwRA8dlxHNFI7yfrdQhJ
1ViRitamOfUzPrkQGgLnW1pKCSmjdlq6uO+jAas89eEdrB6YxRVrSrcJ+XN9uu6X3lUctUg2zsly
iknnloXg2jhIQNcJCyttnSLFmluOitg9oyhWZ94bSAoGzzWjTFuMnjo7w33pXClQDwRZNrtPcgaw
KMIOxlLsubdpseGov26ntf9N1DYzDLIuxmfx7z6uvMZOT7sGJAYocxWjX6s56NUxl1unoKws0RuK
jnezvxc4/j8J+31xQVLi4E/ndj4KYocHea66l8nDQV8k3VsnVUnOZbwrDEnoGt0gR7ZNBiMorpa9
3aGDqTYxajqIEaHRG0ImczlKlW5HrMIcfnpWkiS1jcqBwjyAG0YZl2jmKp7JhhVh7sCdTjutnhiW
+e9fHozMR1KT0FzMgGrdmFzKB3YLXFR+nAQ6tq7+LuFCeFARWkSuM3/NFRGF0ZgY6gIZfG4kQ1Ui
5414SVTg5mdtvlRVy7TMbhr3vIVOAyKqS0yAMLY94042VsEA0Ohn3A6IuYQD1WI71L8OS+TuvCaH
E+bdntspBbWSxXxl3WfRzkbbXkZ12XfuvUaM+SQL4PBhnxdHpIYRhhqRwjG0YiJv5qGP44lBn0eu
/6EuIVEy3eTFSba2ceCHowjcKtnK8qPiaryZSE6TeeAbS0YoJCkxvG4hr52Uqo4Fx5jIDvYKlVDZ
V1Di9OW2DBLCHuc8CrHyoA764WML9I+Co8/CjFpStK4MGe4APKld1V97fLU/ipMzCzj44qhj5z0c
uplYtGxQCRAVJt/KsyUi2hiUg3HZKT5FqGtDFP3fSBDbvmKO+9QE0kiue60tf35n9VBn19fVP2cc
87p2zKq/A9XdWotkByx4pNXrulIDIPynVoxoHBkWb4ih7FRVpXOmX2xj73cp3vnZ/RBndbiSX2va
vU1nYeVgfI7WJ3nGSiwMKZF7hrMC+4nz73dISLH+wCqvrLnqiRao55bZgSUgP+6VZDxE8S/hfMaC
Lsp63jQqbMrGMi7pwahcU0/mGSLcVMDSF0ssKJFxT4jYrkn3sozSQLfsizWEZ6BPknz4+Yxkp/Up
tZqZV99bbwmasDiY462YvwPjfcumarSWUjc5p97FZAJuLOaki8Fy3ppn2mS+lrPKuHtUg81J+Ze1
4/iX8SQ/eFys6Tlw9X0enqWIvVCNIPDz74mNA+4P6pRA8XozqKyLnXfD7Cr2XfFafcY/la1twTlX
6r0Kxt79pBF1LeLmxuprVSdNbsdmKhP11cRE89pkt4XRjhOYcOLO5sjngOVg5ccurOf+s5UT6hO4
Jc67DI9q+Raf15+gxPTC9IE6Egts4Jg8rxCKUhtQjnv5OMaFxN+OEixFCxoAbBGnArt9zagGq5de
Y/n/yvSmi8+LK3z8g3+0bJiprK/tUVIwmHw2TWqmHkgnquvpGw5OCMzp5EZtvGmEZJIl/0AY4MJo
tawPDAySvNQVcYRBlcCuFt9qF8H+U0J2JGNApbbB4zSDtZ2Kduh7hzgQCX/sXtomjstouXGP94Am
FmlRY/Qc9PxwqcOk23lXJjyir1Ed8tq//xOQdZUp7zAPvgfHA53esS7+iRwzJdGykgxigBddDmQN
3yfAehuyfSqmhWQidYHEfQ1aB9+LIrO1quvUazUVNWjwrXHnMm43S/5XBgARbYI3CsZSSxkCmD7k
+Nl/Vr76QwKBDkzc4UYOD4E4ZIMTZz0LlPO6zVHV+Z1z8KJ5Y+lQqwrEd/fRvgQn+G/XFV4ZQBzs
E9sA/UYSx0EDE83vRKtb+oCiFsInp+7WVhn34fyjkFLshp+q3LaJab98D7lZyZ7nrpec2MDeh4dL
Eda5Q7KLzHjHaq7lQoP/wFqzdmFMi/URuJVg/9gOwSACY8Dgft5CSOfhZ3h2urBt2n5RA7ROTEQw
uvpeNbBbDhw41Zt6ZuqMWPtLq+lEulETh+pd9evBewOdJllqpjAtSVbADa3GngclSV/BUggZCBtQ
rwoIHV4UBpBTWeWXNck5GIjTsUnyzvr5aQ7ub+ZdVRWhIZQr782IjngQl//Y0GtDJksxS6SabOYA
fAnfmb4tTdXBdV68kfTlrxeJecraCooY2YWjdCouz0rHG5GT+n1XZn+ZxroUiIAQm1p+IVgP8kaQ
70vXfnqV69zxsZs2bqXUxPzcPHKpTEGVP4z6tFQbhV4bVi0V4WyJ1YmprFP0UfNDW7lV/6p8gsN9
gJqbtkRXD7bRsaTTY1IxPh88EgISZz+Gk4anlRoxZDGQu57NlAAz0xVLhkdJYjqip6IhCaFugZyq
0wEU5o4HozRFMjIr5SIrcdlZzi1V6SqgfJczYuvu+3Exzh+LQ7zPHTIvsq/u88w9wOKmgb/4d4kO
Z8Vw8nyM5UaVZnklI5vYRGtrUe/X3lsaAxIMxKAqpKoxetCWWSfN+OIzJjE79Dk7kvwNyZyhsMhG
CfAUdp50AE8D1KPzD1mNCqmcZG/smaFeSye5U/vTqeF5xoPzwrDYOr4bxlh3w7mBBiSqUAAyUp/n
sP4DcF4+khkqkANy7I36cz4TL0QMtw957N+3Dl/T9brwFIbWBilOCeQ9gSivIkyzPNchoF4Ns97A
v98LGOF9ed2m77OIZ8cbkp3S68rUhawwenlhEk1i3sSsnuMUxlieX3jMmp2USdEhBHcibbIzLyb9
ME+pvvqo+w85jdTvlvIPmTdV6g4HDOI4SF4Fw14s7QG9ATOoWuQCttm3LYjvKPn8xSJhc2idDHr7
Oeku6Lgn5n4pgYvChSOnk8WJm9gqdVN4RiGfTSWU8IsWMAS8HwJuvC67n63W2G6Bu8NfmAJOTS3w
JwEW+dCH2B0jpdmaWvll2fwgFEZGmv88iQ6dEzOdfCksxXv2sdCVU96ZP0jWfBiihmOF5qHH+mwe
6leiQ1ZixEASsZN0I6KIpM9R9qOdOlYX5lLkiP/x1nZhYMcv85PbxP2W5yOT6a11pleX+ODzsBwC
1aSY0uCx8nc5GlUE9WIZ1HAYHbnKUmCDi9NQSHzYMBV+cr1fTcvztr1IX9W342P/DCY7BZdXPl8o
eY7x7DhTd5CBbDYjl5TuUjL3ocFta9O2rx9QzSVIa5XZIcF4oQtsLaeG/0fd4VcZ1MWujZx3YTTu
lwloRn4KG45Mqp7Zv18MLFueKF9Eke9l1D5I2jI8cUyiD0mPRdmGRiQwvn6+tX0zmDzz85Whiy93
YYaB+UZTqY46pNM6rlQpuE3jxod7KmgGN+oLcgEDh/skeq5o275HUy3VEHVvHh9uMwqZvfXia846
ArQoHn8RIENtIaoH62ZJH62ek9fLt10v0DZweaF+oIPV0E/2V8LaqQ6Ih1c/JHlvSYDZtz5uVqzc
XCr0H8AST2I79Uz1r7FrixZg543coPRwOi2PzNFo9yWLVqXo1n8VjFNyztfPb9TTr/Gz/1diLpvQ
wosJokUV8ETLYIFmXZGjg8qfOBi9FiHPWmmYVOo2ewtOcZKrxBZA9RZIGZolqixZFr+P2ZlmHATK
nwPNt7bIgxLV04eKH7VMT74y6TI1zhuwH8XbIsFnPz2WPUeJLFvnHykeSvsynJAsILl6kEX6lIMY
DLBfTAkquv+Kgw15mUgA+INN354s7KLMBnZHPdl+Yv4NJTWBlLm324aAoxDsTPh6BwtoYMg+jYMi
byGlBTG6ZwPGWlZ5Wk2GbbW6u+m54kfZhH6Htll5H7QobpO9iFlsT13O1fRu47XoDAUNrlMVlcCH
cqWzZTwIAMtBDYVFo0VdSh537a5HLw3natitQTqMb2ewNnfBnSMToXqDzo4qbd6gwXyyVskE6vcN
TYoPYRWsL9cIgQt+OMu8LE6cVBVnMC0G/ALVKfsl4FcLzrqid+f6N5yQL5mfqnKP3HjotFegReaa
pGe8fjIfm3wSKMWC3yp2+LB7uZBXtVPk22cbJlfzsq2JgV2cmZXvBhZfO73i3s4MhksSzRNlrU0B
PLr4fEWRB8pEU4oSsVI0XyzBDoMdCzt6ekn5DwzXIUR3WoerRyOkFhTW6v3JzRiGQgAMRHdqDn2s
PwlN6GpbVqz3I8enqHUhOu2m22bJJq+wica+zl1SuzPapAiuSZ6GNJ5jlhTSKbmmD4jDnWV69hal
d+LYsimCqfpN5iLDhBmg2b0euxdkUrZpUnheWgw+LSrx/nPEqeuICD65zmZ775S5Z0i7DS2Z+Ugc
yMG5RzA2B0jElbSoKxN+yzjj6Xo7VkTS9kTpK/+t0kZaTW2ZZ87xdsIqPqQfSQaxc3VJoibN9MZu
iWvPK3r/Vk/9OVArHHKQwchEXYyOjxWMVMrCXJSLgle7dqOZ88JSF3+mlU9kDbub0/pWDRwkrY7q
TkfsEMDI3VzgpcRG3y4ToixPVIM374EfNFYINX1vs2on+FQyJbHvmzCD+qEG5kHVCtI3V1zwkyGE
b5jEp5jIKNJvteXKDALfg3Kf7DtFPXpqYO0Bgj0kPtQt0MKDP5ZECWB3ytJKtN+iMCrLT+mt5XXQ
JjBRnv6831i008NjlPGXmUbQ2Z9K13QPrydsaXJZDgup+akQ+0JN139Kxee8odZUXWJ2qGl4Rn80
2o7eopbNMDfPjJ2UkkkwzJRAL93sHHpQU20jvW/X9xuJlqTp0Od33T1DRvCgRu3yjJ0eX8qiIz5y
uDMPv3jf+vJgmQ7RgBRiE0DxPjUAHwK9X1ruWFLlcgyjMPsBDDCMdfV1KjkdQFsR9+/iwMPgjlXI
tfl0Jszd1uH0mtOoREI78C4GltTJ0HKmTDj/TKZwvhp0TCeptkUsehhGbwJTxoRJ0KQERyt7H6VT
O1ZG5/BPys3L9j190Zjznio2pWJEsLF/gIwGRPTqAT1HIIadENT2IlWeiWXwDRt8iSfPqXO0am5d
PROA9nWvxZFsunwAxIBXdNxniLt/3fTHOTXnt5K6XhwO6sVJiC/RhyfLKGyBjZsd6raBLUK7mQDN
cSHgQR4lzduRfGBar1HGOptTssqPGDxSM+QluptZaArTPWeAu013VCiTPPNT4aSTbgH/2hsanJii
DMV8sjERhRl4sjEqyEDUkVDje3Ehu8KpkU6si/Vxm8TB9YMJJnwOKCVraDgyrA6KW9wQdK8ZE4+I
Bmex2XLp1W0JzAJyOHQJ+iouxOKrCT5ZF11e2G4BaGBwhDT6RAQ6SkzGPdZrGFF89Vj0V4gItww+
APADXcGO/cpawjGG/REFYEIIW6jWq9Tm6Bdys0Ty2HeqiypDN08JNTuzHaAvdIDDlE0OQ5RGWTPd
B0DD89pQ1f/LIbTFRhdTiXNThvV606lLEGi14/qCWQuhMafZheTh/6DXRtIUwQjMzeKEnbqUCrv6
v3eY3iBnGYbB78NQ0cMkGjtXV42HeRpyZpqPFOkStdmEkjgUJ2oth4+7t6XDJu4LktwfZfMA8CfY
KFs14GPc5/I3wE3WYRn3eachsqW212EwdakqoQyBmFG20nu3QnccT7M3jQkN3yH2d39EAKF0GLbd
bVR8RbBzevJbmD4IrNujzvKwWebHw2ypieGFdC3MnBCkwAhOlrKb1hqG+rXBo5UwBcLx5bMINKgX
OwEPGpOiV0DjTfri8xZf6ZW2KdcXveZzmyEymTXXvFp6lzMUK+6s3yluYV9HJzxuNN4d6gqK+479
dZ2Vl9M3BTOEZBeYEoD5fBYuSn8MQhhk/Tk3k31/xZYCYGDtKrwijDYPUUTHdk7Dp5DZaxbg8tkG
AqTuV2Dc+vHLTXlatoZ0a9ELeR+U/kBL1NuBpFNJASp6JD/v1iErvsVT+hYHBqC0uHQepsBGqu8h
NROFGfdqiRRjJGBWyH6+Q9XP8W7LEKerDRwH5gCm0qrEp8PgJiyDAuqISk4SIhEDkQgczhyvPR2a
T67l/v+Gg111TcSrKEzjtIe+bchQgTKbXbOyujJXu+Zj8rHhWw7CmSYJ+eR1spFhhN2LXPdT0/0W
gzAqqbuuX2210PFWSppN5AXOoaM5tRWFCxgBqAdv0EFYQcjg5etKwxge9HwF5UiamF7nZPgP8tEf
tGqBgd13KhPYf9rTGVvCrnbzFeUMtPYM1K5/5sw5gJmIf/1onS+azqOBw7ILfIjDLQWhzESa7CyK
g7rshfShofCcnr6092PxR98ia7LFKAjT7k6IXOfcEH0kLsLpzlv/hNIw0brgFt9WKx1Sq0j8mzRE
5rGPWjOdapMwmtKeLidlRZNWRxwEYF+9i+RKDnTlHxyaFe/fNyYbMFFy12HzctnyQ2fVeae07uU9
AV3Y0Uhy58VI4WBUNZ+1AA2EifI7zJj7TJRZVYHLQ9+6ws56wmTdghJL9Z5CIWt3hYFbqPQmbRk1
lj1btgwib8R7dFYYkeNrQGpiKbTYbYh7Kt3jNEQuznFIfYhRhpsHVEsHq5Jbyzcl8Mh11DDwKfpz
Us3Qg6IsS1RVQ4sps9Hd/IK5gjV9V9ZL/DWvpSg0rhYJT8IrMsU8zbwy3yRudJjAeUeB0RM3QLpx
4/2JqHxUxezxChKLVar96VmdYMxVhu3bcE1UcTE72ifGNzS8crk1niT/MRL8Vg1jSdCkQujPaRPc
XEBvIuCdKxuseGr4DFlX6GVbjbioslbymJnTOA1ARuymRFIPkxRXQdibNQsK2DWaowp23UbnFMw8
AjSEMOo0kwuwsxHThJbgTDAEbp91c6SOP2WKiVwfzeRLpWxSXsFDq+y803wknVA4eodaL4/ird69
evcPEmm+2CIYfFluGfCnzX8Z+Be7kCnGRgiDObvuzkSut8gxH+08G8Mnn1dh9bZgE+V04t/OXE39
KuByz1IFpjC53jU3U0dNZIVz3W66CAYLl9dTJpW6VDiqFdXwnt0xHyGu1CxXiA+LcJaRQiiKflqe
kc6xqIw1laOHiQyDdw7mxXXz1YlKbvZemUCIf0jt6/NtVzWBqPcpJ6uU2oe5q8WUEDbMdiucWvAM
P+2dZPHMISBZ50MSQCYjw/jrGy6Jo2xGag/Ahzzx62fQoXdqc0PeRk1Lo5qecEIFWrXUJ8MLk7r0
5f+zzVSfFNW2PUkVWaS1TyGCzxfVVQEDSgXOsWgq0bwAWR/H5tAFiKvZxm0Y2zLnF4B7qpcZkOo4
rL/tV5mdXySlMlnNqZ2tbMdAGR3NgBBzwMw9e/bwIDQW3BqJM4PeGFOvZDflxUQjxmjLg5nf5Sma
GsgDqq56K1MqYhGac3dZ3PXL1Kg4O9cqKrpbI15BZ3QoApzQS6iqkK3GbPPPSRWdy7yYdEGbzHxE
8QgqyXU9Wfmvj9R0QVgNR6xSResImsTQioN+0e6vlSlgiHZ1+zdn5YdDLq+chrAOi1rXTlWAvOFZ
YwgSz/tqOKxdLRSbKsQINrtyWNX2kIp6jnYxeW3QMX4D+ao0nlJFWaONdQip2KV1vYFY30/5HPMD
b9U/ZfHLWdBQtz3Jzk3gerFT2yZ3W6r760F2BLhpAJedhnrOFemhM9BrTNYhB6U31/BCFczZo/r9
4liuGTdQ/nPtJnHkCgpNskIUfTB4AKhR9std3RA2SH7pnEkA7TJFvgKoRu1329sFVcBFS06ESS6K
0NQwK+NcApgOEUK9Gsrt2xnkf11Bvcll0a1mcYRMaIxJqocDPeMyf0+n3K7LR93mAtQ0P3UU/Jxr
6c7lUhoCLq9tL/ccyFdBp9LSdtbIGmLgBTFPwNvjXl+O6YfDdOhBgWmi4bIsk1SkA0LmbNBhQfCy
dDwb1LiYmVgXHV/j9P51kG+xTwsbObHVguaDpTnDFLQTNT/Ix4gO0MO4Lj+G9CBdFcss4fvKoQ2b
OapdAiAdc6/h5otjuFSKw5QFzTLw1PU0fNNiXTxgEV6PFt6V7RE7FFgmphgSNKiH79ZcU2myd0mx
X7ZI6P4tn0Fl4O7rwdug02YTsUCkASDsIdsxtZm7Gptck4TsJ8CgnojT0Y1qoV4t8OFWYw3hhI7U
Ext969eUYUReykvpUbnpe8NoDCxkRGwpHa3DOLvddU34ekifjqJXOe1amVmeND5cRMT60q8ZzqZw
F18wjN3J5aIhoKn68YM6VZc7mux1LZ89PqVxx1QOQF4wIEI1BfbiNoRarse+9LpduHLU7/or0X5g
zLfQzEpGN0Sf7yogwbAAw64gaMPcrLah9Or/RMa9XGvrCT/gqBzlRwhAR7BXnjfi64uFEPdiQjuo
cEaivTxFx+++gvlGVW8n9Al89Iyb8meRhhItp95dpleJSCDfuZ4d5MI/H1wDN7XX0m/RQj0zpuPy
dulpvIKKLLxdR1G/OhVi6yuHR1pUWxhslBVZKP3naoIIuX0Sa9NZvJenbbCxQ+yymzpVOT+811V7
NFYNClEs8IMVbxXAgOOkxJoqqQ2Pz9pHtgm8rHsa4v3wW1jUbuBqqwC9wFP2wAtbNo5u55Mjg4mg
hczsJn7+LSuwA/hYtz043zcaBtFUoXCnPTTkU1J3ikZ7a9gKP6ANvC+3SRIT6qV9wuQxaHEpmmiY
tegINp2L2hwYza3fdfSeQ+59CMJIY+fUzTGh4g+8cl87kvsb5JlEKxb0kpmqMbE6hRHxsWrisNDC
KhqcpozoNBqE3aTAl/uyxoG8Gsw9NJCeDO+kUZpNjw3pm99leuyWm16+rfL2SLeEiw93UwGsTBJy
QjgYfD41vExrdZAe+Q8qsgACoHTH7mzUAoFiqEfjIwUpczcTl1vzCFEWeKdMzY4dbzI+W6+hvGlp
WBXKrDJ29Nzf60NAe9Zpi62DLNQJdeQhjURIAQol1R/TPiOHCCUPlZN1y6kdj1bPN4+oO+3F1q2Z
tf7n6PsTgaR9ISurJQkf8kUNwf0HZASMyd3QUgfZRNGK9vTqJqJLNZM9iTBMeIm22o8Nad+jVKZz
ggPE5VJyIJw35wXqQEO3d2zM1MZXxyJBSOwNbWw/JfFV1HH7jXfBTZb5LuKPYCISrKBfaWakKYGF
4KgcVpxPtymJ4YdcuDocKdOEu05pnxSehDIDaV8+trjbNxRhWPYgl812RA8EO1aBQdfs+UZ4fw30
SaiQVZ9VExHbmnaa64ZdQe4GP/+x+BOlbvVvsyWS6ENidMbupUGZjJ4aDgGezp1F7kcYOmAskb2k
U4lCbXxQ38M0frc2TLchTJ+0buv2UnDdbCIMYWVs0mz4X9WpbqdQ5sd0vngHX0uO6JWJUHimy4s1
hCt6QCY2M8dqKdcuPhxfHHDLj6glb+GLeeVJfUlneMBUyxmTEhiXMNqDw2anrX+vOnvO4AVZwOdx
i4JHDfmiUZamtS+hCnNny/0tSxeO+0oPs0Pg9ZCG0keWwFgT4vCq1geds1ZjqKDcBaAnHHySdw5w
OOpEeogQvZIouaAns7PFUZMuhupVUoKFt3PELfZtBVYIhEEqSwxXn1uzqbe8XlIZyG7mZ8IXrlLp
KH/ehzAWQVIiyhiSs13EjffZfOx2u9BSuxHRjVj3lVaFPBVkAeglQW0TWqF7PYnLMjys+LQmhcTS
89MKs8bYGVFfDROKHbwW8it2hCetk8VEjD/JSwK03ckSOCzhGe8/ruB2ZKmG7mnYkbwosVKoBptw
80ylXFdvrRgVON9RLRqDqC7aoumstD8TIscluMvjPdIJuj/vcWPQXpQLZvYudz1r4TBPasp6qnnv
/WXZiI0ovDU5716vhBblFtwBXenesX/a4Gl32Z+mTVHik/wmnN2i98lTxQ5usrnyj7rh6bOLUy/e
NeX11bME0f4Ts/svxhUzqHqTyhyD2IuVooQ9om5FqhGarwQ7r5JsnKkyRll6X4+osqilINjK+EjV
n2zkuplGROoOdVWXJbEBvO7Zw3JXbP2CUanhGOFQ4KPEOs6LRiioi7ojF75CwtNP4pkZ0AyVajGY
+7Ey72hp+O7MVNdFSA8ysJ6rSX9oLvux699hoLSS4lrs9iVfam6sQ8a3SLr8vKx6UIHS+s+xwZEB
khyGwMOW+0uF4pESZfLwLbDMQhPTQHPsFkd2TwOrhpvY/yNhV/nJ+wD7+qL5ne8T1e9OsbxQFmrL
JVOl/2RqpZpdNLSMFyeuRkz86d2TAEwq3RGMIa0HdMKsGIXvxwXGasBvDEVT0IL8AV+rj3V5bM4H
9aMLYl/zzgHut4DUEMZ68oPhlA6kYQK1afO0Qrji9wbGuZMUNxCAg033JBcKcOfUrjKWmF2xnFvv
QiMyGvYhCvoGIaDOrEfrYLE84tNnw9ABA3nV4IsLzYbX0BkvmYiOTuhophuAOTIMBssWkLE6eTre
AKEZYCiyPcw1rJcLjQQ7l+OpQOOYKOm6VLRB2EmrmZiL0wuoMXxr74vAb/feJoABLiXrrKYV7tJQ
p2/t6C3A3u5jW3IEEYHsLZvpASPLF1vgP1bgBT6lJb2zp0qCtrtYs0iV1KlXMe/eDhGi6m10rMxr
pupUS0GtW7RDdnI16pp3AEA7YWLpC+ttGbOANNcjrKIzpUkzWPv55dZgbzkpFGLavDFAUkugj0ED
aeD9gvE/JNCecehs/X7ctkHTbl1Za6N2mo49D3tJwFh0CGhUkhPLI286GfegTUy6L9tW2909SNzr
Q9bvDsDkqijGcpW4kbn0sxF+SwWPq5tKn6rSM4k6CnVsYpHyeO2NQC5iuwTQRxdFTC4GSyq9pBZe
tAejOULRVXwoW/naTw9Ir7O4XlLrV9SpXg3bV71PaY/rf6U9aMp5y6xAs5IAi17awT8BqsXnoraJ
HiLDVHp7OgxWWaaLy9AdUh2k1JK0BoukKaADHr4JLpjz4t40iKShuPisxRgYZ74eNriSqzldhDrc
vraulBjCAhDj+3WPDEeNYlse70XMlPOxizVeC+j/66hFAQx3jmuq7GvDVWP8HkYBnYD/UYzczcts
PQaaSaGmyepen2qRpiOIlpxjb88CLfOA3Co+58fBXT2HJE6d37LyfmF8LyelImeqoy0twpRy/1eN
XQwJ7kTY13seWXiA+Rat+kgujMsDabiKFosMz0YZ15lcbc1Ph1xb7EXMCV5S6fyFTZrZsWyKfbum
EjqQri3x2RZaGY1fjxp26lUPjRaD7/dCavCjlw2RABowRJoQ0pRpG8C/80Sa84NoNZeF8kG2eLri
Mhe7VjRjKSkwy2l+FhtS+P43NqcstXlqYHIOCf6YuJRERg4P6tLJikG92+Xx2M/OzVktypo0Pzn5
tjT+yM+ep6sUx5VgCbUFR3TsVwFE9m9sfur9zPt2RBuxVadzJHp8sRzw7hZw54dsWBPS7/sLbIb4
TfQaVvInPkIENbzroIIQj49G6XRRuJvpkX5wXy6T9V7cLj932gLHZsYGRHmt2dSqo/H+iVAL3aAv
9vxluMcoYyVfQI4YRPMTJOw/ITPiwOG/w0CeuAsAA3w1HFIhW9IAhfcZKzZW4WzWfSwtBQ8S+1l8
qZw425tCffZs5kmAUxKp4Q0Z8JsMgOGpJBnuouOz5aqL439hCPKdfnsDRKEZQWWikH3OPOauCp2m
Q5yN07S7nAj0FzH+CuC003eSrk9qmcRtjeLBFovUmBcfwitY+9d2Di1nflkWPA1nBjXh5ZKg7Mhi
mDUhDQO0XzGbZAE7Dtr4Q0ozrub3CeFhakG8F6iQgThZNQBzfQ+BZIojLGDnrPkk45VpGzzCvKX5
rD1iS5KIL5wkJKj/4KHsLh3za710ZiwjPS5GTTiD3Ze3nm/apRiya61r8Jl2KyRNh2a8kayDV6D+
5Q5sBG/3vMpd3M696MswG3aLBTFsXZA+QpUmKJEjB1S6aGale5u07mCDI/pybkdgUG2vzWN4J+EC
fQI1Er7QcOWnL1kBFUvWO6QfU0LsQDuXN+lTIXVqOQKqaDjQXIPAK2SeYLtQcqcVc0UD4KkAbPBR
dVjE4PefhseWIuCrbjxskte/7Q+Lv37l7AY0HrGvJOIc5oPLV4oSgjC6qlOPm7+kDzKcum9c8ogR
E8xt5AAQ0fbxJJL29MOYfFmDQeDYlwEuEUCBFllAzSZSmZa/DMVdRivUQg27iOzI3ONON11NmTAL
2y1V3GCkmEdeT3UiQ5bKoX5Y9DgtdekM0GHDsKxOFyDfTjaILFZ/MW0b+hjMmQpYAKdV9VF4ndqm
+LWF8YYxUbp4xc3odT76rm1WtvSKmQm+zG45dlq2cblng3RhbH/5AoZOEy0ntaYMjjK/RM3VemMz
vTGDrEuUUTJAcu/9uX+d85vQj60x1Q/71OeTGx4AUSn829tY2dyeEaRS4gyi8+eu654aeNpa37tV
RixFC/u7ADeEe7gApdUzBdJeRzNwBJcRESj32ubajRgj+uip8hG+sV2t2WfVlN0oOg6Vvpki/Q4L
MPAxvjHcYQDeJFGHFu+vGRVnSwS97Hd42Re+r8HQ0Zj/NKS0lxiSHgWkazOhZrEdmJKG083koeNA
LB04r5Krc+/BbkGey/873+ES/ulxbH5tsaOyjk+3yUXvNyqFbBqWk+stB77sy+B9nbX+Eafvg0p0
fNS2lwVYFRaBExk7nc78A8fJhfKR5oifFBcWnIvUFhrrCaoeyWzMfkoA7bCI871MILm+Pn4podjE
m0VQzj7ExAfMqic+YVrO1hnjJtfGunBmP3aHVR868KoGzZQI2XZAXO/+pC9iBZqWBtUIkMWGnZhp
ZiA0QFASZyiRALaypQaWx6m7YFNBZjM/XBWikMTJO4dwtpauNZqQtTTn3u1qSgHYVyM+wvSdhDAi
ZA8KPuImjrSUrceVEM8rK3pZH4kNtwE0OcWy4NJ0VOYeHVHo73wkWDvCswGT5hUc20QoIqNLrH8+
YlKMBjTqFe824nDPLulRnUE5FOPv+dGFzy56a11IL1PVeb2/JbkTQGRMqwdt9/0TNOzi5Y+DI9pp
5ARyqPkqFLe+fV5YijkLpIHYL/iGDcV4El795+X4LP20nz8T4h3oaLb65oeC6W9ytp+pLyFQNH8T
BfDUPLVKc/LO/bR9B34B7ziAgxxVWyYgYMmxNKg7kbYMwVSEaEVSvxor4ALh2GXxsxKXJ7gL1VyO
RmQlhGAXRoYLbFrByCWdJxxTYcIa+vRPLvXCYvJo0NVwmsFkyFgytaK/N89kQR9Dyk7esAyOMW2B
7SMTKq/6SOcsm3YoWVNPzL6dmdHMgmXsOvQKu17YzhYQ/cGRepfapQAy8hoKtWXHh4p7LMzTbeFl
RXZul8+6genGDsMTqA6aHEKqBQViIY++K4HdL17AV+U78cXzxwNqNvLR6jOmvgNjaFZxVrcXQrpn
fe19pnTeXwv+zoaX5zEWHNryNHW0bkhHMat9pykpU80BsDZDRs/Asr6uqy2baFKYlO56C6LEI5Ke
4im0O9W1zTDJMLa0IcyHjTAVVpL44Fp0o0H0OCSSU1ZEros0UCpUouKgW3XB0GdqSrfgqI9R7CEJ
/BUvRvDmPH3yw5TyjHvoGTKRVXAUkr1Ux/vqe1Ezz8KkKfz4+2350xcnD4JA49txulWk6kmBwhC6
jKlK33RkQ3vy3dOIHqPFRir40BC1s2EDU0GE0Tq4deZYbb19wfslD0Mv4D03i97wg5WLkTd//sVd
ymHbKbHiwaCfl+nDZ2BhPFAl5KYAUU3nltkfQlOV3gxDPfqtiFMOLhrpDTUCqPFgTWvnl7CXmbC3
Eunm9qfk55SNnbz0tsGtHNzb7lrCSj8Ifn1SEFcH8sbbIOyMXC5WR2P235jkFvItMYGH6tqv5HkK
k62WW4d2o87g1WYQKCahtuYSMUuYaF6BX/bK0V2nnaESSxmNCc6S4Z1aKDx8IhntYKKOh5G1JwJ2
maxxiTOA0TeEOU2XKIZlrQpqjGjPXWabSdrWrHFSrljaYXGRsztFwpkE5q20LtGyXynGhbPWKAay
7c+oOE1/47YOkKV9p09WbPnDPUHi1N2UXrIUQur/Ctzww/6ybbBy04LXbGUQH+bxPVYAuE/6DSdD
IxrALQasB0Q40miNARDlFZQftgaOxWudn9q1CZYt1FT9JELu1IWzs3sSU2mgGPo/qZ/guEKO12IX
0GKi4gf35IBbYEe1Bc+c4q1FJWOScd6dTnxAkHPU3C0IMKusxfxVkkJ8cly9BJFgAGPDCM4WdN2p
c1u67L2zwPbENVWMK6FLHYJlKagRxpuBl/zj58UQmQcx7+YooUm4NZOZ21k/7fnW6oLYvVhs/33h
FCf25/A0fQ7iRrosAlb7UaDVZc21Pz2V4r7CLfOeBLGMZgHHrAMg1KKDkGCZD/+fwW4Ln6ZjzR6c
n2kzr64nAypjev190Vd0BVDYhJA1YvGLWc32QXqAbuMkQdSVL2v/rcWU8ZD14DX6DKWZ/auGbFmG
4RILWwE+MKQIDUS/4LpFmqd5nuZ33SCiRh0ul70nepMzVduDEJdhhzkqbIv1bYPNs1Gwt1qibIi4
y1RPXjqXO4m3LxEJdAhAtRrsBUCI6e9V9ldXX91NxBfv3FyPDZ+JsMuHtONHWckHOclX8yVWh1gR
5cvEIjsu9dIEyer4yDfqF518+iksADadFjCp10L4V53T78ojeCoJw1pWfxEhVtqVCBDTdFIldEUs
6crXcWyH9EezP0YRi47ydwqKRbJBLSe+4a/T9xqbg7bf5rp+mrLl2DmM/Ql+uen0oImu+1hCNu5c
ovaQsPABqCSHfBQJDNf5WvNzmIdllG3LetoLuaNKLP9iaoNEhn0u2wea+udybzPEUtBUEwf6DDua
on6MC/nyEPtMxXhIkNgd/rhlvFV9RpiwnBPWIlEfX3JuArxqgHBMKDVQ7+j2CgpTzCNX8N7T57z1
7Lsc9Z6lWR0auOOBAqxqobjZ67SXSzaKs3l3/z8wj35p/xMTlZ4dx2Fe5QLHayFBbSDeyMhUQ3bp
/Ztv/nL5BEeK1S5h+1axlkli1i49/2StWweKehG8rHvRSGi8QmjJ3ySW4YpaYKbU8wYu0iFgVaJ3
gQ4irxWmuhr+mlf9fNlayo4yESirsZ4cpyUEnVAJ9pyuBJJpAFGRNt7KRdNclsXoAuk//FWzYxhQ
4TZXlnv1q1JEavvW83BEB6GZ5yssF1S0hb7RA3N296ZoJJDVcc1Ca601tgc/GWEXzPC6+abwexlW
NzPNxBdJiypmoGHDOkL0ypIMq+uxcInNvIIkYZSmnohhyQKWLiEabeBnYbAVr/wARt5FFs7XqdrO
PjEkpoc3E/nvD/Kbw2bEAqPXBIbLsheKNWt6d4mJdoDv+BwQQ1V5l/mowtAvZGibolXj5LJD5MSL
qEvrDSPbDhJO0UbZ7bSP7lpqGYXhiZqHvBzOJ6KZmuGU6aJ+vDHQhawg9Nq6GvUkhBb5UexZABTd
MgldYUyo5bochA7AsBbQbqnslOYllpNu2m1IZqFpNhcAgV18CxVxrcsLzpLe5ZAGzMAE6NXCe3jH
XIISfb8e2vVLybBeWFRmlhnWMewRlTaXAoPvMUkpkTsgjQSZJAC48ruemG6K+CiPgbDx+O2zmgye
wa+R1y5E7NdOijkhU8D05NUPpk0Cj2RMPiZkY8oFSsDWNp/h1R6eDXBbnwRFqztyjU0YvkcSsjjC
GxneKGtYtoRn9Wk7cI2pvXIv0+iyBMsAhYRI0Ytx5BwvWa/d8fwV81wPMYLyPiohYbrKcLtwKJsA
AwM4hpClFLK1z7mYrvZQS5QEocn3eYB1ibzbpF1w/9VdjQq7hEz9PdF3t7UMfq+X6KzLNAq20eO2
rAm1kMe7NsF/gmPSJmT4cuzJ5nwaQVJvRzQfPUQefnJvV7wErtXsvwvEvupRjfbeQoEePITOOhej
VpdpwIsyUYIrPAXifoENr2BcDhtpPsxdACtslPaZMSMaQUGYZf5UKHGT6bxxnUxoWQEUTaaJlhEr
+A+cweTeY4/XgBlHjaHr43cyLmCAxWZ5sit7llUzA01PRAQ5BOn/fjW9MbMGVwOOCg6d9ow1EFhp
R0SqUcT7HnuvJyBPePaw009d3KPH1eAsNQf1e/T9oP2qVznicTmutbePPn4nevqdW6HKMYFAHsPg
SZZygWgn2mlxUJYbrpiiOq7KkkvBsJnaWNmqhwf+o3YxRaHi7A6UbBtH4R/eSBeAxxbG7LuomhBh
9zxFT9eufrAnY8u466UnMLaceWDdOWTTRS4TBHk0g6lNaXJxSoXZzt3ZZor8HjWx2GaM5RjnaLXQ
uCmIZOfL4VpdZ851q9k8BMJcNrNt5m55RUg0sFsK//FpBd7fypKHOjis544elA8UDnd0oKihYInO
s+yl37rvkKj82alZJrmvn7rX1sXXfqIjRcaQyD2du9ukrUyMiIuW2BcsNpq9UsbDjMr15FEKfHhK
MX93bdgTh+uuVVkcEFo3hFgz7e0Heovx/AziBrFNIV4AaKEQ4CSb4KSm3XyRWBMn6Vj9fdh8w8JC
bdhKdWbzz/Lwqcd6rV5DZvZYGwNdwS5pD28AqS0yVWq+rgZ9r3m/XL6uC3WBJctKK3/ZM7zMOtbp
yqk2rfDi6EGZF+sswEGk3EXJqgSxyTJJVO88egeEd0atYrk0UMrujHiNp59q32nocJZeot467qeH
4R3GAw1RQkFF59HaVM8S67mjJIgSkgcEohCTxpcN5RR+6PKSsWpKJudFHAyLorb4qiHpQ1GK61IZ
Ad7bNTTNfRFHZyF83E0lldy5XdqcvHDHmjh3GDGib+/3fxqcJOLm9BUhHXNSAdZyOmp7JYDW8dHz
uRvQ44h0W6KrKV2vTi6YrUaKcCbVf5+LcGVnb3lR8VNWGsvshLNnunnu3UJIXWn1fcqa/LyDnE20
YAes9wF1GXZc5ctp6od6D0brj8tr42WqODCuHszRUxtiU8NN6gqprjxq2ynSvLGouGeklsFTnESV
OQ6Z7Ek4Snw/ZIJWBiqC2q0oS9d36Q05SRERvftId8UqG947LbtWBNLtO4aAEyCWjZnNfRYsx0bB
Gd4n249+FJCmkE3yT/XhlxTedZknxL32/n/Pku2LNFZLAatZO5eQ1JvrSgazaJmLAd5pD7hY8XKN
DNr4KXQQc2di5vQmksJ7d9YJNIim8OZAyfEB27Yr9s7IU+nuUAyGlyZsdwJRjKY050t+lF3Vz1FC
6sYbglDgny7zl40amcgSDQwtEcX/wdVmN7e8+MhleuVSqrqA91YSj8pXSbWXOiTXk51S/ADqAJrC
w5YZPKwffpC7PDDz3LT8HuTeu+/zckAYCncSZR4nqtRIYLpbInc1/JxnXY7Be93mIBla3rMnjC2l
lpmL3XDYudOsJrhH/Jh7Hj075/QJsRAFh6YNcdGo4sGkuhexd2Mpa/5hlDPmSQG04sZFqubn01oS
BQQ3DHaE3g/7c+e05zpwqJA2MnKi/u80PlL/LS3basm9AD4qrDCVhvzUacXookWeiOL1r3kwIeI1
NfpAZOC+dZHoLVV8PvkPHzZvv7NYBBXylZOFKHrq+GOoJlof1DiNGWyxDtpMFxUAmnQEYiNryxaq
5jc52J2QwCSY52mCNDcFlqngeZDDmKIJsBgWXEKg1KwDE0A4eyTpkPWmiI+HjlZjvfMjnSdl2SvP
AnRuAdciAN++GfVP6MpcuV/LZNkW6Emx0iCC9ZKpvmIxAiFmffORkRrH2zJJM+mkIBMGYHIwqtlS
RLAjYzX8QWq0t8hiqIC/5MhPeHzKZof63LeoPwQXhVfObirBvLMG3Sq02vjfj8/w4b1DYbpBq4YS
+94wNkHmJXFdmUVK7r6o0HbbKY41i7Rv0wWzyIZzO5TI7PjJgilP/t7O9ITFFv7IqTTd22BHIxMQ
jOIzYAlvqJ6GRO0lkb+mi8z2mXlU4t+mAyXUa9myhXa66m74bcC7I+PRNRATShkW4O3EVXcXRDBu
yJI+hEK8ynAIO6tVkb4sT/uFCgiI7QPUjXJY3w3OE3vPtu6hjQeF3UQGpGYRIDKJyYygT9i3xnUu
j8uLVLC1/8Yad/l3KWJb5QyCcKejXam1yd4u2N+w0frD584XXCabJMhHAHH/m6jZIeciJtI/qPh3
5fKIGQqEwNrYu7FZxbZSZuDLMAwbE6r/BcsGbNb50C7ztBR6IHBMYcGrX6jZ/SuygrWIkgr6bRVf
J491BidPkmm2Dh2gzGRTkCHXoZA6XrDmknVIzWTQ2paBxAu64auefbCOjYeCBWTbWqLQU+9bMkU5
b7QKpoe0X0l9D2sHa/dJRgBNYS4OBtRKc/MIQhx2OYWVrAxOuU2EYQTe9h7891tN1aqUZzpf3zI0
FGhHyfqH+vMVqrwTvZpP8PB9EQYaLfncCfRXpH7gxjFgA2D1kQBJ7dSAGAesKArvjQ+/ta44Cm/s
P0R/fxBwWDdYwS8t1t8afoV4j57rNPXzuMaIk8NYzfAutK3gBvkuPv/hv9iBiRB6uWDoXjQ6uei9
R+BlFpfwimOBf37gKgfHqDHYKtq+b//KkfSoaUD5V4E9QzGRbTJgdjojxNC/RT3f/S4w54bSXRRJ
Sx4ph40aFhtIhy8iyKP4L+NF2pQvcCdEnDIrvq3yZnPX4STO/Q5QZjmvTDn8TCZXVfS/CuUgV6KD
rrLHdmogFBbUpqmvHqeOyAVphIJic3/24AACsoIQZOGkFe+6qf0QhNYNhSZhWUYaEKv7tzoONGit
Gu459ISV0EpAHC38Fjva6evaqF+kp3pIey9sHs2SFrItYkpsTIox+6S7hIWG+5zfUhjy+hFiblDF
KSwI9Bwmt7rKPTqhjRsOE4WEgiag19QwNielZs9o9cAY4Nlm25nw5dHaFsW2DY8UtCaoZd72B9c3
c7CdloRGrIfhOwsyi18LrUQhKfBhHxCJjPO8HM18uDccwMFFOisgFpEjdyjMc90JTGF9O95ISnge
Q5knuEPwmG/z4uFs47mFHJoiSxPXFH/XLsRboMysKajQly43fLPFFV9RBCC71VyJE0TyvyJN9bD+
mmme9k6DTLq3XxkkWXmfp4l5cBKgFU4FqCV6U0ziDJvq1+UbsD25jJmne1VpqF4CYpTlJG9+WQoY
W4CPs3cuWIQhuZ1BJKwpWDmpEsX2R+twbSUMjbPtS9e5meGECy5akgN5VtbeZWc0mN5eO4VDaXQm
dS7YGC8DsCSvH4hsp90Ctn8XUhEU5lEXh1SeY1XnrmbymmjCPEGwLzpfHa0vvgniwuEosdoE/TY6
+NC/3JQfs/ARaUZtwoFW9WMvOaAKLFJ0u+T3xSg1Pw3JYa3261FT2HdNdzH6grJfEVodwkU6tEHu
xEN6ryVWCQicZlq3fjcZWLVhCnCJI6m/BtI7BXB/aGLULVGiUtN/UuDL67NVgA0ZiW6zGJy734Ko
VQ7ThjLhYwjTu+I2VZk1Z+UImmyS9awMZ+fQAdbdw8YxqcRp0v4yeQsEcxcllwG8xKi2uIC7RiTw
jAqHu6EkGYeAhvMdg9Tbc7J/kZPACMWaJ56Wqfn5ni7wpSlxDj7dxd00v7W0wYUKQwVr56H5tnv4
ycZamS5uz4ysrFZAXbJEtyqS2rL26rR7w1pDLIpyedKg1IavH12g8owui3lOPu2F9j8ofFAgy31+
G7pmfNxB7JYZvHfLUZcvbWbzNAdVnqyyQyyL4cX5iQfkYP0ZGD5FDkVumKA/W4tKCnhqLxkPOIAP
OlXlQ1colXN0+O8mlr0CtvFWf/bZOlmqu7SM294dMXsh98lGSWV3aAT7IaBpnpKIXwhh2mfLi1Z5
R6rpehCDXvN0DZRXBF1MwwY24PeDx/H5UaRgR1GjNsoHgUWQ/PJMQpVo17OR7OUyZSRtVt5iDXbh
HR6w4M4v6ABhcc3J/vulz1fwRTTmAke/6ruzeY1zm2wU9BzghTG5/+ArWTJsylNrSZeOBQolFMUT
AEq/lR77C3pvDAMBK65bvvs1TJDrPqiaiHDIaAvhl+oYtLGicqaIv+3H2lMWiz7CCq84rWAjhTlf
8meUEDPvBiwAlVf7PvnK7/iXaMw/CNfz53bqbGTZeLR/6tQ/YRM1UEtbpvyExRzSBVTl8EuFoxlZ
LeArTBjsf/46BTbvRdtIo1NxbtfjhzteXYpcZyP8IvkEe8LfLhENY/MNJhytiyhqQErP21Tj4vxl
YwgwOxqICEnqLiX+yXPPo/a+ddKAOg2uyOG7R34Mg1/rLNOCHHyykE1YKNdDHypB8aHe/jXmEkNe
XnIiLzYLeNmG6P179aTFV+vbNNQRxDi/HuyYIIOLAwySEnSh7DAxLOxqYl7NM/FYq6S4waYie9Kg
nxJDfbeBp1E/UE5d1tgis0p0Mc7jnifS/US3h4tJhzTkbVIlmh3sbMMKdj1tQJpCiD6vV/Qbe8TH
8EcXFY33VCplN1f3KMsQy7IfnznxO6idYPcQ+pQ8UouOJoUL5DECTZiL4sSNlDSn+YGBa7HZ9jbw
h3KZD8F1vq4oeSWiqKH/VI7O/aFE1UdN3w0d7xE6cMUVFuicGccEkblhZMQx0GadbHJLWwwMM1Hz
+ClSNOjSDBgJjGdKSI8JOeJlZArgQNs7czkZWiNCaQcsrW7Zu7ExDy9NFLqc4q7T+ElA4xeCuWQW
Vttb4S3NTGPtFYKYrlFWklSa/CljkZ/+WbwMRZgJGF7rq4BG7dntSE7uwr3fu9r1XReM0zBvu9ii
ka/ifZAyd/OtHmFhg4IWUi06zkgpDiUOWymzauK52jdBDT1jmGsa9g4rxOSS5PeZPc00jxsJPHmM
/c8H5rqIC4e/Njf4uYamhjDR03gZlcapj5Ut+y0NAAOCYsfuXt5RHFjAZffuCZesoo3IJiYfHkVR
KdufYE7MFvP+AWFjkiW7xiwfsc9ivGmbjR1zR+vdHpA8KRqVc0PkHkrqM21k83YlrHbeNXFMBG6c
HZ0/OSJiP5AY7fAbaMkIAIck7a8uL6Sby1dv0xrLnpWPWMl5rFFe7j70KOLmXNNbh9jUA5XxcLgg
uembL+RcifLAqZ/AGm2ZaGqGe2trc5RtO5jx3DivkjouwbUMSoP9UojZIPSFmkEHbHmT4C6fspQW
RwqiwTraCUFGQZoQmK3z7FD9lKInKFaimEL4EaCv/T0Ct7BHO56XCRok3Mdp+CUaum8x4lxgh06k
PC7OUv7pFgL1pCIyT5X7ToJdoec1kRST0Msn/zibkaeY2WvKo0om+iEu8qMoee1a5DN8WqU5u/DU
udkdHDie1AZXrKcaL6bPtQZzJVzNlPN7/1JspfvIZsFb4o+myB/rN0sAY/RkHKTcmYZcT8pLEUPv
PvIjK1PHLIw/NqKDcmnBnh5GbdzxbBZ4I+SC5t7iz1YXpfjveO03p35PLGUVYX+DVGpfnlG8rOti
bUaAIhAQ9CtqU45ek+nicoe+Xj1ITKk6mcHXV409cXFwDsf8F3PQupFvHWN6Pq+u5wxyG/XSvxHF
TP+lVNqL5vU8Hn+SfBTFv5QFJCSf3GdsKP7RZq7G3bNR7pxLmSuDLqMm6KA+RBvJ00e9cZQymaSj
CQI54B+HFcDUBsPvy5O7yRIqAXA2ETiE5qxKMtw6C9P0X+AeOrMjVe6YaT8X8dQMeGBdel9A9l/6
zbkekJrwi0sr13dPYVCufIYl3PFMlKgnkilgkovvz17WEl2uwFrBzcSmd2ViQtFnpwRbC4i1ZhRm
iQyATBEIR3qX6Ds9Zl+mdTmNegVMkSs5e78QjLJOac1hn4TG9VAzUye79yvwnYgtj3uGHQlVRovP
LgMK+eR+FLdcJXJYhyWb30mvHU3Y3yKa7s5l8gDc2YDX/QAZedz6/YjLPIfP5om1GfbnXISAkAV7
zHbFRPI+SenaB6P69xwHeoNXmCsP+5i1TNy5O8wMjaMeU27F28fh5kAZ9uF4T2zIcE/Z1mvMDsBj
+1QltWThNvPOL3+owmp6/dm1mcBVnIUG7vbZ1pgLdyzBR+tAHr2SjDmeu7+caP9DdntL3KCemLX2
8ZBhDitJ0SgKfqohjq0V3ekhTEbFP3JPR4yA/SBms4eCeqPOk3cY4Tc33zIShiPcy0fJOqQwiQqs
mTzJZFg4tmUz1owtN5IhrIDR5SsRbDcExtVdV4KQfWwBHyAEqvlfainO51r4MxJ7ir2Fu2kOS1YC
S2zr45c5OREW2QJN/DYbdfoQUaO2TLy/hJhsh5V/TNOamu1XQLDfiGPuoo+4nJqpm16748YXiGtJ
PyLzBpsD6UPXha35r2WL4A5+LmkJ5xhJr+opwgnPbF+lS4B5um8zLHv+tADltEPO+4tTODVZgHsa
D5WiS/2f3wTQn8z9xBr0tmVJrtp+JO9ALporv9t+/kopgK4qU7dhJLSMUZbKRmDvOtTUpYmkaMGp
lY6GyMRL3ISrCTreoP9fkiGBtacTmz2C+VFj/wHooVB3YFrWtVRZp3hbpOW4QmWUNcpaZVT+ExZP
sGYwKJoXu3uMINpERLq5X3rwH5DZSavBRxAxzcjOzNTm97fkucSLGjKEJGy3IcsOXiGAvq4Irfie
e6OzQvHIPp2pXEjMusO2FA2JC8UeKA0afSHxQGFy+CTz/AyLQ7GdB0XKFh9fq4Y0x47EmLCS3PX9
nVx9xdL+ny1nBJEIN9B50xrDRzTV6Qbeh+9tel6C7zNGE4MgeJfO3g09hlOIhI27ldh9r1DG6zDL
+paGQQRt19Jza9gR0JUQbqGxFcK5FvGSk7yxwO+nocntGF1dd9w4Lk9NA5onQbGdMGta/TDvZSBa
vmHJy8rAl7sHllqOOyLKr2eqkEu00oBWn9nzhwDK+2zJq9fmOqvgqO1UrNvMk3KyMt8eRISdcmZh
/B/m45SOjIW/gQu0mzaDJgnXzimxEFK7aML4eZ0Pe8YVFnFpOifoRk6Pgql7FlFC1igbiXHrK7KR
JdAdlg93YrlcGTd2Tb5+SkE0NQMGKQV1QqIIqGIxFRd/6g5TPPmiagY306ohKvUE+tHfBcD2JNDw
3nOufC/sHw5HUZNsws6K0h8VjrpTm7ff4GWxvAydJGLERk27nSvD8732G4jI4y8h8od4AgLL/Rpo
TzCZHOUJHfgqNPpo4IA4nBHzDiahS1MzsHmKG/DD8X+9qmor4JKOI79IbCmq3shwwTmYiQB+WsS5
5oyZS9RQVX2PHiC0HpgEnYQskh61sSeICWdB+WpkEgoHuS+W5ZCuw+RDWPr7oBlbxVAPfnU552VM
7jBdeBeO3BBx05Yva1OHDMfBuZvdfYQRAEc0Y3Pl2WYsUby0srMum6U0oqaEeTg+uobZUNIE4qAt
0HYXlGvaSUrnWp9YfmcHknXjPpagtuOWBjM5wD/hMpURqR8hNZP+uhPI0Pw8RiOWL4a6g1Vu7H7n
v0u57oeUmI8uAzBE9fp8JcP8KHfQZCK1+qC574qlwzXGPGIXZDnyi9O5ijjxpBfbIulNCitPeOAc
3LIktg+vdS3MSZDiK8EL6aTQNCFU1+GKVppfXa73Azxd5ReObsY3EvZG76Bsp+LNETbqbn/UP87K
CloTJpb8/rWX0cY48YaCaFeFF5Vuiqc8GTyvvrCncM7ikDDq6s4sishb8ZWojpkbSM+Z9KoAWvdM
vfpzkTkCPxEPdlX5RfhmriKgHIJ8vSMcIEH0I0cfca8CyDNfzqyF1QoqylftuHP4rl+Yd+Rt9Elz
1sDESm/1yMzUYYXWeg7N2p0D94Av07uyy4fi0oy/Ygf6zcloZzAFLigyCFs1WCyHz6TInnfV5e3C
/NEnkjXXsgzUSwMHErjQ+342atcFqWB5GezqigaGgVjdO338zjKtJpsfQhngaHj7iuCvinB3R98+
F2iW/BnZzgPga0E5yhKmSRzrpozx/YWoanAZ5yzxW0jaDhleAojAAgeWOowIGOxlAF5tPRzLfB61
lLLbhcQoBFDuwxebFpHQiflFq/avWLhnJ+wxeCEW+utf5Smxm7QNQXwhv8kqvOLdsh8YZKA0m4MH
7FkxM5rocngaSIVQn2ONWGdoPJpIsDpiiBKB8ThLZF25o8Pa21NUfrXppQdV+/Z4u95os254PxvB
kckp9Xw5Ib9wXC3OogKAJhxLyz2Xs5O1PugHd3Zjv+RiLf15b2pnXbAkulZ0fJZd5z14+eDAtrIq
K9hJ2kimxT9q8WbtuVicEnQ68K+m6mRNRHierC2JgLfzL3JJONX6gAYTbEGsrV1lFksTKvPxbJyQ
CrlXjbf3tzSuvc6MCm7cybTiR2jMysly5LzHWh7bpXlLbnuLrP6SitiLLe2TmZMS3tQXqRwHud+p
HkX8XLXnLEFsL0T5g1Ep6Aauy9bPO5TCZlHDtlr0udxrgsfWh/HWKzRcENeCzhBpR/WEItoShefV
STvt4A0IJWs5GTtXAQSoLfhzYtxLA3jsGCVlQleGOcV76LmpMOWOCd7/ArsTjZow7dxlgSJGHQ+S
qhSN/U10Izzwsp7Y8AJ1hjoof1sMRGA8yBWUigmuvfBq6TksLJCVotO090ml6pOBLDLQ9GhNfbCF
N/qia7Qq6ItFzzKgSuHdnj5fb47+n1Hp5Gzsx5Tn5NJlvpzd1p0e2xiTCDH/6tXy2jpFZpoaJBzp
noej3wVQg1wjYBcb21U1t1h06ZZ74ENrABJNKJ1VnS6hVhseXnI7acHX3uQXyimmPb8j79qLH7rH
I2VWnozf83lxDl7s2ESbVZzMuFbXYqn4zVIEapj5UjMUQoTHlogGsh8m9iH/x+DWTHEF/boygdw/
jAQ6hWAHqcVEpeZ6DNBYZAPsOr/uvykKcUxvx5abSjNATzplf189j08hWhsERiVJ1OxW2baA6BME
M0cVj97orwSBt23LkdniiLx8clZA3OXysAEaJGfTQg1AGLWS3NbRq0y1KZd9GhHgiifp48b9hFrM
dX6No4y6asG21+G5r4CE4ciPNSddF27zY+Fy34a0VYQxeYV2Dn+akqikXfXMIGcyZomZWMyB5lwv
9Yb+bjykM1OA+wm391I/5YolQJIADlHS8F7Dwg2MdxYKW6dxnr2LQOb6TLhlKcdgl7CNbhLHrsZd
QbfTVILWIX4Bclk+ZigfeqnkOoHsGemG0/cx+rG8a0QJ1GU3/pBR7aJbZ8wFXhvvEKX0GBlzj07D
ma+CeLc4ARtFMjEP2ROOsLcQptBudLW1gMxJiWUGcy9M1Ng1tRy9R3QtXD6QKqlmfRVZWNN9Qkpj
sAzcJP62OJapyArV6n8q74K3LB6hwAtT+4XYIqO1NQ8gktCrpfN8+4bQHTieuNzpSUMzeFp2hwHH
KoTyZ79ZiGXlP0GgEpsfaqXwkSjgrAIyBqI4BhsI4rwqeqhROz2R0oEzynkQsRK6TEjG1+Ph3XKu
oPoVU5qUH8UKOsxnjJVCP6hHI+tp5lCpq4Kiek8pEFJPR/1sVF0Vcxj9zgdRE9hLNdXUafUa5uVx
Jn/X0EkCb5tnvXgBcUvR/gzN62wV4X5MN3C/UmfS3WFgZG09qwNr9kjheRZhNzSvrErAt0yYkXjb
50sEDP6WWj6DPHundHsk6o62Z14zNJBRRN1+O0OayidcRzAHM4yvbQXNlc4kYrXtregHZyTcvB6v
BIxqdy8NIRriP9ZHe4zos67NlZtoHLO1+N4APmC28viHiB4AiJx8Qk5rYYaYYon81DCFGviJI3Uf
7igIHAsUKCUFwP0D+San2nfaxHSO7UtXKQK1IvQk/fgjb5LmgVYbKNN4qAuT0m+alQnlQIsLW+RB
WSJybh+jk7n2sr5xVt8sriqhJuhQileZeMUT5Ap6FaFn/V0w2LAAvC8wccQMGafmdgKQeeQcAonE
mDsS6e8N48DjDSl4EuZqp+8//X94sRqBsgV6d3GpuC7heTvhWbsKyXwFsn01GGzm5kDPRcx0FqAG
uVQ2jITucqlTycPiaWgvOGKJw/X2lF6llOkvMcDXMXm9pIkYR6S2w4zmh4T0GlSy5oGPVIrcRzRi
qOzPRzN+wnUMyzUFiW5qM+x4Ly5J3xC+kDLgp/oow+Fmgdhs8zwFEb278fYZneBc24WHQudN4hJS
TCBtgv2IAWHm+nc+gl/sMD7lwT7dlwy4wrGYx1GtVfP48gYCI4CwENrbv+ddjE7Ef8IGBS9f7ljl
hIovyI6Eul0PKUumj2KSxpIloOYfZuBRtM/UI7Ft/h4jwNjYDGoRZZ5ncJAM6UMfmvEhlWT9LHBp
ZM7GeKnd9zzsgDQL656kEUZ4/g7bOpsqntApLfjiZ5JPkdGJsyTSDDevYLHEz239kydXyP0LMObS
CJVocS2ZXgpOcVpi7S/WRhZzCsvs7q3W6QJ5Suv84G1rmBG99xqafuQroragrejTIHSyBl/dV7dz
dJwJAiCpp2gSpppLHR3kdblxHzCdopcGeaAKfGVyVVQ+3kPQK4VUCHxbNbrBOdDTTh+Hauth9YCT
D+NbQH73/yC2k8QKWzeDxNLpkOz0T1VLIqNOLRlgF8xuhg9WXQbqwfbrclHKMQPnIv+UKXG7BEJe
hGwxK9WF2bXRmoHbjeVOT4rdshagH/hIhpFgHlUpCuwMpX9G8ojjofhIZHU/iVa+vV/IqwrZwdrx
3HpUmxVTHv07uJabkSYUAMB/1d4HvY28BPftmn+1UbUGV/nAkNNRmEJCs6yBad95RT3wA4DCAP5c
gXCTNT4SFyhEjKPawD2JVtlpyMaUdKHeTwBru1OKnGISuNMltC3MPDCT4gzA1YMHyb0AwSsU00H/
NJxUOcJ0v467dRKlW8ZV+nklN/KnixDyOTDxb9+BJAFL+27OPHp/rWGdKZrUGhPYSONSdADVnbuf
KHts59RzDIeBD0GwPkJWG++8+WCwycDjYatDaTZw3mVFn7YP1PUdGXCC09Z2r+GmTVot4UYk5kSj
gKFBfHh7v0P1OxEI6N9Qv4H2KlQo4kXh8onATCmq062fQzXd2VMiezR+vsavMNsbD1uSMmtjZrCF
FOSSVDItZXGKn2zY1i003FdzfROTRnq/+93ffRY8BGKu8KinJ63o3nnXeyLjoKaGPH+51RtrGNJZ
bWoVavGtSKIHH22KwbY3enBZwWkGmx3oQntTwHOQeG+S6ZOBiJQ0PQbVjoEyHxSHQ+OH4y7ST58a
U5YEAY3T8u2NUVpnbVaMhiNOl+ysvlQkmZdfQ476VDTv1n4Q2jUBvsewNYEuxK0BVqt+I1WB8yeQ
+aeR9ciShS9gYuFIM9kdHCLxkOCtodz2ft7eAkIEwrJxAlaV9Pygvxj+5ECurzXHBU3U1s63RB12
Emx1MaqTJRP76qZQYocgRVJWKyC3VkNeeaacFFD8gbaLR8ujeDlOB+247y/nQo9JoScf2oUkCTza
N7r10mxg58J4PMz6GuriCJUwqFt99nelIYaDB/z4Ww/PmWrNIULqDKjuQVttbaOi31zn3ojKtNOY
/JYI+J67NuCsymoer74gsZUbEowJemvEB7cfNqoabBXBjGLBm+srocNr/FX/6+vE7wW0mJUa7efT
h5R8q0mqzRi9fOvSoVvf2BgzZv7F9gg1csc20Q8wrGsvXd+cuxp2Olgetw542WyGsTq73Nk8yciL
qLrsv8sgtA94yCkZnM4sWhyA2iX7uC8LCICbHfE0pBOxDRqs/LLHBFawIEbgy+W5zbRtNaP1mpPR
VjR0mzUZqUH67HdOL7AdRYa/wLFZ42VlHpAKK00DB4H5v9l8kJAku6yXdj6DOAMA6EvSphib7VX2
mfxRf4yCfsVrQk4DWMhcDut9Ub8b67mEJhDAZuiefSIq60Jlt5ldCbr4vAN+N5SfdKB8O+hoLjyX
ih6hxUGFCikKQ29+pmc2m/9pI3rygZJew09U81PblpfUjNSAYuvQVvdFdLIVYkIugQmqlHujtJsF
YmJLKe0rjdJBcHiDSf0aUtvwdcYU55jz8CAtORb3Yblg9CCkaEYPiJBU6kIT0fzKbB9YYqI4dMUt
7UEEOFpkaJHr2M2it4ytXU+kOoLoEXCCbwWACThqsHKWz3/ToxJuNh4ybKVJ/wfiWTRM/TRPDB+0
Koi6nuwrKawFKV/CExSv0PyetkoSsS/ZY4MmTVROHZ6l0yQnsggJgIcSJNZ2ig03KpZv2mrOU2R0
I+z3RkJqfcMiOx3azsE+z43gQnI1qofsnGMuOLiwpMEuYcYweQUQPoY/gxrPuTabRbCHFPybD/tK
MXX3MrWzDXjKc/s7c2HAB6QR4k5eHdPp3dWG3euNMirnEFzaoHBpxPi4GVatwcNV/emHEq1Y62/+
1I4rrf0mjtG1RUEk3grMkQE7GJoxtNegUYIXBKzewmeGgCqx643UC4M5N/kZTMhYocpDepStcyiU
flP/1sJH051eJygcFfS0gntVpznBOM4mFp+sodIB4Ooum8xCksI+5xUyMsDv9c8cJpDJo6BfosHX
i/xABOsBZ1/2kqTkB+/AKn6aUXiAOSFzar1woyCwABIHEd9EMiQPHq1Cypga9OARpvV4HoXWxJuZ
yfTc2qkqTf8pRsqBYCIE6katTE+leclL2KmzjTZ+KdxGVRN8kzB/YwaXcRRhv+B5FCGnfnjJ31C9
uFuKkda/hhNjUn2dY/KWwPFPLuQGDhOqyv51F69IZOBNEKeVJZaNjiuhOeNjBspLXp+6OOXQoQfd
3PQ+CILVORCIK9JOidiynr8W7dCPK9oJiHRgUBbFQlM0SS+KzhNeCFr3jae9j3wHciB+uO/sDCfS
C9KnATxEH+oCUUBaBDxi+02ghLFEXvQW4lFrNKnQHqu3hmlShWaT6ln2DwDWqnniuHz7siofVyGh
84LqgUyC9kqJgfKxf45CwcN2Zv8scRqCm7bZTbvmpVwrtpNxmsd9OXVG6bYCGvovEZHVyyYE7Wz2
TBKMCQxhETaOPkJ33qeP1bsk8s1q2J/u70ytVw1d6RjCGK4F5lNY5UFkXT05eKvGS/KkuH+vypW8
61eYmU8cJFmTCgRTq4IeuKI2++BGoyfCQL+90XplHLVynaiItvwbLHWLZozOaqBeVS6EyJMFGbGf
5HsZxbLQAgsGJOnZIq1Y2ysNYClbhxA2FaVHfklYCFiJCKAd4R378fQqoVILgP8Zkoa8UpTWZ4p6
KYU+zzBNZSV5d6WPtXfmgYL+BZnQVB0LyqF3b/YZ/7qCuysV0n3o2hd0APjBOGJtUYU2k4Fqwl4B
OzEBw5eafYHMFSLXH2HMs9dUc6dIpzRH89n7r9+fIgXv6bMZ0QsfClGhe8ua/VaquAttpJn22/70
UT+ZUsFVXq8sxxAGzvCcjM1PqLQNATS9nmfrh4SMlrKbDhKFeVflRdTwEyoeyVwZH/k1D5/gzw1g
IG75geKn8xJEofWXzBDEHUsL1f2aGC7osyfaLXCCRjx4bsJgfcTrSdyMN3DyQyuE/GUOfdp87aLP
ouRtcEbBGJ31DCYPbwHQvDZ2Kf9G7Z0CcvtAbyq4vSOCupLOu6QbdEhdjzL8CK1kPOrV81VrM2n/
8hBdbBXPuVyik7D0GBMVgg+4NsmuV3mB8YoUuO85gvcQ3E4RM1wU3K1pIJOGtfcir1JI9eNKQiWH
NeMoxzOTiwIwOofE8XkdGoxb2gs5txVSwoNgcRRJb8BnS/QNNrXzcYAWKWI5J3A/owkLMwn9pKB1
98RgV/HsF13xqUJjeyXdY1SzEgAFajwjdzpCP6z62zlRQJMlnRJyp0JL3N/1WVN1ZfY8wlWMQiW5
MXXjuY4b+LRAWb+dLk61mG4srmRWgpS4rDniH3/yMh5JyoCVhO3g3xaT/y59J3PLqXEmvkv2xLGV
+Ivq8ZmsiXFLLBfBmq9eRHsHqlJowUVlw2r9AMqZnVzYTOMDUfV1CTydAtUaU7cqnXDJG1GhsHAJ
i2iK9KgEnSYsfPvW/vt8gkIfDqlXYymGhruaS49YFySPfLJZL90VWXGTTeAmzdC7beQYa+gEMpJg
wKzf8xUuydNYSKVLot7dtiEBPELbcZLbuZOh36I3861IGa5mVRqYEjXe3xIart+pop4LkCwLiu3z
4bXAz/wNdwZJ9qTYpRwQalOwLZfCEUHJhVqwhNz5Co0ce2ZRA43F//JEeAjqXQsK4Ij7f+qBEbvZ
HFzJWEqUytuaYSSReDx3qTXAs1+jZ+fsNueUVyVUVXDUxY7kwFV8BwK3CcF7LxqC4LkeNu1h/gI+
hZI2KnuLNaqFAa0goN8BQW3iEy5JiM8UhatyCquDppADdFxOnw4Tqv17UVbIHYx1sCuacgWnDoMc
CE1inaSKaxrgSd4yVQbslsAQmdTSdt57o2oSZb9msvx2AREfyPSD1TYSXH3d006F+m0Glmli8dAx
zUM5Di+V0EF82d62KUO6rhopmwAyzoELsZ569ojroSmy/5Yft8k6VBQzhHHUw6YSXPcITbDl3P8f
EJ0G9O1MDXQrNJqCwWYWOe5ZBW0swFgkDki06/VYys3rsDEHl7BKN85llzTBo/cS5lTJGoOVdAdJ
y/VZkOkrJwTuU+S5aE5YcbbHtVnthUcSWiq21fY1Ge4I09Kmdln1jRnLwCYZGF43VUgX9V3G8I+H
u4/Y7syC74A7ic165dTkEQW9FcCJo0QV+6HdizEA9i6MGu3S64DX46x9oSI/xML9/a3+Iae8kwM3
ugQ6IfXAS7EK4tP/y2FTcTklhkCrkZVsO6aKW2krda1V+/4y2qzLiEZqWPf5cWR6WnTXQ+vo2Mhu
UG4tfeSBt2dxyRosTZdhpI1WTAhDjSWdKOuCuCrqtzWUN50RK7H8fGz+Jh6Pi9SdBVH7GfdKms4t
KC6B4bEvsm6ZfSPsCTjTnxTQhHxGICMqMU7MM842cPRSX14ICfkJSO4loqvvVoFpjlHm1sz0IIEi
5Fn6vzX0jZIZq2Ga/EDBVZlChdtG9/ZlU+af359xutZP52sCWCaEl6Gs1W+pUoSP8nx4gdmvIwUP
4T96ar8uprXXnsfwjSL5jyhof20ba323XFdbxqwAXm3lKSV92R6yK16k+W80/A0+wRjegwukon7F
FTWZCPPTprhJWxL/IBFVBEYeBigPRytNdVs4v08UunBb+dku6/ZTBiBgnfMADRkbtDcCAfe4cMvN
jv7JRWR7wV6pPCGV8a2WvD0vChZpg3XLwt6PUfmBzw+oKq/BZtfLvRcga7NTsxnVhIr5IxjXr1XX
EA2cHDiyBxCGdGX2hc1EapyX2Olw4ob4UhWkiY5z6Zzo7RnyeD0z6qxBD4FIBPQh/EWnlHOuxKnd
UYURnbGcm4Nl7dCHCB2eOZQ50hCBkY2QlwpWec8Gqz1doXln9f8Zzk1KS3qf3kB/XGDOmNYwzAld
IMvqoVNqPzdlC5S1ATXfl1jzZmpGiSgug5IfPYHcJ6QoYUg5R0NGCh8tyVQn1k/RCW0pR23y4pYV
BLwgtlTNm3SN+AT9Tfm0W1a+9bT5VVOjI+Z7ppAAmyg68OX5kvqkpyCM2sIbwIU1C3G75/5QQsq+
CTps57QcvH21RfMP5T41+lo2nwDIuCaBmVDD8YB8STcrnED2PbOV3GmKNNMlLQJCXk2OqL0Lpcm1
hjgHmScFYm2okaKlHtNCgrDzYjmQR00rYhj0q/FyLXrpW4pyh9PfVIFm41KgxvHAIOkzd8giwumh
/5ulKis5gB5NZPESgn6kE+R5JHuTdRoZgAiKddTlVjA1+yVPiEdrBA0n7WAWu3o/7XRDHtVLGAuB
z8X6SmLNSumd1dme4gimBjc754xGhi/vo1NxC2ybfuaRDRwKD8BXTRwdFLgC0uH1g2o6ZCrOOD8D
LWiW+0mkbtfNFdUZC/sURzxrOq3SWw8InFrMZbyK7HBWPYEkNt1/DtIgW7nwdkFl8hzHDu15N3hr
Uz4slCOhNv1BCH/xdTUVV4H/gkIfWN2oYqnPKd2wpuIjo5hdQa4dBO4F0tgH4459I9W5QMiWj5Tn
mMOZyeSIcW8on2pGHEHjJm6hlycD3whF9hMrueqhZGK9C8bBPHDVYrNWmIwP/CTalYZ9AUzEIIPI
Z3KuBoI6nqiw1Kguogu031dpApavVDQF/tb7TcjSYuaVL1VO0S4fJLAAuA5zVIHXljziufHv+Q2j
aRv6OCfcZ7uJMjpodnSCudNMXANeZ/J5JtnuJ5AP26IVv0i+y1E+D5KHCk2Fy1UcbnfaW28PLblY
d2ezMNKVlcwtvqB+2TioTk0G/Zq7hCa/97XeB0+0hUSpMg1Gk/NLtFh+AIkmo2NVgqHKJmhnt+lG
8SrpgWreYXfbtgq6TyHu622oEa4D+y3q+VRvp1qpCO1J5nlk/DBeRDn2cldAS7wElfG7l5KqUq48
GKO2kL6OO1kAzFFFDFhL3QnLMA4yvs87HjTl/pys44B7VkIRgHraiJvCM0hDkJdPukR4V5G0Ff94
FZKnKnm5b9VJf3ES5/+Su+lSzyll8Az3Ttzfyqg/XqFywv0SCi05bO5spWCThjuCbikgomRn+Wor
XmwMnCPClAxdbJ7Gge+elZiffDV6JRZ6vQ5sieEie5NpDLIw+cwxA0NXPi/XmZ2rnnn9YlEebMSu
JefbLEiK93poCRtwBBxNrBmA1q0yNBdWzi7A8grX64W2kzOXip57MjCsm3+F/lHF4SvtVsG1FhTH
eZxe9h9z8MLn2INu+O3ijU6bXOnVX3B757IzUrOO732ZKfL+rQuKmmoQ8fVN5wxly+d1DYTXf+Lx
pZXjm64ks3i+7fQsqB8r9N9PdeMl4+UrYp73iIB1tds8+Qt1SM7mKkny1eok2YuBWzWrQ1Sh+N/V
t8n7RFgfuJhYbTJ0NkKEUNYk9ZuZ9araDME8eQvkH8IbjAxwzsh73ojnU5trAQHp/2mkU7QC/mQS
/EY7ELtNp2b6pvfUZ2weOInYln5qqU0j1hGTMCXAj91EdHNFFlJ99uQUXhb0+joY6Pd6SnJW044G
4yl2eVVeifumos3qCQusiNqLbsxsWoOu/7KtV3ZLG9JeT10o3YumYrpXfNOXroBeo9YM35mkjNfY
EkfzdZSYIXryyZTCV0Ctm29j/ZFYSaEXf2dCZHfWclCIG7eMJ3Fj8IZFfSKHyC5GxAVR9kn1CJ8P
4cdDolfgF5nPrHtQBLDUIsQ90XH/iYmK7CPaAETGEXPEvBO1waGPmX73tzIOAI/ce60p5JAK1vXK
owt9RPNkcKMpsfc81PcvJVVh+feWa1bjNyRuM4IEeaPKgnL/CD8LsIbPocqu5tRhut9Z9NU/k3vc
VkH6Fk5zyyXZh05okQKgd4yC84n92Z0MgfIzTAxqyoko8BC1A93lJczNb1yt1GVpmTv5OCn5WCY6
hs9wM9bdo2LhHp6buxKXtiip9JMiBCC766CysckM6RzT0E4lZZjo4AJ7qiLcOUB7VAmHP5Tk2vDS
n6/wXLbsRrbNBvBweNqO/2ZjLASwv8RqikEo/s5bWskito53/2sga1U/A+9kH1ZNREU/91+lTb8o
HyerDFP94NAtgOLTBMSpNxLVoK7/eyYrL7judbkyR8c9g0UC4Qe1z+GMea8wJrC5u3GKmZb1zFWx
4bTOk/nUYNO13nRYQ2n4kfYX+2lM50SOon9+BOt35YFm9i6qI7s/a14nnBiTYTwwedm8cOvw8g3a
PGyQ6tgCSUYmVe4JUVGtedSBVpjwzosa5BdJOS0bJv6F/UDt2a8iEy7ZO2Pnwg6JV6Izs4tOS82r
PW7UG6xxvsfuHcMhPJ9hU5E6ElgwvmiuyvE2rofySN6ZZFALSUcB4jB4/m9tluFLUgttVQDhVwSx
0lEI8eA9JfHnpopm8MKW2soRhOedn+QMQNsbXZqQEMYoJIfQcbA8tv1d40VAhoxv4o5tctYxadiK
EKF0U8IzQYfsmupxfyxXdk3cLRKhIvg47sDs6zYgelEyf/2ISxJju0ANKiKIa5ltOR7XAlMkfGsY
+c8Las9HcCUpOATNK3ZvA9jMJ2IRksNCgoQAlPVRQ9MZDH5pKGByy3x6fEsitF1h+YzsuKxU6uMf
Haq+aSb4j6OdgBtL2bbvxDRUB5FLmdeSWIlfYWI82+12IMSYycWDIhJPdhxUVuXeNTSzreZWtJBn
sQaG440hQb1BegXwbBGdu7JCE9Ogq1DasVWJUyBIjcl9qni7+wFF0qW6loxSrIB9hf6hHpL9O/8r
6L04cngS657CGSJ3d6wd6LjFs/frUmskFre19ipJwt5LIArZOWT7qegBK9uRWxU9M61GjoIECDET
qIIz0kXWJTRlUrGIkA5Bmpy2oMEOOKlrlSKiSdJW/vfJlBv9cStYEB5s50IjxdZHXgS8URCQvYJm
GpqjGy8zrxB82mfOlh+vmZxv7mRghSqPTjoDBXKt37q1vsuqwlybWkyI6rw/w6IT5Lg08WMl8gF6
rJD2uCJ5Ki+d2ER+8iiZMpSVsl9NBGLJlX97zE16k7sQQnxC1pH/4wwyOfovBavRylFYJ8MpY5dz
EqwKSzUWpCsR1Zbc4540nF+XZ5WzEs/ZIv/5W+HPeBFCNDiArVnmzFDC2ADYG2ogXIL5Ya17GzUR
aE3+NZNCXxLtF2bdb44VfSUBmut+Pc0ZH1vqB4tr3IPpg79IYhWc9/mIukItENSO7uSHFmLggLTE
/43mEOsEtfM5bFBXYrJ1xDBN510siUW3fxLk/Uz0ciBFD2XLmQnP171B0Ar6gfH2ojBdD/UrvV7G
TY67PkOUrl0BAU8d0aSGLXiZS0dM57F6OXlcjU6IhKtoj2sL1x0rBFZBztRSHkOTYbi9UbiR+ooV
UjnwuZuIfMRYxP2hANbk4jyCvXrpIjjwOtSfq0TrehjvX+oDloEsA1/Za7v/1y6r97GTVnB4HmOH
ajEn5U3qy5hBshz/2raKxC/Bd3gZUBNFXn6eoyvnAdHAffkYTF7ukqbyFCvomtUQu8q3OlnIzkO6
VwodIPoEOO6UZygP4TjAuKOv1NamYXDaBf+r0DCwPE/Vv+s7N1wgk9dmnTTDihZ0IvMJKqm7sjep
3iJyFjU52jqnXaVIE/6TNon6TSmDgoupIZCZ487VxLOyyJ091XARktOeI9+9iOHNkS18BfTHxTEc
51YagYHCVq8WNbvUBX8+YUPgjrOOw/FVG5zusRvLOrWOacCACGA72rlnYQ691J4KmJHSdUJK1h3o
fp9Kl6InbuFIjCBpkhX3+8Hya9gsCTR9dDtblTS5X+sVnY3QdUaUR2BsLT/Aq1D+r72kaO7u17oR
NDcHFa7u6cW3HvosPrAitLFLBIXiUUnCRu9AHGu87pVn5G3WB6iAC0G/M5z7MfpGGv+9yFqionuy
7obpMOgPN2tbnW9pymHdXaym5tXTCpNNTS3UcYsein0cifdq94/qFVylRznlgferb13fEc4nF36n
jzj/eD0JERMZy6JfvYjDw/ZuD6MwRh88PcPMWxeehtiEHQwUj8KVt98I1EC3hhBoeEYRkvFPkvaT
RefhwyHDvNKvf8FnIRJMUBlDPCuFnN95ovLro1NUAOEGAN9NTdslYq3a8Ro9232FvexFMyXOZn7/
BR0svipI1NCQvVtU/1AyzF/obWZMe9jl3t0lxsT6Y5oe/gLHSTjoArNOgQGMFj5uA33l0shpfAkJ
5eiP8vNhYzcuS2Tx9QfzaQUrZ8iq6COiAfWu5q4R38UZN64Ys0ixZXJb/r+Jd21My8RB2OVNQ6N+
XDWG6O3Woky3jafrFc0HzISdPaJeMe6CpuBklqUsg7ABckmroHHp5Mc1xgeeHBwgu4mHOaGVbnQK
eeuTA20DwpjbtttkIkeepMvlqdNoh2gpVYqlKvB4UQz3wNc5ydcM9+vGG3316rYnRzBbU3VKLFMq
iSJkR5A4ghp4ZDFBptyyk8Y6wzdUg9L/Z+UNv6RjoOvtCZur2Gyms80jMEqn5bLDV+xzZQpAB0Sr
lXYGSSQekOJkMq+lew9Ab43yttD3k4QgXRk1BWoeqtWA3hxMrV9GqZkpnOfJmZFBOzShVErGbEI1
VJhM7u3krS8KwkOUuWOyODAc2h4K6QSesa/4TYLs9KmIiAjDWrSPxYlbL7NSV0r8ynJQp5oiYpYq
YG35fcpLS+Pf20GjqzVAJtxMqMsyvNpgGp1II0+GIn51KN0F+MrcESo6xCYekAdVbYfkCStg30fo
ritcuSh6QxkqQ/tL/StV3tbD/WKVngdvTJ81OSwYqnny8x8lZIlLYm+fhaklRGtJ1pwX48evAKip
3ep5TbkI6fgoHQUPTYPov744tJTUaOP7/aO9e/VYdgAPCm71dhQOuFLezFn+TGYvEuQ3L9IJ+Y7P
Qp87TiqlQlqQWDt7pLC89kxzH1yJ4I1DejIkTilv41+iHFiY70F/05ZIHYnGBdxLdmH/yf+9bb8p
783ItAN8BxtUncAveX7wyHUEJmF1+8PaaFeR30lA2rNs9kC++uUvjNM+c3w5yTt6EnX/IwVf96kk
Xbo1a1VyZ4q/ECjWJzZMj+QptN+R2U4uDYbcsN9hLJ1hl3T9EzocpP/B4N0sP1/d1ITbqYRZwzhL
6cmKqIL4gyNTOzpwnT2NlFsdQn0JebplIkMOb/A4XeKh1di525MKFA067YQqVIbq+W2k47GD9wdN
4FiIFNvptkRSPtmv8+rTV+uRxkmDlJlZB5l1Jet0Tw5R8dl1G66SJnEiZyWDhODhjPI8jprnjF1x
nkBzDG3Y0kc0AouN0AUPc6JTPOxuqAxHuRy+Ll/nQ7bKu3jjqbTnLykNi6YziyJMUS33x2EWE2Jh
A6FD94Yw57RburQqdiZv6vZSQi9zd/xZ6fqh7NC+toNa5A2zNTVMBWcfKYqIUYiNBmDENwzr/+jb
+u2VZT9jVrlzGU2rXVo5FV1i5WfATXhNu52ysYNh0yvk57WA8r/OPaJgdsvUXgMtxc2aHFOpeppC
TR5I8KTcJb56yiGTZ0cn5gaIqg5rHtdnYSBPCZNpCQwpSppSHJNk6JRjjL/uOK2/Wkj2VHuJW9vD
OSmXd/26j2B5zb0grZ9wTl9zwqEC7bVuDSEf+azrlegHWv98ubHczK/FacBFpP1zQbfgmnluTNkP
fTp8tB/me8wRJWrAFoQRnKQ9GEhSSb1iyNMDd/Tcb5fPX1wgic/JNWsqvw7VMelS7tnUHyGPVX9h
G3xWIeuMrpW7OeiQdftpH94m/MK1YqwBIGwDSXfQIH1lJM8M9hFHspbja1cty8CdYcDeTXxDhk0s
UPDInspTmcCFbNXZMDQ7v2vZS5CzLeK+17o2xo9FFx3cISknre7x+BlP39rtit9lk2flcXZnCSRL
M472jiJoNDGdye36x3vquFZPkrMKwlhgZafR5TJayQAAjNihnOSwXLt0UNc+AGH/ZF1vdTayB55r
PPKBqtQiGbMrx1X8pmFqWswTTe74wA8Z2C/198FqNn1FTR5yBk8uM4M89++Hrptfq31b01W0bReb
76r0uYCF7rGcV0/AopJC1tamiL71QpAjNNoUIGzADUPVlb7agUicr0hjngVQkvlqH6i2/zxzNWxT
WlPCqFSymAWysl6qr2nZ+bl1akji1g4lHcoMMs0MC98Rr43WOJQptoqMBi7DySX6RXqto6EIoDwy
34sq86GTA/PeSV/gY9swreUu/wZYzTeVMb0t7n1vQNPo1Bq+n8ZWqH4jX1mEMSjnUE6Wr7hZcnEq
lb+BJeVXbqPO0oxCK1Iy+llFDZc5LLfBjg1Zs1VdHva25fLtoyHswroI0SofwTwLGKXJ8YFMv9l4
hijrFfzpUVtSpVuVUWG9psRN40o/EZ2t6rq8WQkRYXuCw9F8dbhPQsvCGvzMGPIouj8mQvnuTsGJ
kCXTbbyI5xvXbBQL5UIxPHXXYADwm9X03yrEz8/pVt1DeuEOmwZoL8kOfuX7HeXNeNrpKPdgBuN3
+4OhhoIq3CWSIj6WvvQy+8ZMcsCmI7NcZm+WwA6KNvHU4CcAXiZzrIH4g0tYVWk4R7w8l9y8tmWi
+Hat1xNfp5cZZAnen9jEX2Hsl8hSHZAuu2ZjR7RiS0BuTPCiQuCPBfBRp2C50puGM4T0gkxiR5TF
33kswdYTD5lLlyimCgs2cTZmGZLTRNnPPzrMy7zviCX8KpL9W1aZS2sxytxcvy/p3qrA7Bp3cCqQ
S61Khxl0oRDEYOAD6wuhNAeWt/dItQHRAMB1r2U/80jt3wYAnf8Y74jnCaw8XxDSbHmmdFe702yx
A3eXHCIVZn7kYhIl3ECMI13efOiDSiMs791qOXGLukWuDlWE1PerKyf+a3TZIHf0bDq3OfZCWXlY
QbnkBND/rA3Yi4i74xOXDpQjHF6deP18ZRPXQrDmDDm6FeM8o9AjeflRmyLD8Hey2fICBVqYQjJF
06YBsu6eutbhLiwzC95D+1yUi3DFNVBxtjYp1gECjMFFR86YhsJWYJjRWiovDEvtdrv2ixrh6N+K
1OcG2c+P8117AfPU74Cflpn+f3XuuId3LrJP7dQPrRd6M2LsRCiSswgZs+HE5TRZCOsicNoJp/W2
le0bbxdYS+3F3N+a6iVuUU0cKHuroBGEtuPckmP/frPdf2zZl493wtw/PrMr0dAMN+2ZYBU8RBRO
WQq/igAzwbx2a985gXsqI5hMEmoVTdOeQFOlW5QWdbK+AAn501YX4DBGG2d2/G0jeQYOcoA45Jf8
ULlL4JpDaCoSZuFDt1CvRYBM2izjvU0Sf5MYVofN7MbvlgQfpxFtmZwQtNZlG357hc0oSN0uRjTN
oxLjkSWuf35Nsl58llmusrQEEjLMIaXaAd8dO+fS8QfAb0AQPhQDAEa9pzY4eqcLvzTV3nxebUBA
kBy0sMHqNKMjVeIzgRhM7BPx3pYGNrGRrMjoGixlh4zghoNloJ5mcWrecDywEkpqrvGRxw4UvtoN
9ZL9S2FcxokZTKdCJHTfEo0Awyyyjb5mHi5YjuCvgz+cSvUe9CNacdt2Yf2LYiy41Kyndog682qh
PJMS0Ax+lKi+xP6bg/onTkdw+ZvcBXmGTK15pVYeKGcXa7pOag37J/GajB/nekU2I5UBNwg1aVGD
5/FqYFFLFRC1mYo6E8bPjYfvODE7B0SUtNSLBHi5A6O6XwSIYxLn9Rxzij7PHVnCddZTxSWO7PXS
RKZO25TjHOGsFOu7Y0kQChVPGeGod6eMCQXPsobxheKQtsb12SViOotnLx/nUeJX0p6GeZTQZFC6
Vg98Ghzr+13IINztWq8X93UNVAR1K2njToV3eahGKsdo79aivPF8Lexapz6r2xGgE8RN2LwXS5rH
SexFohsqArzLfTqqKD1MXTBfR+X12Swp3PqNgcYMY+TASUcpfxEy1oOquhF0cpU7Wk7rK02UF/94
EwKhjvGU3GJr5wLdDUWW9ztqqKJnjHhNkW11F5agREjlcmhcuIhyj97i0tFLAq6aZBg7mfHvJgvx
UVDXWf7XqQZeoDlEud6aZY7RB5AjrkXA4QcHv2pDAX93CAjV9Cc6YsP+1N0U5f8hFiyZWwhKDPIu
FVHz2A7xtShMkS66Vael3SE7+bdE4WtRhnlApLEAzFH8svehPwy1p86PQ8ZyUMf/8D0ksJtV1zFh
TTqpObi3XhE/B/D6YPewnizFhdsHxBTGLWb0SLaFCFPgSHyMrhQ/CmPC3vxkyXDE6Am1wH0h8eRp
jBU6rml5TmwE7NitKKEq+y6TujMU8OKv/7a6pfoizcAHGsiEmMhwbARAedTSr+ACcU4Uwq4uahaA
c+2vDL10p+1i5Ot1RDKBj6uW+Ot7uOmyx2o1rXFpupbbPRUXLjZvCxUL/PYucPQdbnub1tauhEpH
UmATI7Y5QD2s5cft2tJBtNb1bkHHSFbDShF5xi1CmLuLgkDfDxlrCyaYLxizTLIIilXVBz/Pu1xO
0ufuFK6veE43cug4VwovOoC2cDD2hgrp3UvDAqsiFbAt+d3vI4oLSNyzkwkPzas4wchxkEGJ/NdE
FqHawbop5KK4+S18z1nB8XV0OC3bxfcxfBWUEKbNTz6k6OhQTT9sgmk+DU8Lfzw2oZByRG11FQZU
OLNwHYfdgrt5GLtpeWrRwIXMxfoxpaz9u1zQREzv4lnug6UoQnmEBNJ76JynV23yDvssvRJLoaZY
eeJj/TfVerNhQPPVqsPU1cvb0TZCWJ01hSVZvhZnYbMxgMHBZVBFPeWPzxOb2h1F1Yj2UpYARR2Q
U7d4v3a7SreEqry3cMO9trxZh7ZRP/roGISBQuFDfropwXy6T7KYqSv8o2zAy88U/YV2lx3qfU+5
cPwKOK146X6tFS6p3SlfE4JhtR6sYoiixVqhrP/LTOGjHXW/yW9pcPuQF9BAx5xLTTgT8/CL9SwB
KY/E5+zXcFsTuNq7ZIvlWu+XRJR6Z9yAOw6DQjAhF7M1Cl74GGlFS9glWw58z9vIKgXkekkrqYIa
FzWRmRPEENQlh/OIdMN+fuNWXg4w2yQOtViMlQOxjBJ2/U6X/xfbjWPybzJzMgDmh7+g6ird0Dvx
NIZ6aU9Ty8ImbOpgqdUs7DVXEYAL4b3ZTRYeKz20saFNCD5LlBgYwBPCIZuX61EKN197336X7YZZ
GoDBGdDJ2L6c9GumbU0Tf9WaFVM1/e8iaEvGDkYKAgJsXlNviRi3itO3RQQfm83tJho7Y2t8l6Qu
MD4xi+pE0OmI8CsBYyNveBFjLq8qII/UTVmF9e9PSOfoMiO+4z0lXIMHCCTGxXcq1MNKbi3iNz02
C/OkfdQ3PrzjMQkT1zyPmrwnyzptOsu9mIKCDIn07zc+8LCGNkUg0Vt3x4rAKG7Dd4jT/aEPEhZR
lstb8R5gfP/StgV0KZ2AGgQc1g8takcpAzj2uqQpRq4sd4t2tdu8Gi+4x+XHmc2+d+ZJT+WzJxMF
vTwwNMOc/Tr6CfvTl5M9qnk51FoXRaxdG3II1EvS4+F5xtW7lxlK8JLe8fAaq4XB1ySXR+/2+Wei
L9Ecip/U07sAm2B1lQvoi06VwtA78CnB3I5QMIpE2Yv7cYuv3G0eW3wICOnz3qEqs1Bz/VvU/4ev
TGxwyrslag0dLChVr/sf9OnCyvBPGNtHa9DYv6P5qC91P1eafuVZrqHmOjqmMD7nFsxuny1/oIll
13XIEaS/vO3szeWTWlbCgysdhpDkMCABwIjlb9+gtJPBOIehpqEOC2hMzmyD9lMmrmr0KChmHhSG
y635ewuryVdFIazGmjfRKzIWmyd9yQS05K2XK1xO0sHyT9e38ffyrTVf1u7vtMKHBPQHC5CKqu69
7qHN5jQ/8LrLncX0fiSNthjneZ9PKHZjuwvkK5YQRgXLySMIBqwGvcMFZFTkZ+m8vC4AYEAIeJrg
YSXbHYYbum3jkhCqTDujQLKVtlXKKbeBswsTh6zyqAURy6JuWRyhWQGBOsGFZtWC12wgocAQFBAR
B9tEWccUR9cFP1KP2IVGC9G7wMGECYxaP2d0LOCFmTT8fCfM6aVia+H0ks1rkR2Ll6chQMZyeiKa
TKNySbhXFALMRvXzhdn2n2OIU6NUd84qoKhildxtgKD9xn7dc+zvRRzxLiq72TxKBokpxULEp+H9
OZ0Df2L6KF0eVytUgTJQdZOi63/fJQS/ZctbhXO56AQ7ZqLrnmU69tbaffMLM6F7yfSHK6BkQQum
avR/Rav38RGrajeUI9kITG/v7zsBKHaqeAfcGKBqwEQGv6OUJq+bJbjACG3dIeNvPlLeyEfiwhsA
9ziQ1Inbt2NsMHmBsmRMuTySXdeTqE9xfnJqSqodsvUpxy8drsAEUkzEV7M5d0YIZOoccAqPKiEa
9N9NwYbwDQ2bWGSFxSTjjAQ+2gSjaXXFEW3BgjnjGnV+4UKAWJB1UJEe7mhBn7F+8nn4NWhrbt7V
sph9B+l5W2cd94L6BoDDdixYKrLEORa+X98V5HprYSDMffKMohDlRvf7CTRM8F5BN8Hi2sIXtT7S
VRZM8kuVm/kyU38C5HMWsVr4uiqMB6y0GBfcGR44sMYoI/RbSngkjbGLEC/q3EkiMs8BiVQe87ff
HLxZHSKzC30tkyD1AE4nmuk21FbaijV8n52ss2tdXaBV8YZX1J59QljB6ixFXa1VjS2x0zKMAQq6
hqQmkZO0hATQdOMORjJ7Tj92kTfH+w0vtX2B42GTOKHk2g4ltezF+osaH2PKJSCCiW+m/+fa4dIL
7c/C3QIatMeA01zNlT+qfxiYBMOVYNjCeW4P/r4O+W4xuX3iVEDIeGiUejc9yJGCChRwYUsjxq8+
C8fkTNIA4kMFfBiA2jvpzJBI8mbYlqkYhRpM9Dvz6W858l7NOJSwXrRTkQslVoUfcRfsIBeese5Y
vN+0ZO/c8zhMJgHgX9KoO/LN9Agq1vDuQtFP2qMY28zMRnzDB+Ic/Bi8Li7s0/lhghXA7qlbtn+O
4Slbz5eqXIsrOWvxVbfihiCy41Jpzh/WIWCrFNy9QJT36xmWhPNht4bVTfC4b66UCiDOR01/px8P
3CS8OvWTuJc7GA+P4YVjznktjertnTGo7zS3zzPkK8ANwQCt/ZXEwkfrn94X7mWOER0ZalwIiLZX
aOT+i7k8Pka5CYSdhpERgstvwWaZejhX4n9CmPzc8DRTUcq9q6jFUip0wD/Zw62ivBLhMIxyLN0m
iblCe+ZDyCyq0DfmYtig57CwPQ+qL6KJvFiQSQivJQTE710xIzYeav/tpYfyRN/TomCSbqf3uKME
Es9p59lPNu1LoaygzLtmsj/rCTw/z8QJ9pTf/6LQcxQqSNqisaag21wIVWQ/GX7KnGB6JQ8CRNTN
CoM7wv6ZnFewRYJtZVJggq7xtBHKUb7dlbMOuhsxV8AsPpN9T2sQw3WP838cGd7SLHwbyjxx/sHl
D+noVebfmx4dp61/FZkrudG513y9HnVGd0o72BLhlQWt09i5yuQe7wZ0Rjx3G1nTLhwMFYbtFREI
WTP7p7+YafJN83pN5ipsdFl+vMvEzoC2aofBqgZA3pxWATs0jf/GiImduTnq3/hglvW3IA3mLMNf
XW8ZqC7/8OqKNt8sU1LPfCtEnkTe1DNVlbr6ifBqyXq4TffhZ2wODOnqrmlGQIL433aAbpGRS5Gk
ga0CBvATODt697MRqaWzpJRFdOEEz58O9+MEREFGjf7j5b6JOEHm68B6dkSX73WTnxdWcQgplJXz
b4cmbn987nY6R6ZRbenM/ZdNerbTsBvXKNUZ0o6K4WMBQPa2g9NxyYn06CTpk51wsAnIhYdPz+4T
WDdrZpQ1BEVvnDi9ldy6dkM2JbLjYpz8YeYqkxuVPBpsXsehmBVXWMkXeXwUec8rTHeYgRI2qTUR
zDIWhBJPHYrbFyXxLRanQfEYLtht65QxMOQfTQo1sOlF+jvlpWqiint95PR9OPX/J+FP1OcDNvKR
Vs3cOwYhDFRjBNleDkGdTRjTavJWdBIGdxFurmP7wFFj6k5eUzCYmgaKwpf/OdcEx159og2o9Y+A
9r3kf+qUdWD02uMNAKn37aQk6pao26Js4bdnxIsR1slZddQusotlCDpdxsTKxRNmOx7QlVG8nB2X
e7S7EYv7SZocRfdAD56AGwVkG2ptkflvZVrXpp9Hhpj1ODJL+LfeHMT4YfQvciqvgaqdYZpfykSF
3p3Fqfq6Su1niA+D+baZDqgEROHt+wqyecaATY+p6XzPD5/Droxv2acseeHL6Kl0oiVYiqhL7BHh
+hDTKFI3iFNmVOdvPd0BIagnrVuNBYc8qhyVeWoSA32TqCjWwLy77RsMoTklDLTYa6DhezNQvX5O
uZOHQbK5gNwm37nphzLT5wHfurSXKiec4nBZTAvWY4FpbF1dAeXZcl5tc4gCN4Q9nt5PAi3wweSq
3mVYWE7EFAV8UYPCi4FM/yNRwUyFoGssHQYGFMLTfv9rHkzXx439Tc1Fu/wbS4DFGNN7jeeda8qB
HvOWrT3CLUfP74Chu5R5ns1pscDH6MO63i3M20LXGkOy4HeP131xDU6z2146sEoz335KlvVodMhr
sfYdNk1Axoptcr2FtBc7x1getfPdsSg1JI1GN5jO7P4QFZ7U9b4uN9naYMEdKzO+lGykC6BkcPN5
I1uVhtKl+Wpe0Lt6heS2lTpF7gtLz3Tf9gF46O5c42Sn7tywOKi0y7+44x1PhIEn/64g8I6YHuwW
bXSj6OYEfWCeaM8qKOFmKVHbHKFA82I9cTzD5eZHitXJQ9zJ9/CSVASMtwQDmu8myTpCggnpHQk6
gP2X2bKomIzGxs3AG2tGU/ahqm6fzWUKQw4oHOkL7IdrgBcC1OuV1qdPgiHBcA5bzMbQ9CyGqinu
U9e52Wz8+vXg4oJ4OEPFkad7lN6qt9o3YkBNOuiKFv+CYgMjko4YKhQGcMQviJchmurgI9OJ1tS0
81XhG2OiMKgvZCKlMFnZPRPkdsA7Vrh7yY+N4j31mAXIml9/GLDvTUlTDcNPRqhKgh6T7wsbwK1o
lVS5rMtYibHKnbLgWUWSeeyfcXGidUcqbvgQ0ebvvc5T64E9TDphSuhOtIab+oIEfZ3xfnBVjRO5
D/g0z7wQW+f/1GNtHI/qivCU40+7YTbEpXmUzp2uHEu7TAq5B0RV4ugG3UL+X6vBp8RZriOzlg+f
koxTE4hn9z0FpbScSSpC1w+TOYRaijWqt72yZNDJ2Y4dsBN9CgRZvqwYQwEmrKTFk8VA0XVdYR8Y
2ZNs731SA0ok9OOwzVX3vTiTHDerI55+E/EobsEfFg/uFxdO2O1RzNGPQDJArtsvFbqxfdysFLsC
H3Cj2l8CdacE7Cz4nQAzNUZnPCyrDMG8ZsKuO1vHuM2Mtw3XFWkIBpv/V9EHGj+ly/pQbDQSsPbm
Yw2DW3VUJS/sM63+aEtiD7+3R0heY437+w6kKB3ox/s3Dpcor0fLyr2hesavCKYxIm2v9jQIqYBB
aunZpp2NBZuF1QppjR8a09EhRMjGwoX5DlA1c1wZxcr66UAfum4PxWYG7vSEguuymgTsvi/vCPKN
SVZIgo8GQxGaIsx7BIFvm1P49Jl2pe3G12/ZVPdh7wWrpG4+Mfeis34J5hUj8MQV4wsLfEQLjg/+
slaP5h4NgKa2LjNZ6jEb0yW4koS09W2tZMDhs+3h/cc+An0ln6kJ8K6RUxGMIpgzwiuEAgu+iW42
GjoSxX4BQaJmfe7G6xoLCdsBz/Va6A+2BCTfSTZ88+zO6jFdojjdJabpbyeC1J5O5fKvVYxIs+g1
qhheKuXt1rtQPTPBzPCcRtWiLPXXXjkdlFykkwvdPb7zhF/Y+ac+Ig+X1z+eQzJuzIGqY5jB9QXB
77VAINGUMy1NAmqBIsKluLIsE3aKgHUAqxUWTWzBkLoznZkpiNXnLVyDS/h3/d87O/CU3GrfmE3Y
rlQc6rc5qJTpTZhlw578D6l9rOjRMrOt7k5e7VS/XDaIMik9vubLb9lVufJHzIrXgj72JVsTA7BC
VpPlhmG06+JngVc1ArTzfAllWUWif7HCx/tb4XG8V5VPEyqCJKrucZZHq9Zgx567LvpXluxKQhfH
y06Cp4l+fFFfKB5NwYoJhB9Jo0GquH0opwpJm7ejAumySC7hNbfc/+zglinwi04Ny6oiI4LNQLIW
QNFJR4pz+twncBUoip23OTEKK/oC+sMDpz00x9bGgupJPAnzDpxedj1ei38LmQ+TbAYlEzD2C8o4
TC4rOpJbk5XldpJyL1k2hqDHOjCr5dtOaOcTQ2aWN6d25BJEfi+TEQrMaPIwP7r5QqF7FV8YSmta
nJCe0eVM9QPHXlRovlfTtntCDFYRQ3hQxuS6yGVYJRLfCvX0CtRh8YAu7s4saiI6Dcr3JN6GS6sd
rdgMHZo0fFLporQGDRqfA9QEmdj0S1ZbIjPNrqtuvF5TQH84l4Nu7vs/up81hWZ1cMLiGeGF0Xfx
9Wt8zDtEhKoSRS5aVFyFMzCW995Wc56ufoZ/Ma/7ILa/p/UOVSgJvuLp0mlBFziIHxFYCHfS6wK0
OoBh8A9+GwTlFsOep3A2rJEQSkJSrpJulvdO8QZbBzXl4di8yoy3J1+0wtW5ZKlRlMfEBgCkMIIp
y3ID6kt6rgXbjDOJc5pIKGXmK1X57JRCl1aisyoR59J2XHWM03N1+7l3pqYtqT8bipapGOHukzkL
gJVAXymOZ8XnsBhjK0HFPpGkWuDh9iKj/VYuhBt7uoXVdf49lmVj9GB6YKfkF/TRvmrgPLlWvSTO
Q3YuXhTzG7n+aGNLonWnluKTbA1fp+6a5ZoBslFVC375tt+bYLgEUNHn7HVILECN4rsB3ll2TfSk
Ect1ExLtn+zrD5uoiCgmGvmjpG7P1/bWFmqaukdSBf1gHcLnflJsPIbXZMzDSl+mvtfXo/wl0Wb7
kSv5TlgUudvI+AodQKzRQ9x3CjrXOwNu1iQHESrEPAtD/PPpprOR/ZESMLGdZGrMyNulm5qdM80G
r1//G8Sxnra02W7XG8Jv3hiCCkg2CLtDSE/nXzkcTq44kfpF1QXGGGMgbyDDE4jptVznNWwd0LOA
7L/K7qc+bi9X76q9tsBJXo8g1Z878ucGCl58+b82ZR8zdvjeif3DikUHPqX5dnzs3I7OppdtvgeI
gbkWBTZzmlLnMH1bazZa4Y6uLHrXOe3QZHjE9A33Mm95rTmhT+3b+A2YiC+LvVJfau1PRrjDRdDo
KnyU5JxuzilyCNtyw8r5go2NbJC16Xdkj+E0/19uULFP/bVMU7IUMIYYNCqb5gUOuB0JHJWP+xjp
ZP/Mr6O4BrSQww205prRfNiadqCzbFzu1c92NO7sBCfC2VzF48BDB+u4WLkbpT9Bt/uy/fJj7cGO
pROrWIw4dDYnymjHuZCDbMONQcm9qW21pFm4yM58HWKxC9hcmTZMGzHP0+ykNegqT3fpQN7pdR4M
qsSzTTSo02TtvZb/ag6+1OWO1zthc6dpBvKFgwg9WRp3//522cqXWgIRdhcx7P6vZ8k7UfbzSxgJ
6f0zIH+FtdKWCdG11P+v3eTyjj4BANTCR43/3qZy/ZsT5Zm3cGZUd86qQfZLqHkx8FkiHc1LGuv2
yNCrQYZZeJKntq6vQ/NYNHFdAyeMhhsCaRVj39QzivR+WqaYSZuNB8rVUOiUxiDE2J9/tPmiIKGB
1XcZ2ier+dTgqQXSN6JmrIaaX6x8zr8E8tfsArq5b1mWf2rbluoO3T5tJ2Q/gYbkzLeoHngnAjtM
cuS2baMe5mLdf50nfTyWiFJiuASUFFQdWdqAINQHEcbusLlmckkfc5H2sL/0CapYTE4+oiaD6ZJT
mJZ6lRdZ43/1ZRabf9R0WObfPzEKOqOjUSvdatbHBla2ItaI3QVuz6GSxIhowrsTJNTevTqHg5Eu
0PWOqYKA2z0oT/wA2giruVIBX55HhaZCUhbON0hdaGOYeYdKnzPGBEZSBTLdKWQyqJFit6+LUi1j
kOFRRPRbKSZPpfBrRlxwB5rPYa5ye8lHyh2mQ8wi/uvsTjLKOCQlRQ/dEw1Jkb3rQgNBawdjQ2Rl
b07V5RGWMN0FzEerS7J91wt6dJFj+tYnNwdxeU6wWMdZQ7vwNo3cRYEwvj22o1tU71ARWfQiGCti
t970b3FssEDPnLSVsZrIt5pJFp5s8V9kHojnLTh3l11eEQHPOib0Sb+jVXprrJzneGF6ih7PUawN
kZi/rCcYOyaHhB+2z8vZCwqGNwDGyXAnjyw3WeeWvu90MwEt1h0zyrx0R3SfVFwECWTB6PCi6CtA
oNSk4P21rVOHW3Dsq1luBVGFEjlYh2U7xJ4Lgv95I6thR5i073jDRB3B/jmunCSiqphwhdRhswdg
iJMDLFP2hvqnfrvBTZHxFAFGez3WbTBxUhCsQotSImE051USKHqu4QpkGu5nPAgRA97Zh9FocKY2
6sm2RXsA3iiYyeRmJ47vh/iKunyW0zq8YrI/F3K/DWup16SItqa4kdaaomU8byBc7xDSMEnaBq9J
/4vKT71IjYxlgeTEwokPD4OlWiNdjzWZzFd2vo5bUMXQlYNX/as+0tQ/xf6CbxcFexVDFLdeX0VA
qA2qlvWcqOorWqFe5lr1G+tE4WpPwCqVgeDui/nXoKh/uIDbT7zqnGvy8WlLJKoWF/YBaQtH75c/
Uvs3wwzy7UPNWMpp+OE1u0zxFM0F5ArYTOE+vEHkwl5o/l6sgrsnzNKsPazl125Uj48Vu7a1pnGN
1LlRci8jctO9SpNDXfwT95AwIlLe/2Zs5pJeNg414cIg7lzpIcIvx6d7m1Zp0T1B2ygXqoRYNIQW
/aA+Z3cX3a3nE0oK6pCOpkxFgOPbc+sxQgChh8djWQuQzant+xQh/6NfJm3z1oTjwVZwx4PLVdPF
qoRwst5B9BRXnKRKGchrBbWikhJWFSVDUqyAoHkK1kzWSn3TH7YSqdbF/VcnxiRJRqqhd3ABBxhw
KaYrNGQksIlc73jSFVBGN4v1y5VsUPlYRroHf2WVl3cjVgslje52r+UXJcE6JbVcoazgPJCR12C8
CEsNRpyNZ03MK1PHARaVp1aY5vW/udVK+i2DmUzGorZO4uZtrAO03haIWEJKLFmCDbb7WWMfrUgA
E/6gAGYNUDLFACQ/9jtm2v94GBsmNo1yULXirxZxlExLeKqypqjkreESbPC6LGuELxdwqwjzWUXV
KAMFcTO68G5pKAEln7p62ZztD0YKlY0rOy2oMATHreRnys2nenENQzfSo0wk2zzVFzSk1HNJ0Dq0
e9D6//l3CRD/J56dHyvqO8RW+FWVnF5qvxIR7ICvfHtYbVt9ulms+4ghkW/olZz78SDkRgU/4+TK
yz6wE4pBT+e13UDUn8T3pkcT9B3HTLSFB9VNTzV+62CwaSSX92Ran5bq6k9zZohviPmCcfsN+hDZ
Jskk9QL4oNdtF/NX9+9S2WxrY8/ZzNOLgHCf264/qnpTLaTAld8eV7TW76dahAgoXxZfq+1AzBVg
f3qJ2MVqfnqoBNEja4vu9O2nNtlvgB3sfpGGJREgrxIypzIJ8pwvYV7W0+WpeEggA7XCRYUqYPd8
w3iGlWKCLsfSrk/jCVbyrFfXDS7n5RI0AVGRnSDuC5j6Tm1Jx/MR974IHPBL9yVHM7DB049dHNS/
mmuSy0D1bZ0JJbKmc3vGEetlwing07U7m5KAed9E7+sr1ME90usCBnF+W1hJJVDTqL4SARrvI7RZ
DNf1kZNt6yrk3GVVyU3BQqUtYXgOS8U8MZKbxVKQS1Z/yP+nxH11vEO0z9bzVTpXNNGQoYLac8r4
VZScLk/FfqU7UNU0m79AqFCHs1i8ZmxFGWnPOook8ItYFntieoIHiY64kQjobe5B7imP/9Pta9kK
Dm7D+8Vr10PgG+u17UXp+ngc4O7Iae4syG4qlYW6Vs3otJQPqF5DSkdeiUuBd7cnoLAz7ADOp0Gh
QgEI3IfLxiHZfPnCUmlTJ++9/cz2ly5XPFXdGdqgKISc4MmspdLicYnpYgfAW3NgpLCGcWgkHqKa
Y29HE8anJnn07aLR/T5n517hlepNsflwsH7kGJfA0Vid+J4DALvixJiRFyMAv6EgP1SiminUuyut
Yxyi6Hy2QVWfYrdoX/gSIZysB6Xg4pqM1+x9AtUmXOqDaiQzFlWJ1IIk7vrEJJJjwRzbKxQBcjUe
6LjGl3IkL8GNnAQ2enpESgPrIb/s7kOIf8dwa7xhqadSvJU3W00Ycd74Z7avzmxpobEPiEuazCHV
OHAIxRhM/lOiMvqy517bDEMFRp5xghlpso+UrouFQeASoBHfJSFBOs4Hh2wCNaTaMcaLmiAG9SDy
Ti0DtxtoH5Re+I33ruKM2vq6S/0EaVAco0dUJ9x4dz/aoS1TsMr+4xO1VWDvPl7g76Zi9c3RUgec
ZWzkcoop59vahQA46mSGylAQGSsIbEY5btk7UDhADbYxoUvjb2ylRIHYAJsVjtOl89rmR5N9H8CN
fxDXQffGMllCbJOe23F7zPeKokEoi5VgeyZv3zpwYIkTulX/9MrX4oRx5bjO+S7H1CMY9T36IOgp
WMCIjS+bfiMIzj4nVnztC2tzQBHezJpt2Z5ifcUuI6vBS4i4kOoTtIem1eZUjIl6K/lD0JGeVLgt
5Jmq16LQjaL/SUuywDqbd3N9gzGhaJdIZyZKnacQscZLr1ouZ0r2JTblRtksznqkwCkUecyn8a0n
/6B/+1OYmohidkqbtvvnvO1FyWUxy2fZx39Va46Bpl6zDC4K6DLO110mZGVhml+AOjFhhYwW6+As
H1kor4/nNmck2rUguwL+oepEZ5MGA+RbhMh5WuEtCxstLP2I5qOxMAEyCYL/DJecSauLiT40abqz
We0/Bw70lm05bxs+0pATLJ9PcDYoXvVmTowRUsM8Ch6vUEniGhUjyD7igrmKF4FOL6WgFiSSjlTv
fX6DzVad9qrDUvMtZPoRD8AoufO/oJQEnWy6MR2cNbibtXSSXb0+hauFX5dURFP64qwC/7UuGM90
f0Q4JyHlwrdDcUF8d19IyFttRY3BG1I3jgNdWyUr2d88hsqwFOEHy5EMx4QEDJDEZwE7GH/rBL4c
3+WfY6Q+31vhg6g7W4HkKWL8qlDEwF/xYTaqTOVZ/Jm3KEIQrVnwmncEZmzBWdTiBvVvJPKuovGY
I5cgQOsb73sGQX1KW2BU6HltkG4DMvuOdztarXtuNKT9D0goHrquATE+QBZPhcnGiQtnnkz+1ule
PgsXW470FMyMkF3PUazEimLkM+15FpHKZa7BjereVFwYzDN2Yr9UvPWr2CCTBhSDuvRa/JqM6IOi
8/9o+7wxR2JOwCbh9n49DRHhNkjJMhbViElJA76oV/1L6kxpwsgJH6hJEmF4huGDGEYREaY/0dTy
3jJlaXaPcDys1YaUt9XzqcXadzt/sdwGJ3NvNWRLjCMRFVqRinK55MCp55jJV57YIZrDS5tCpjrG
1gvpxuvjtmpdodYAi+ys863Y1a6QUe7XeFg/WXzWL6tyxkh8KWzc5uAzWsgdEYd98yG6vjnOYW8I
9mjvNOjhwSVHJpJy/IQYqzB2bDjsh246QmlJ4KcZEw5tIzUg655ag+pHJaWTi8rxcHwxVZuDOD2Y
iDFla55LQxR1q4OBSZUag5CWRVcyB3g6subxS1dB8XAjeME7WfTrBavQTR5YHJV6yvu073uTelKU
nxzpkwfhDSKxwGsaSLxyvSMgkHLa1wBYfhBcNB5uzFi4fkX2R4eTVEYrn7JYfIWSHHLSPYrrJwPq
Bfscq+cwjbLH/jQhDsxdVFehzgSdP09RALs2fktoTV7gZC9bxzzQxhmNzyPcckVoGtYSusHj/cmV
BB6F0KGG6xMgWwbg37vUqwrwNfXKGQgOvsnmx+q7bcLz4DDBMiuLYPn4ay44nYqKhmIqGyFwvj40
h2xP8iweC6wt750951nYHo0jnlSCK0q7TR6a0CWZKXggzYvcNfg/AwJaG+id9+ciiYWKv91eaV70
QOSin0XUa4W/Myh4djdfyqULkplrQmgFViXuaNuUU2Kloih0HqtOEk0e5jobnuuavz+Z1mLpd+IT
fNUI6YUK3vaP5zIdYShlLR097wsStoGH1hAtkxew/VK9RonweeMfupACkeQZXXIx+a4K7tlo1wC2
oXCIaYfoYlfEY+W5wRbgrZDdSDBXwX/Jr2eg4dPh5sQ+C6hlX6VTYYGkqls4z8Y3m0zhINC5qTKh
w6hH60n1QWg+TMQrUYidHACZZzy5fcUbcJRNePekChtzPR+ng9QZ2Yy6LaZ4AgW1sXDrd5cggySX
DzIV2lX6UqcU5GdSxBAoSZ18tL8VnH088pH3d/3BXOR6OjnrXo/teVl/SLGrdCH66nojhb6BwOgg
/a3ccxTdRXmuqmjmP4cvSIZuCEAoqPd+q1ytvxnXVKcPdMSlAbRnIoQsShb2ADRA0Jv4QnkI5rkB
HhBwYjKxDMVmz1VHSc27MgelIvhc1OTniHxCL61ID9kvyUzTJNxL6VLuJa+pjuKD7PLEwIsyM03m
0N/oNQijYzwsHf9P86MX9FaDnZDdScghQg0b+gAHjJ38HLSkkkbPhR5+mBySRbGtBlpnZxkN+NNP
E6po/rgtD1fRNdkgcaRyl1seUwGdAWUq9lc/DxaKnL8IXCX992amD4y1YSloKI/xmDOH482/gMAu
1FrEqiTjskwSAZE1HTTzzBl0C4G1o2rMfDWwhCGi4Fb2Cpul2NGSDoqXtdsOBsZYRqBuZhdEEB41
u59cpBKEDXQiYL+ofxCgX1F43/B++WkVdyZBIgJoaNUTjlg66JAtqyy99y6Ulho3Wka+JrwbHffQ
N/Lx0XdiGuuIA9T7nCBekbf4iPHaef2N3wGxOrDGzdvEtvbrJi5btWUVEKj9F1YEEPiicwRR0qFZ
S6YxTd6PAkNvnBcgkIw5dRuQ5E1nr+MfciW5OnmDJX9oAs496Q5+00ygPyfRsT8jyKkh4v5cX6Vn
D+oLE7Ok3Nc3K+VTAqMLhgYCdBqM1FjXIyT0Yjp0mJCukoQUdLkp5sOsnEs7cSZYEwa6d3V/RIgD
nsiOszht1Z6YnGkLWpp+akUzkm9PWrIOOQF+tbkGlxffUVKgrhz9C3OQeUVYFbjYAdZIIk5GGcwZ
lsmz5zAXxYsMc104HMUlefHl6wMEJH1n68qdw5Ol1ELfndv4gOeSjCOraNcgvQzP+NpF13bhINSc
yRo9kCzYlyCQKatR+oraGfRQci3AZAzYQGv++ytMMWm32RzxjuCQ/2E8EdDQtp66rTZcH0mKYHJM
uWcIXK1YzhNYwUCZZCZWtZHOT6U7H0G2VkDC4NA1hTZuAFh8EnwspZII/Ev1zte8RqZ6rKUXXo5B
gBLh+ihhgST5MHKJ9sD69LKVpt+zGRjwbBe+gDL14wd8vhvBhczzI/8FfuQlmiY30FKmKKdJ+bmN
i0dRRRi3t0C2cyOjLL3ReJ7DOzpoHuvaP/P/HT8yutDEpD7KCmYOu4U1apv8BGIMiBm44/d4cxnI
sakBau+ZsEBrQ7ICjQQtV4yGKAjnXAnCT+Ak56BIQc1urS865V5KVAhXVdUvTkg4NL0mfmHATKab
/SFDeQRvjn749WVTevUfudcP7YVFBlZdC5pbOY2ABMHJAfsTaj59Bl/QJTzDtKBd8rRKCM5Ghb3h
4XAVUMKV9SM7Cv98+YxGWsv0oLBTaTVLFiek2OAyGapuGegYO8+ZPn89xori2xwgcwMmUkWAKHCE
CikCI9XNVRhqiPiJUrZ1DNpKhV/UYRSlpoQPN7aPvK1K93DV5y1faunQCU0l5NiejMrCd9NTYRyl
wTYSB2XBzIvwg2w2aZJmo4N9y31NI0a2P/ZdNiNtVZMkR6bxFeIiy9hhKJHyE6abRFmFtFek3+Vb
NOyjIlTF584pPHX9MhaQsuvuWwZRrNJwsiClfph3V2mOWc+ahCTSfL292m9AXNCKVYiCZHBKva4/
4tYArsHAdn6WM7S80g5nyCRysiYcvhU54O+Me4Jk11MiIvW0yJCJM1TIS9Wb436pm7/HQ48Dm1N5
D+3QoOxmMS1J2wcMZgMBq0uZ53YcpW+AAkSiviwjW/7y+pmvKe2mtlGdIf5yJIMGHEQ69VGGdWcC
onFH5tW0iiwJr1/eeAALmE9IvpPs1rucExgN/s2CQFmQsYy3s2fkLuag3g859zahIfufhzicbpaj
Lx+VFy9JwMZEwK1bgx0P5Mr8+m0aVqaeL17gLWn7ipkPut8RCAcvOMjchv3w3hBA9TgoVB/lbH4k
xPM3S80DamqU0+zwYtt14RaH1h9ofQQo31lXoTElIJ1I64vY8l25QV9kXQek8XkV1QLy9eZrmUht
Pw/AQAWqJ9mdov4tweEF3A623lNg1WwIJDwmKQ/27aaqtB050pQpl3axRESh8lS3R8y9Tb7oUYTR
vSgzKXuClnetpDgBHgtpAnMHHFQLb562FERsKoYMS+9m2MQCFuDH57ps6f4dZB0mLNgHI+GALkXk
OLLut8ckmlmoLJOFZWqeK+DggwfEBrDbsmewpZT126vxyNALl5eukATh316UxBMFTg+emp2mwNom
pA+MxJnP1C9x2F+B9NbfbVuBW66DyUAXXdpuq2IiKbbc2Pk9lpvGE0G1veQCRholuj+5cP3Jh67S
rl9OQLJrpdXbymynGLQ92dfuYbtJ2vUViaU2L7vO3qI6cdw0gWwPL6649u5VaajcvJnS98kPXjOd
WkMvNwJ3KXl3JZuDX4yaIX5hONu5UzCIQa30jgXL/3XujkXBSv/HrvX9KGMsATRlnLzz/sz94IZ7
GSSuKyQWB/fKc24+5pWIJ5zyMmdaaoEzYOoe4DiM56EAnriiTAXxFDvY5T8dkj80+CM/R1OFcRsO
4fXrU35EfoOxO6ahHnLhMLzycDoHhyndIccpcqzkf119ahQEVkVfffZwHPty2YNBP9beEnj0IBYy
ClGrJQwuzfxv+Khn65SofrGbuUlV7gLKh8fzMMKIw+rJMMfpX7hKY/UXf060UYA9hL4HFJiLhfQj
KM9i29+Nh6BuGPy0z6Z4WIfyFE9zhFJJiBYGnSXbTgh9EnZiDUmW5+UW8u4QolEbxHEL7XZo/sxX
PZdu81zQi/br3Vjc9oo1ewJLmK0N4SpqXcWnn2CvcnO4kv7hyWb0f9GM3hZHleKEoXo2V7DIU3VJ
55ZuNGoxSPwMmzr1HYoRvaKkSXIb7O7u5IpngVDj9Hn90zsosi+oN8GD4xB268PBvq+K2bzBAVif
W+PM+hq/N4TWpZhqh9ZaNzkFTdTCr/nCOO2hMvD1sMN0EVXsD464Ex5Zk/KoOe/TD/87vZ6bcMKO
S9txSTH7Ytb7q9bMqg4MMeD/m2mZeraYRxPYSPbDiIN2QIBronHP63RsIIpTQRdr3ZRqpHravudK
5jLCInaGqvUOQtO9rT6VFVdT+B4LmsAs+ieY/WBxTgaFBuD4c2d9wAMCSHFJ4BNreogOE6kXEPa+
tv7715iF+MHvCNzqV68UQDWML3h62udNUFxhqoa2H3welb61BG7I4SUVzuu5ONNhbG1mwHu/WKfm
kngCCTKx34tNNt45dvMCV0J9ebVGJCo+NoF1EVnHrxs83itezdnmI4Q+l5aKA4Mpxp7GTq91zpI1
LEgTsSO5R0xDfJ+sNAyWKawdfVqvnIEFjhrJQyZYZy/c28tZUuJo0DSkBXLvhveEUGJlahZ8NYG4
1x6CuOJu4zvLx9gezTyeayu28wrQFWN+Kae3bljVOauIOZpuxGc4kH3KmDnR48WUvPXW/URBWPpk
ihb7iHFbIx2WV8C+WPHSYhnYymb5CaLXCt/pjO75JO5OSX+1hvWCe6RwbZRYF7yIwO68+9UeDkcE
AiUg7+vwCtsd+xENjTXyllU+DgTAYXuODSPN2pUSnts6/GJmrZ3wbDOk8zB/LU/gcI+7iIG3NrFr
dblzqQS2j1XNnuJwj0QupTpG2zdLKwK3FVpuOeaa/M6NsLvDXIwCxznu1GqIXY65NKpAzWJk6/g4
9S24a3doRpMV1VDecnu0Av5gDmm9/xQnkRZIKv3JDo8oYIR8+MissocJ+4HgyW6RF7XgfWdwDsKO
wCAl/wfIJFZYsvO6BgveJCDq8bpamYvCP0t6DV29YQaIP3lUGMuv/1mCUEEclnx+j9McQGpx8wxZ
+hrcV//CWRFi/Emw4gBqhDhZ/0z890XuwXKUWtrDbv3tXLKgUpfWF381rX6+rBBY2fjFHFfpu6HY
CQ8gjuCmenSFfYEzJoBR4FO04UrpVDzS/9vRKIqQDhKyAj7TQ0SI6NEOREA3tbSEHjWSGQuvorNL
5yTg4wxwtYINNMlQMZlJq7JI/qJbauUR14DKLw9zJxCJtCKPzZoS3DrWL8yIqQY22pCTsrfXnuSs
cJ6+oHrrLsdmCk6I42zhm5MZGlFUkt5vxvKLuc6+azgwXewLzeD7RFBRa/ZIr64ZaneSNxNK0Efs
lr5gLKRSGRzcIbowesR0xaOdbb+VqnYLD0vn71rhj9TUdMhnJA8xWn38p1yXN3JqB7u5ESbyxPN+
x2+djjhI9yZKfT8qcn/ekvcH3ACqeBIP9Kg5+WI6wqVOCKdoC8Llrb8H9PmtoaPLImuPYLIK/Mhs
Vof4N1Gha23sgdCTjsDkM5+6F3UACj6qmge7g2GhuUtvSDt04WFdxTu/7DK5WLOvi0Ruk4rdmbx1
wqbXYB+veeQKxD2gsPokPIk+/NP/DWYcOGsA8EbeadGrpW5kN+GSUof2c+U5pXfF0ofxPy7ObjV9
xIaaoIjeOJrBJBAM66CngXPkL+o86XCb6o65cX1XAt/fTDh+KCZraT+t594RFlGAhkYwIhijntyf
gV3S6Z9a0BGGkEK4oUt1t3FRqkiDs71ehOaTzdH+lrJPPgQQgpFLz3l/Dg30K9ms7z8oTXBuFC6/
18hxfm2cYEJimS+bZil0Beab7jrcyALd7aQxmfV/k4Bt4/cCT3Ge3Ykl48cRIeWsQy+xgmzbUb1S
fuB1YXMG+X6afJk7B7YD29Gw5bzDKLrJyOvjsvCm4Z4jZU/4YibwxVx58lQZT6tCo6qw09wVUs/O
JW5cMHN8X+18mHJQHEPWf+unaqsmAjo1vPE4rwHkvMb+3rOG5KhMqgwuqrwS7WVW0lkBffq9duim
+Ev1kzMRHE2pG7Q7gZEvLJsAZMiTfl3G9FUXpZeWUYCXR831DCyaQkYHJSKeEptyGRdVga/GK1cL
WEIfDp5822DbN3xSbH8ucUOOkesA45hNyDmCPvFxi09GiBBJofCp+pg48tCp4A1pG/ctcw6q+t5S
0BSoyMir8cTHrvxIFDGV2eOfOEpIOhFQo7/upxpwLv51zB40ifrRilaANxsYXJzr85N4NY1CR2ck
BsuiOj2xZnzpV0rWD3B0Nb7h39Wy4LYvirUjxQ56FlMAHlU2hV63+NEDGoHX7pAprterJb+5fyqv
LzMcn12W/d7DV6g/ClXp6p/hg4sHC7fjn+jaKMM7eOFHV5mTzoTCeiKlWKQxHKKQxbO/EFM9xnUr
llFCvM0eBBZjNty9fbsnLFdGPE9GFCAn4vryO/+Rz32//2UVtF+bR0Rr8pZK32/nDh7KKt+Lfniv
5itkNGUvzXoEXJ+Jo9BmvHtTk+Sq8BWD7FflAqQL9LvpdG/wQ9fVHgm3PgohtBG+rvM95obQCsHD
MWYgWmDxloaT66HyR5nmdfOlB3ERo1wdDAWhpvCfadi+XtNDtNEFYtjq8rkRaJNhAQH/JBhUdw9f
aRifMj/jgsc4ig6hLpxAF6B0i3LANUxrf5eAZjQJiE32rQJRrhcaIu2fwQSITYF1yBGsnxW5XjLe
etiCq8XNDqv+Yh5wEVAvQaDoj3Zdvs/FzTS2u4AzFAZorJ8CF5j+qpAQjPKlC1itZiZBUdw+tYdD
SDrfnCLJsbStC1UNxHlqBAPiedoQ8MQz2bDU8FYi/GU36kxqOAvWZTws+DioG2pmUs8dr6jj2JHW
rg8y2/jzIPABQk3bamy4LdtvTgM8kF1JSg/lg9edoUGsIfbhT4VOLJxGrXRVxZ+416upvATJUr7/
eM7mrkTLfYAwbcSnFwbNh3bQBZTWL3ub477huILybtcj6ffN+3zHXY1GQOF5eVzDL+wthxsvCkkg
HDQaW1NGzSn6xBUWoxawHAas5WNhP5sFhOeHL840cBGG9ng0doSfTUf/vLSqRJICOgOYhF2l73OA
an1Sw08PPcd9ALxEovv4+gimcXJzcnA8OH4GdT4o+kma0Td0rXHJ/cP2baJcYtsAcCCoq72wdRT3
RVnQx3qXnLtgN5grn97XdIeokZgCXA5L8yW/VwHH5dHeBito4CwiR9Rq2D1jypuBNXPO1+bLeOFl
WAuT82HjEicoXZwVpqP+j0AShPFPf45Bazs9UlF4UWJTauMstz0E4gciqJkgSLMJuTJ1VQZ9ZxDk
u/LQX7ZfSySKK5q5cxRcE93o32ojZUr7TDlvemdQtFcdrS83P412feNVSeYSC1dy5V2w4i/aEbFf
CR9OVOyTMTxAYacRbDr/9O1zokbFitDCl3HXw6ruLzql8hvyXM/CluCGcVL+FkHJvbwQm2WZ8/Ia
t58sYPDPGeYZVZE1jWWwLMRtFWWOFdziEFkjSx/uGD4SAdLX0Kayg/EQroqyoT7rAEiGK+fxNtoD
wjn3oL6k0UaYJ7QNMVd4Q5ZWgAjlG+gbZwPL9V6MxGcv9vUxKy9XEABcLBwV9nm8prB6yRhsXJT2
wXkZ7yeSIhs+TyYIDj5Vo7jHh32cI9r22O8JuufJJNbKDcgbczLdNL8amymL+UHn7YoijDiMIC61
xuWbudmrRsq4TIU+4nC1Ajs21hplgm1ioWYraFNlhwJPHi4d6GVHOpZB8S9Ve1ghFwSY9BUXh9g4
Futw5uspE08va/Iye+Lht2h7TqPPo2AKNjPS81kbLD+7g2/YLz4OCMEP4TIL4oyOT1LmON7KF4vB
LqOU6p4OaU6hP8XYDCbXNN8LQMwQX2XoeJn6blxNZJdtAO6OdKv38FH2cduWDWFQDJhnKnCrchQf
NB8Sid5Dl+lPwxKDC8AjU75DZm1Ak2nR3dGoHfkcQeS9GzL48k2mGO0n6utlrJdPljyChA7m2Bqv
qu3OPigc+DR5+tSL23hYD42tWVGF7s5hnTok9iFJywwiTTEUYOcB2XeaOzY9kzrrBxcyeyRj1ybn
S1ARDdHoC5IcGAlBV+5xWTg/Q6nnnLgn5O3cQC73L9vzOsEqqWXkPERU8KODX2nrmlYOYmwzqjSl
qAARuW83A+aRNCUqdAiywm5h8yJ9ZuGd7GQWzkFcPGA/eDNPpsZzUzELtFssrXag2a6fx55O3hJ6
GENKO5lPaIc8dGNjM696IvdHMrdWRU/jEUdUdf6GixOa8zO26Rei24RmnNv0V8ogc6EOMsXCOGy/
LXyYPjRjhi6mLxFys58KVmPu7nUa9xxIa7v+OHD7R766OpIhyPUZ4xfY6sG4sNfC4JC4sIQHVOmD
zU/AxFB/FOdzEm+NTkn+QTzdtsl26XUUhwKKsyykjV+ToCiH/SvOstRnuQ+ilInzfwMdTGtY/VCR
iz5ZSSdRNV3jvNdw72I4xPYQzTX8QtfQbua3hlYur0r89lZ7P4H1fkfN/Y66M+qYCS8lf9nhuJQu
hhFRp9zbhX7iGgYOL5CHcYZZrsAvySozjV+L3Edn6b8Xv/VznQrC/UBhbZLgISE7qIH0pR5pAS/X
RounKhKshruln6VuJPP9AjkF3/2dzZFtxYUnqbWrwgivG00kM76rW9BKSpebN/rEHalYwOtX42UQ
SvAoMnQx3RrcNQzgLIsvEDGyUHgDqpLrLCYmjf14EEarCyhD2nBAFrX3Mmx2T2GWOvGwa+/3pgSW
Yn+1ExaMOk+HLn6rLVZsRZucC6ITlTdP6ZIrLd3MmAaECpKwEvXrrhaiUxdUi8qn+4ff1mWoofip
i87yOe/YrqJ+CJX2iYXsj4otDKFqfa+8kenlwHioNS8enC62YcxtEPe6Yxfk2GM44AglopW9vaZE
O2yjUPTBsuXBauiTYkwkDoSUNujZ98QQsrewIuNTtJc2AVrx/rdA9B0kmhhDxB1KpBkK6IU5Bogn
Djid69zPMwlUllYJ78B1tMmr2R6JkfRu1X+v5nbL+r0CRy9lTv17CLECCDAJIyGIt/8e4gIhyX+e
H+dFHX0431+hMvC/QvUj5ly4BvgN/sglk0Iog0XwTGqvBK3BrYKTZCnpmwbW/rgZvqWWAoGWoyVs
Pd3Tj2zDnO0r7idaY6QPiUa9N4q+1Vpz7/9MeyV+xTXNQOVL69y0pxZheij+uh8unTmBzfgJFe5M
wmyW003sbVSLP0K9zTmdF3fi0y1H6dqbnJ4bMFlu3ITzNsZ/I7XSVHhQu67KqB++xU4tjPd9jWwn
zHhUQbMB5GonHo8bJvD8ftUdg/QxjTity2gslOkCZc2bELlZ+AejJtdVjQRWmvFcOaUm+LgiaCRL
tO5o7+ngrKURZ3M7kTlWP561YRcTYwFtzYvi92Gq4EnHhf43fcR8kEg7g4Yphk8CLZmQYjDqcUfH
SjMJZwsFZGJFABd4hScjmfWEq8AcXFaBYupCb1nU3rWYIVvNd7FpCT0jYOKfrYEjt4MbYZiN9lBE
jcHLbNnZndk0r5NuTKnf7NngAPzxGLwax7f1dHRbraOrEFMLM8P6NlCYw3wKMV3ksQpMEgnX+sHl
R4iLF9pusS2+r6OV6zQAewrm6r/BiAPDBAAo6f7rUsWaQrXCPL2CArqiXRtwiRcO1zFiABmV3gcR
rljWprnLphJHCOs3XraCbdJvLqJ/yJ4UdXHpo3dwO/MFy/PUpE5tKorf05qpZqCBc5OGk2pPZRHk
ELsqiuHuvOka9kKfDGwXpIN+NF800BXR11BBRzLCcRb0o74SQKmsG/v4HVkWlPV383pznlzMP8vQ
Ksn1t3NT/3RSOMrm5T20T14ke3j+sqhC11f5Tzik/PEx4fFA613C0GQXGj7P3UyFJP4feHkWUpS9
IjKeC0HbMqnzKmfzb3myyN8SzkRVHHSwOlS3n30qw12exAeFCmw0V2OWmu+ppzLrG4fN2trq/fwg
ZEwSxrSv0SAQGqpxefzqPVjqogK9Al2YzrpUq9MqRxFJ8xyOS/1JqzJ+Fr10Mqhov0AJlSGAl69l
rBN929Gx32IrdEG5pxGgMQZiFAKYcb7dsuw89EAswr0PIyUH/cyBY7q7i4bP/TsyYUl/eSjPKSpG
K1OYHM3/E5It7H9VDExGAEC47cVqq77MPR4ORm+r5mei6rd76OZ6cbq7m+n7p/6QAtMqFfcoklLZ
oPevTIkFDbcR0luXnW6v2l7atyRg8h6KEKBx3ZCG9wbVE0Sri/eKHgd74JCAzv+xouGxjzunaH1p
3TjHlczOeQ8I62sJf0F+IWVZvVM2Y/iBZAPd5SznqbhuQGeaw3tc6W8rOeOtgDTsjjh5X8gg4UMu
19o7J7nRCY/nmgeR55FjS2KJpnoJa9bbtOnFi1LtddLkST0/G1ocia/TkD1DG3UN86loAzKS6G5b
zWO1Db2RyqRKBiv+u8Qcv2PzD9IQ7737uxi68iVy7Yu6xXU0CMISZYmzTSTOl/usg1Jarz+aMlY6
gkrKH6wtO1tnbp7jrnuBvdP3H4vSn+Ki3Qp/N52pcJauHf15Tw9b8P0T91emqaV2Oh2oYfGMykey
gqRPmxpCkYctvEjcsD3AUdwdGVA/8u9keht5/LuWonMgl0xD3AuUaL0lseEg/OdPa8FjSxiiJgm4
eiBTEonVR5W7a1/bE4lZigmQ5nRWAY+1MGGvfLw4aP4d01P9jBYJ5ZXDZ7xV819pzqCu65g1c0K0
fVv05CY/fvVe/wsuixCzBnw5f6VBvb1E0ioW0N4piDYvf2Bb3PZ+wE0p4u29mHQVoaBQzh9Hiomh
Qyq38CJUV5/00wn7EH3fsIOeFJmqEdoYlENDINW4YhXa5V+aEcSOz9iU+4Vcyr9fxuGuXhTQmWuM
IEHswOcxjZ25H76WfrSCBaqt5K15ZkUUGZXJYpV/TfYbTKm8Lagz8lu4Kakt1gAGpk31h2V40Iz0
QzMmPKYi+pCwLRYKNl0eG09CeuJzcbzf1XCkg83vLPTlSiFDDib50WZ94ugkRsz6Qd1GbrHUMXVr
hyY350Jb1j17x4JlWdLZeBqvKF4SUPkONotXU4vAeI9a+D6prFf7FoskHEt+8tCDpyyEJ5FMhMu9
fI44I4DFO99hfwSr9NDfZhYm62dg0jHQAeTr1DLmPLVotlfexs59I4CPWSr5BYQRGZN83jcm2PvO
jev/KuZez7w5GVOkk2JTtWl/ungpje+s2iD2zKWxA3w2cSwWwFRhv+fwmrAw3VGiKC5x4+ULt0Zn
V1omu3UjQ3bqfq2xlnouNoogHKX2qsmk+OgA1PZLlcJ5EtmorWT0xhQNCxgF6pMc2y4BRK1J8aWf
RInQBoX6z7qUY5ib5ktl0/lL8YifTfgVB+9IKaYCMWAugSmjbvfLbgx8wrlW/Mf9obKjf/cGVevU
2qDCeAQ/pA94AoH8oKc0bNydZvpvb91IAq9hzbhklP930XIbaFMFdVTy61NmYYPS0bsm98N2qGko
I9wpHNW5sc3Jmq7anlJ8e+DmF4lFVoXN9dOuN2XFhBT1XnPYhySrly925pC0pWl7XeamKhtV7wWk
9ogTP58XY6kp5B8548NK5RNn4UUJc5ZSGVHgcakElchvf0tO4Wi182n/Kra1dYqg0lzUBa5R2G1u
c4os++w9c42nIXuu1tkKgF0oV4RyDnkulrdzmrOVQPu5jyJGweK+JODQd2x+RKuzm0RA7mQX5Jmx
CFWXoJHocPJoFcbl4AF7rFfC8tJVQcn39tzeI764Q1B7PvucEK81k1q3V3M+SYj7aaBlm+UsjOay
3XV9z7yHKssVzqTTcS9mzJHQ/webotInlBNN8hSPLV0UQdMSBR7y4VjOmIoznTZFN5XKyeWHX+xg
u/IMC93Yj6Au9zkhppprqp0KBgC9SVctua+Qmw70Lj/ZnxBomyNcu6O2aKESb2YUOyObwUOXDVcY
d+HXJ0C7ynS7GRCagPTSmatBOiH93pfDdruxo+TEnKXjqr0M2qdt4YvsRbTOhOCRqNMXhDxq6Kcw
fda7gfTySkUchbtSr4tUdbqCU8gFj+TjPepX4V32/jolsCHJGHDc2xr9dEX4KLP6QRO0dWweKcsS
rlUfWESMuhiGVoGJ1nM8Rfk1lrFfc8vy6GVswMN7TZnXx5ReZ+eRA+Lj/02rDL25ASdrlXv9vrzB
WG94+rCZgkaINEVAqORD+qETni3QC8UO5DguYAJDrJUDabahE24MV/Ty0pBHRGfJMISyIgSbV4ks
rBmuFEVkPOm1E35w/uEbzqIScwKRWw2S0L9xRCorfvJ7lNBUqDjYfJ8IRPJ/qYROH6Zbu+ESRrSO
hqQx2XUqxMJTOtV1wGlKZ79ruzjmWTvX5quzrds7lC43zsBccXPGUrL7IMio/B70A9Ju32WRRtz1
qWZKt35aBnsvASdzDYXjor0BIlW0uqxLOrdXa3TgYVJYkG3UOjP2rzNsL6naRM8viT+tvPuaB8XL
iUboSEZYbO4AySJy+OLufHlrDZG1LH9Fx9yuFYm/4H1cSlW2bYXQcKzzxl6ATdnfoMU09jwdBNPe
cmJBVpRKqL0+cn2DH9qq6WMGI8WldOWmezbL9I0gzW/GrHmwo8+twFUvZdIL2VJi0WEXEyho1Xj0
gUv+26WFybmiIOqElLkKG1LAntDJpA/YFpNZCRXRpL6B6c9f/L/jJYDGP8bN9FlQv9cF0q/BiGkv
gm6RQiGyW5W75XmqnzAZo4q+UrAMPlN/WXmBUwiDgt43+RV4aBpBSM4+/Gqs8+8UYFG+ua9vm75t
XJwi9OAE0ACUJodI8m6o61dTVsNrXCCARGuo5Vgx63SdGzAC5Ogmz9/7ejLnE34pyJlAcBlku7SO
nIQRL/7f5gna4BdSEM7qntlTSzLTf/tvvwYF/j9h7YSrVngk8KfjYk/XJu0QWWyqA+mjdeusFAu6
NldDGH6J6Hcm8VSe77Pvp37fa4HibAM+USY5qMFRTb2IbjUt+73stSm1yVPfMvJ5NWK9uwibz4Xv
bMZUtnFCk5T05U49cpwfDOr2Vw8d48nrqgDkQe966ZqsnMX00mMX5wFFJVC5D9oD4nnuzeFrI74K
F2yP2s2DwQMimHPNJm3g7Qy2D0rFsdb6wKAUxVd36dXIPttjRrfFbnm+XRgCBGY9Y7aUPWg03tNk
e7ulQKxv2WDxbZGy3IjcK2fJC9kzAdNHB16sNFEkLiBknC1yDO5uZG3hGtf+gSgv6IZ/GYYRILe+
XaijHZ0PyorxGVca7Qu2W40j4cn8xCIaT47PTDh7MKrye2ROr2r7/dsFaBxQ9yjR811oZ7dtAlwM
HaXS2wSqWFr1L5Tj4xcflCeCFLsC+bBhn5/deaiLxqiK7488yjDAxhIJMuV3bP/7F18BhFp8i30q
xRvSKhaO24AIdH7kpUMGE6KA+q4g8REWA81ZA8yzHdej6xVGgXGIrLNogA/WMHmpE0P3/ihsjGqK
A3Tmwbjn8QnhHCOu4YEy0AVs+hLsWhCA4THF3eXFs49xVLyDufMd5RlRHoUGi6t1XYyochPYpAla
47uIpUu3l+Gj5W1AESOQ0xUw1MICk2yXzWjD29bqdNdmCO1Uyl2OFe2uORR8h3As74drtBj4TdqE
WR36sYQyhjfs1V4CuWeXbai5ktfUzvG+BN3cRQFsGrQVX/teMBStJ9nhoOz1cvPIzHtrjH7Wrj5b
S5tcREgZX1z1UTsNrfHHB09OxvZhdhmbtahKHhuRjXv6hQkYr87TuDB6xp+5GT2Zb0VwA50HJ0GX
1uYzfzvGkA9VmLm7WpdmvE/AYhmVyfmzjvkTVIHLLxmtEhLLGiKmOCRYeayo1Dk7yoJaW9erlxVH
FX+GVPbsXvldfc4yW5x2Juj8fWnTb1jJ5ta+/V50VtGaFMt3YQ2qAjbygzL2Rc4t8LLEEIk5Hv1l
rPoLejF0GmCs0fAKgDI+865h8HoNFMf1FqLw7IGYbc/aQahBR3RjJ7mOl2qJpnscT8DjHUAaGCPh
ZL3qM37K8xBfKNAMaxr+SbbvlPsZ6OKSvOgDSxyR3rih1+F///EjrCiEI08iWXHnWnInb2oSS09Y
DX/INRYDJDLqG4l3y4kl1z+wUqAp5D0607cC/i2kzS0okMWbG2tj4zXT7MS4DS5rYHCRN7qpsGpv
4n+we2xSI21O8Ln51frbxN0m8rMQ5I1LNt93h4PfQtiZs5Y7Oge0dFeOV48jEaJfgHLD7dUXZjVs
SjgzyXhfW2tYrYPbDJ3yD8qg3W+9kmBJNZFnpqIWc4MGnXFtmjphYH+X723lvF2mIGuiWQBMJ4g8
5W7H222L52JyvHhn2tz9QC/aeCY1eob5U9fdZkgGHal4F323WqE5Ocdb6BE0s5ysBkCu9jjusEPc
cCWXIARzAoH/WohUn1OlM25ht4vKWzDeZk0FQfhJ9aIo1NbQHkM02QO0hurIghn5WxgC+NblIhhN
RgEU3z0zjlXSkPHeibBdDHYfM11xpraIGkCrDC4o2BhdE+Dzeb0uVMYhmjoaeiV0Q1onW/DF4m1P
77P9jKx8YfrzHKxgIupYUQXAhnldBVWUd79DSMFnCTvRokWkBFVYNOJjuMPZUmBDMWPG0yIOgCY1
7Gt5vwzT93YLcxQ5qN7Ab0n7YPtirROa3b7Rw6scgtW+ULU9AH/Ujre9EHcCTP74dqswGLYP0ALH
bNB6c7R+HN7r/RM+Sqebbs0YAylXS92Pmibcj6HuL6SO65e/+/Vg/ypB/vYDO+eG4pAWDX8QZAch
13W+IIjKkqrRZl5bPnAncLyz9MpDHyL4xwCgeNhw/WkmKxR63Z0hQC7WYfTzqf5Q60x8DFV+Sy27
9DOrgPs7p7lALvRl6HiLl8BQiYfqlqfoC88H+1VwsItLrKGzCXhHZ51fPzC/RKirHTqiiG2sau16
eYvH/Yvpz7/b0xGR3/DNNLuewuyCzAhSuZ8l+EHHi2tJ0XMWyvH0/thG7Fsrom/iHGD4RBR/Ux0F
67HalVnOdi8N+LYmPUwWJFwukvP5axz5LiZBPGDG1HxzEDG3iwtpk6kqw8XAwFE/vxALiffWpeIm
OJfDbpcZ/31ByD0lg4PRGtKsI+DspYV864H/gJ6w+XKb3/yaHd0R7Kwn1UYMFGjAhAWmlQjndfv3
uPPGolez1znYMvcSQHuJyU3boQtFLN9ip7rcD1L5CZKs83yF1Gvt4BJETAkpbkJhAqxYnNsfh+te
Z9S16aKBNQxnDmOEFUOSFMzwS0Ewr6THdqbEtU5mSWTKAHgHX077OQehsH493Ob9mW6eJ3W5iGqn
+8eI1lXT0CJnGcfr7voZe6kpFHxRD1OR/B9of9CG3wDTrcK3r13ohWUdXcAsIImMz94a1NWzwL5Q
x7ull6MYEpgw5eLmkY2kpGG4lTIJikXN6B9M1nTxqubiHzW7BaEHoSFOwxOWS8fKEFOPu91dXgyE
ufnUNsUZddM4lGK0tXHWlNLPqMVw6ESA2h2QX+H1BEJRNKTQHgk7QXD9HS5HhGb4AUzgyccOwH1D
WydSZIeeZ+ykkOwSoT/NoNzJ2R632e5r9xk+8gptUcbtwust6wFkOQeg7Q4S6fLhqtMWQXzaMug0
tdjofrvGaKw23hzEKFg8mBX5PmD2e6yeHCy+Ng1oFveN96DbHLkpVa4YPyA+mDL+4tgo5lxIGDxe
2jx3ef9KGhP3D9eyM0TahCh7a9coJpxFx1CFZshRxlM9Kou9XD2GRyMB5tjAOxThl9V/xtyeJOTU
jDLWENHkH5Madzz9tVfHAkQE7UaiNE3f4sr67Fjb2Iapp7bkl02EURyZikziQBUWHH/o59l3iqmy
QXiwBcJYCqvN0+56yRTlyjZVeP02BvTpdolcJCwOSsiMRUEI/Y2N0AdouW0wgj83SVbOOVJQ/xM4
x44AhMxzzQciSJx23VT9ffmz6SDP4TXcbXzCzrBPzAPg7hTtOZCG5K97UoOHFJcLv3MqbM6eJnsP
xDBGNPyBqkGg3yYTaUVy/swi+kV4wFwEkFXVhvFDoVOlIseglQQnx2J0neFZbDk6x0SNFwV1lJkB
b4lgcCE0nNJXvKnGiah4OBHrZQah7mpM5oFieDERmI7MRyT3hyeLq8VClf+Gd+JqAWVsqgy/XWSN
LXzC3hHzmUUP5uMLcVuIHL21RhcTw/jRNRxWMI5po4zkqJE+dra7ywymAgabrcPQaoR1pQ9XFzGT
GpB5hgOxAtlFoLZVsSWxi7dGIwiXlYDMvO4utYZuFY1EjrgVgroc25F3nS3kXxAe19lJFn5n4uvt
DUbP7yJ3tqBU+QKoSXtVafzSWqxEM5JCD/5IbScbeTdWtB3y244zDRsxUyrQLNq1oqa6EpAnhIQR
ocZUpWZYaBnlDRU1uUMRHix8IfT882OUEN4q5+e8PwU8jxVo4cncyfZXwBKL2z3B3VEk3R6IebBs
oMd4A07X5WNoKULH/fyZyHT0OenUe/6+kvatgzuay0PYt+vAkhd1LD5OY2+lpTasgz2LkVGrknC3
daL8GfrjDyydstlr2HSe8r/stM2xDbDCK6KIn5IYqu3N4suCoKVcJlL8lcgfycW8sLh05ps0JQ4I
MSc85qX8+gbZy4QLm6alVUuC+EBcFv/EeU21NyGbY1F1cLQblopWd+re7h292Empi9/mVDvlN2ji
5iLfOKJbG2Kq6IRDulgbGkhLFRlMd0hvh8AKzdYc2U66FtZmp+kjIlxTGbfUAyU7gWzSowqnnDYj
kxFcXeN1admZ7NlsaGIXoJ5OMUS5Tm2MPpprS0p46ipF8/GoZe+5hn3ZwjwRG0W2gvQE5biFJJA0
BmeY6OiNbPKPiOc2RX2Y0aACkK1fqAbvl7MdGYxpzAkLfYyiAAvHORanZeyGEbaZmnbldnpvAN56
c8fn7xTeYFm/b1vtSjasEeNGqEiavE0QKCyPoidLN7+QybYbDUP43HbpJswahdjXqTjvS65AmyUo
8I5wi37kCaZJCCKpR1mSJs3dMidEq3foIzTGcLERE8m4Mpob/0vcxrBta3SQ94lTsaCYZiUKrYlX
WUkeFHjMoKOqY52TCop7afIO+cFffONxN/LOpU6A9pyNpwL7ILogVi2k60IKQPnyoLRjmR+0qKNL
XyrvxxSd3fRRdXjvsO/2hCPB9Pwwx/UVc/Sh2xJxH5is97YxQbNC0o0O/AbAM8oo4x8ioTNPqwbs
hh8LcFFes9kxLyuRgCWGpHNcCzZMsjLhQt72k7WZ6j3LP1ra4zyDZ1eHLs1CQpKP6kTPL9Zkq2/h
SKfnTUhblSRzy07SQAoI2LYdPEdk4p/bNI2ijPWkljsnQ3/KJh7AdDkQ/9Ux+NclfLpJyyt7aFPe
Dtar6xkLsLuKlFB563f4jOzDVB4OwyeX8iLQFspm6QUzgUpADHohfR3c7pMtaXJeGNFfRlI2qvkT
64ransVT1sIdUvNKNbDYlPCfVV7vTTGu8+cqK0YYRii4JRFs7oeL2W5hPJtAliFvjZjCy9SJE3Rp
d9Nw3B/0LJ9F7y/njhOrvImbJTORC+C38WDgaSxFnOcB5D+tCSh0g3GxePZjt/4HzSg+KTRXXoFD
eYm4oAPQxfOTqHScRhnyt1ja0+U2VnfyOjXGpANa/v4ilSAk+oyD2HUdaEJYo2udIlxlVGh14ibt
inYUG45f7pjPgzC5Qp2vdmnqwdiIXTGMcHEOXG8kCXJpQuYzJEqdWfRinxRqIeQYfqf1nX1LYpQ4
0S6AOAMiwnm/5O0TIVliYtK9eMKLPiHDdRZcueVIbFhxjMesajzFSqSFe/rR1qd5LxZD1gHEhyFD
xn8x2VSlLPZGccD0fA7ltAuViLWgY4WiWCopS1QUvx3fWCIjkHnsYG0XzKbTnxAtpggz0g2eQwDQ
w8/24Q4WoesJWMFDn5PX11hXHS+S4UnHGqpWpJMEs7KZ0NPIAVP4aca2Z3IjoLVPCYz6d2x/Lc3K
CceF56uqwJln6gqr3Ftw1yjiX+h3TstOqx8UneyqUXfUPARp+f90vwE0iaQjGuybYNWgM5krLD+N
KlwCjNmJRdlP/tNd3121ZjSNCQokV4OcG401+1MrA81OtTy1EO6umr0Ttj5uFWe2wdAgoJwl2aC0
TtSZWimqJ4hFWg363B7jooH6rKxtW7WppSg6ebRm7qKof50O5bOKRnLW2ed0OS106yTCPoOv8LW1
iQioo5Pj2D/AZzAD+/m+T+W5afHUgtVeW5cibuj3iLXhXAl1pnRmi1WTL7Ei6tI7v6OWQ6ugY4G6
8eNfktx5kXl2D+jAu0XtXaSorM5Zd6Ji2QVUOdij5DKKp+ULXb9S+v8DltSMYNwvhkQmDOh8m+74
JWSk2uYuQDzHaVC5TYFTKAR1HRbyMxYxDaw3OOSAuQyhGSQZ26TJ4weiQ8d6ts8sec61IUBLmhdH
094cpU8b+5bTcqsdipOPWVzFV/dcv6Mv3E6wsj/BMWA2B4HpFsdUG1uLypyWZB2lU1DB0KW60UQD
pssNClXgrP9SGEO3ZJiSDeNPeqH/s/stKI4WoJGEZV3IR2tm54oivsxt8luFdDSMV1Cs65pBhIJO
SEjic2j+Z6SnwHfXBe4Ilr+DuXgMfta+fdkjdlFox5p8ME6PoRXNaTSUf/7ncESYXJca23s5UjAf
fdwQMDyZ+MNTj4k5ucnzQRWR7ZVtY8bcvvl6OEosljPMTSvLlo820Lvctn7gDpTnLbLQTU65vKhB
wBXJdWCUicSxBPyUx0ByPKFeVy8mD6uR1X6NBltaLKHdt/aL41bp3kQPN2/CiCZ/Z8IPC3A1HvmJ
oA4QzbIJlqXqiBirKnVR0EzSCCjXSiXaKGIx6zJiwPp1A0maXAmMWid/hrBYVEjCYun89DEEWYEo
bfOkNx1kpKe1IqZuvXOE64o94lPYmqLqu/V/Tgkbegb3//uvMqBo7MqdMZ786tH+X/j+34v8msZp
fZnOeR238rznyheXqCXq95pUzZuBPdpawYj2nRzyJYP+p4uhcl0V3c35+EVb+NKP3y9UsErugZ83
EucvR3qyPSs0YYpcGxB8Y5LHcSa2xGd3B2yotBSLiMpaZlXrjvcd+Lrl3GiKuxpkzy9Ohxw+frJy
5MdGZnODLBdEoGomoDllp7aUmWuDtRMnQ9UaIzni05kLNh1scf0Z4idwu6tHneuAWZKammzA1vMU
qiQK1MzPCe0bbTKX3wgdkXWx78YjVJ0P+i+pBzRp1pUB+bgVcSGZxWwp/qRywrjwleDc2kZ/cJHR
tT6YkuHlmOjX997YLVvE3FMZqyYpaGPpT0yJfitJq2hTsDy8XgfNkIAfIb3VQA6l0gw/40x2u0AZ
Sd/cha3e1+/OS7Ew9Cjr/U+22KewS/dytk9W81fvK9kn9UkrGNu/HjMgpeFVYh46B1z5MMckpkrp
BOZQGytbVaZht/Cd/mfjT+zyZGOonGgG8r4m+4hjA4Aj+gA5YynPUgo4yVA/zvadBLLLvceN74Yg
VaS5ZBmBRgDsTSi/uU+ZjGXCYEXj35dLij/fLqSaRJSpZFQHNcLhQzuz5FHv52Q/Wc0rXYboiynD
cHzU36RQcENYPKLX8PteqglL5tkRmjSUcm90z4uo05/8bZQRZybbDd5NJmGhH7Z2ajxY293Tpdx/
X3PchnR7QqLCI7BU/UJSrE5cRMcF7ZWCrtRs0ZEU3BP26Mjauh/Zkr3jK9+LBT9LO824T26FOx1b
ijZ9qOme4n2mPjFYrZJzf3Gu9vwIwAnHB2b6sK2SxIXxLQ+ENh5g0NHjYJV7Rco0ffZqYzbUxKRX
TfCdt64HzaGbycX1Hzrp5O41XJSVGFijwbpKR7HAcqJCeSEWfQDYB1uY08kzwww+BwG+HaD0UCoT
kzg7EQhAc5ZaTeDZBKA7CDLcOfP8Ifxi6MT+Oe5KJUWrZGzNsUKV2yUG9/HF9nwrS8XpTgl4gezn
eXKJdoMM25WKoe6n7ODkJaVJKo0KfG5NXGBIT1grEW4c2T1lv/f37FOtPLKYE6GWDDmx7PEDRFpV
a0mG+EXiQ1ktPkLiws4//y6BSVQkaZc99FpsO1BucC3ebQu8Xhnyy8A2bl3GGwpaYqMgTFM29P+8
3qLnbBJ7rmivVXxecaxY0ilSUD9OW4+qN++0/7ux/nm0Qjg7FpmPe9nTrPEe8ySfq7W0QHw31NSf
aCSXanfRSq9UMO+Sou1KuozjmS/nm7R6WoX2pIiV8YWfFUJXu3odZWBE/qaLxsYGnw5527+EUycp
+a/OOOS5+g7CW5yBUhNctrz4Nq75sV/U+PFi0s2szcG7J7VfT/drmTQ41dbeK0SwJT8LkwtEnPtD
KKCtpOEQrtvnW5IOeJVpSaF3EqPTxRUbfAGXxNE0E5nL+hIR4AE4k3oLmwBSJPnbiXePsEv9qHHK
G9MKhQOW+pfWTSUDFidntFd4S4a4+5RRtR2oyv081y9qplRuym9HEGtkSQXqXVxs0dAs5i8WS4by
K4mo0XfeidC4cfMBI0rfvJF3LKaCEoAaYzt7k1U+n85xCK4bBxgiRv+jaLYmdhx2HdxlimkSe99T
NJpeiG/P9M2P068MVPcKGebwHyBKhgZoyVK0ML9EpPfmkLVLoZEwNFtejpMRPszc68wp6u0M8XMN
rWL7QpSFv1ed7m8w1Hn/J8yyCQ+JlSwO7birgfEeEGrOSZwDQRjxF3jNYlWlTsE7rgU3wUXD0S3k
hxKgXIUGbnXEMC9Ry30a6CZQH26ac+SNMTJ6q5lwGs7+idQhXBp8oYbBEzgdZAy4fCB85boh0yDe
kPVwUAqtC7m84s6Qfh4cKdAssg2m4QtwrcQi6r+3j+ES0cYDZ4Dm7XmSa5w37/ALFmG8vwj/E4/1
k8spfmNKMmPoZDJyVI+0ZfyjLzJ6i8dCooW7blr9Wn0UYWRbtMRwEl1V9gVmi51unEkTw/S78w2j
6ciYATIiMP5VN66sFn8ooLlKVgKi7tL0d4VEZ/88qyjS9nJB3LzE4h2qGnNy9tol0FI0lsUlfeFZ
uRS6wgLTBBsbQxzEW9piEzstQNoNEOqukbo6c2n651J4Gds2FAJI/qb6JKGpr5MTuSAa5NjI0R9t
zBhpJPoBnXkCS34iXxtkhe0DwQGRR40SxnCJ/CQd3pW9/GfDc8EL5A/CKk1lMs1mPm8PoR6WwlXw
uImqyJYDJ6fiiCw5x+XFyXjFNC+4qKkQ+nLmn4N6R33/eyHha4H2KTkfWPpbkZwJbV7bvY+vCNs8
AZqrTSwGfty4kJRox/svC1a1YEUMundXaoYk/ZdsDP2gIucQuSnbvTBRYtHAT9u+/aPRdcQ/ai0i
R/keDGvIcm2uwXmH+lNZBa3V4Q1hMIJ+E3Z2jhixTVeCTJ3B01fmjWEVgmSz3yXbpkYD+g3d+tde
ZdexVJTI/axsaAut2FdUUcsuY4OX/mVf3Jk++w0id1d0ujjl9i51zwGBYRuY1wpIUoB4OEyugp0V
EyXc1/pKb2Pz2lZT1ewDWwByaerAuFFeCdVpLvkbj2SHLV9iWhrYdQ9c1EsfFrk9BsyMP2XFPkxj
E2cPF+ptSMzPUabYWVUE5kb9vsSOg0JlG8b37hGdMmc/ulPjXQzQUaT9kwchMI902RK8Kti7U0nj
uV4L91I3Voz+IKV4mxH9zWMZM77I3J+YO19Qvbete08WeQMbHaH0TntUVvI3Ph2aILzqVggq9bfZ
2TuSJb2NXppjIzfN0eQ5l5hqb5jHb5JoEtOjmHZEdnp0dKtwS3HwiCBR0VIwgUrYxprtmAK2UX0N
mf5DMT0VRnagcvZU5QqE6jwKLTXF5kKwRCJDs61B/xtcKHNPvZ3MBUkgy2vh+hKQMJnpu9bYa+o5
qFJxAu3Uva1Sj8zBooL+u5fJ9dJhoZN90oJiSoSPUzPy7qkYSbqZHeGvTHDHXWG3W1NlwjooWbWb
6iCTlroqv4iBUHdyqvdUUv8yPzc6EYxdSYsDnmyuZf677qOfO43P73/mkHZI8p0HnGUKdO8cX3Qz
t60zRgYht/12MHZfmKpXSQoqhfemVRBEDC0eWhAVIphI/lL43KD5OIv5UjIE8CaskQy0cjjcLkns
j9FOku6sAbzb54/3hYd9GmE5nBM+uLpzkGzIXMOLWsY9HavV+nP1xq7PGR495F1Z8uHU95JPEKXA
YJVxXT2zGHS7FyvK5bngOcT/wIE5P8HIk57UEd3qqjANCVSktD0Yd8enMo+fa6+2+BigGBulrfbA
fZcNMRDr3tkvalIoBhuv6qodszfwNi8BylR/B749irYSYgwZFuinClTbwKjTbuQ4eQO7X4BrOY7+
qzs0Uumr7peG79mBmSqqymT8ZxYML2i59aHKGzZwteNSJfBxQ+LXfrvULS8rIYzdFnpPSz+R68ub
cnyD4zeAOdc1g13+NAkfqKo55w4S08O7GYOT6B/WVC0eylnI3j+j56zGO3v3AWz4jrWPN/eKI20/
Txlg06U1hWZUu0vlWMAPQ5Wj0DHOYmkKwS9phRU0aXDbW3iQQDUz+LJ1VytM9Brl+IMzHT3RVqKG
1yvqVCohAOLsGz3y0Ey9tWPXVwFbrfpPjadRIHinwOly8lVhFy2CqM0AI3XRuBZzz0XCRdnnhaA0
6paz2DGrE1maCKkO1cm/0GAepKj5rWMTHmNjc/ySq/ArTd9kOU4+nwZx35G6oZ6LhDMop7qI+paE
x4o+W+hZL3pUZ4Xqh9uOhwGe9CacPeVBJ38Tw3QMG/jdaBTThXxFK810/ynlrEYmNGTyrUIwKC9c
bh5lgxXFvzlpwqCJDsa7Y3mQhjLwG6h4/fNgIHZy61zDz9B5f+RUHiSTobBIRlF2Kz0ytKhdrlrB
JLpQ7amayH0G0x6jzyQU5IPT1hWXOmyaohV3ZIX2waumakhHU/XWammvWuoOsTT5ExycrVhSJxlj
rkFsXsoEO7PBNihNEwwPWpTv8zohVbVAwCD9zonKZfg4EemgbEPkyhT0MZmYjTz32bGj/PzIP6z4
OuNqhm6xr4OnCKAQFvrAHuERAohiZQgrL0LXMM9kSuD+ijqe2+Jw2fEtVI/hgKXch7b6Bb0mhXE/
4N7IBUjyxJC+j56FaOTELWlZrUlnpjPtyjHnTNHPW0/jVtfW0Ztoss1HcCCbTQzvdB3d0HalkMgb
7bWRTfY2X8QZ1rjWFAfEOOO/4PBy2B+rncr1sQXg3vBrXwK8IpIYNbiwlFfHzBhtyKMpXUlCHd4D
CXQyt06/Cq6gtV8y+BmgTVqVT96JbC4+G2FomHWmOQytFYkn9mwJP5id+aaiGmeWydyNkQH7LKZo
iQl6uAFD0A8cfMC4KdVGVpE6t2U4ZtKWuo0suGC5C6671332zFqK6K/JjFpCABgGObSj8E83fcUE
Pw7Z4U4CXixTfSn34U5YPIRbkC1aE8kTBsSCKtfq8QAc0s/VOxG7wgCcSmTfetShd+NnphUrtZeN
F0NEkyvBU2OHU/lBSi43wKdv4h4ITjY+bQuCjJNgtxjRDnm0biib/+Owilx/wKLcGC0g6EPSXQRQ
JWU/EdUfPdFP3k3yOiYO12qG9UpH5aUH1l3wTPKNlKQoh1EVJJAGBjyJ3ZK/xl4Vh+IqN9flRcUh
LAERPy7TnSbJDrg7WAFXyrEbBFoJKVdjRxJHYhOlJEf+eDi+0QikpwYgpMELPc0POyxweofPGzxn
DZGSR7aZJf+ZoOz8oH++19oL8GfffXAgIX+/8oyLsl+4g2w+Jj17I7jci0JJA57sVNXJ/k2Kc3vx
K6y2FurSQFiVttBBISVmpb6LTy1ufCzSFvCXHamL+E23ryDh607/tPzwpSiuuhNZd7qe1IvBDl/a
sR3tMMui73Pyp0Iak8GnNnwcPmo25Jg/jY89N/1QLVgS4a7V9bOKUkglyAP7rmqRwL2N3KFxc3Q6
m7kMC5kqbTBxK3n/Fk2OGpe00BTn6No+8tfwuqBArIKsexVcnDHF4DXgCLcSPeU4ppcLXyoMRQvW
qyvAJYfv+pL930qSLVaq7IQ2F7z94JWfZPv1I1D8TkvZP0PA1qCoXzyuD5TK0NBPGEHcB29EhmDi
wYjqdwB3XEbZt8XSVLOMmKKzEIr4olsEyXue4PH9KoGVyBHjyVanMIlH2XrvlTxaQm728lGzbf4R
Ibtl6V3SvmrBfv+azZQN3S9fF7pCbLxGYxefv/Eq0t7DduLTUFdDLRsVzsXIYfdjJYP761J8dQvg
gI/WPXvQY6MVa0wfxu7hLD9ISZ1dWLooGLsenaqoaZc4P1dRbLR7kWYpC3KXllvOEtmvXzo3Rjgw
AqDD/MAFY9gUBC6A93XMziKh5YasJVW0vAPVIV6cd/QasmeYqHPcoa54Sok4yuILeK8f2T/WX2Rb
GSBK4fJ2DEj3OMrqbglguH6HTseQG+1MBqWgBX5ZIkhR4r1EH0JsH7hU2sHtbvlUD2yXCzQaKI1h
l0c3mz3jVr6JyC9s4L0anQ6CeoNEz4hjOruuVT82rpU3tFMQA6u7L96Q4+kmarHtVJadHTh0u4Mt
8OLVwMZFM8O8m1PGo2IXOlUQIksci12/hfJPuzeCjIjK/ahYjdjX1C/TTNT0KnGZSyVMO2GMk3NM
mlqsb2KuJVjL8Dgb79QrTM9O6ZqsPRHKMQe4nnxfLkeM/y2s38jPEyC2ZUXPZh/a2+6jsCj4/J4l
s9rvgGpHtrJ+Npw0Sa9sEVxkaekFwvZcP/eV6uJ+jAg4eZzc8q/v5on2Ho559/pmxl1xYLAGeLtN
4nvEigQ5p6y/yQPnKGbHvAAtxZtXhbk1PvwII0n/HtofqfZsoL3+wylDs57/TY4ZsE50Bl1LjfnY
53J6XjrbQisuM5GcmSPsyCObsLtAPTlKp6aUcl/PVd+WbixdqYvS9Y7M7y5S/NmZElj/4yQqNR0f
cPptTFAj/5KVDLv34QyEI7cd2TyT9MXw/MsOo+RqcsLIl/ESf3Pg8NHd96wYKiLTyj3vDvRT40Yi
BcfZxk3MtSnCUoEA1Q1tOSVe0O+/MJRI4B27lHPmPLfIbTJDu6OL0VNQD5OKiFussAbFm5IdwFIP
Hp4mlXOCXt7xLO0gw56nIOXqnKo6QlXIJsr4ioasEaeEt06fT/1XFEn9idkc1W2HEgmZ3keL2TI5
qevJ6WsJWDZLkHKIgzJ+Ia8A9KrUFBuaps1G8XfTdhz92QHheMnU87LPPtkmIMhZ6kf1zW15ypYJ
5E6hyoXclyBsz7sh7KWfMGFEVfo+KuBUTYh4crYYoFCWSCL8XRIppK8yAfU/U6z+x3IucRATfR/r
6t2Prm2zpbNXKB1v0T5R9NA52c/mLHZQ5kOqpMGnKgeK6UYQbYxCbuqRc5ZSMftp18W+xcrfKKUH
u59Ywawra/FzbEhwcEinAUMtfFiKNapTKrmxpa79iIzkO+tQJZJQZ2J1Bw+Nc0NtCYsDb3Fj8QrY
m3AJShTI9OKpxDARC+tkQrTZqomaHj6vF0zoyJxfYfQOWVZvpfE7XGJJznW7jLW36wwUJAS3/hGr
SjxvNQSYAWAWxNZcdR05E2cFmY7T54pu3XEOzhfkM6uakI6ivDZ6jz55f0iYsfDWSkdF1Bj3vm1M
09h6Hh7ZFgYipqlVmHGcoSbfR3JjIQlz6lHWyIg2l5ul9a/R1oIWhFyy9g9hvD0ERUIqE6A0Tgsw
WpT/J1qGsAElfmr5DzNG0f2sSgtWNCwHs09OB55MCzR7e2QsUpFZNv3gYl/k6w5EnE6kM8+Lkys4
57RxhHGG6mplHB2Ay+59JodsaC4qg8wcaD3eRhHrFk2GulEvBi/KcDUsyy87vJdcWmFxiEJ2Wqo4
43XBDHMx6PbKLFg6lsv6zfHJeb2DnVrCjTCN7am1jmSsciFam3P50smRsJ4CUMRRtXl/m52Ah4xb
94hAttelfc5KkoutFqt69nbktrR1lA40BqYnw65etx3aPczXHGumsMpUZxk0uYR0iAmXunbQhOuv
+jHekmbMufSQcD5b4xbTdZMjHw20BqQcmC50mk5Q1c4knis0RYPvfQbK01X+XWj05vB3ZA/QkfYU
DRM9gx2xNvz02GbflAT+Zo7owm4dGGvc2MPN+Afowdx2eKCNVe2Rm18efKCq/C8OMYu6PLh2Ex9j
lAxRAOYV6GfAY7A6dSbJumcpTcKnmwcoR74Xp0Bdkl9+28CIL3S9U+8YaLi+jf+qB3veEqn/kB3g
3q8Ac4UTV0qqNFKhEvY8677CTJI6XX2AbbbBdRUSRkhnJYHUti3EimA3Axft9xzJGrxjnyF7rcm+
FO4vClOZ2eG1lhxaXvlzG1Ofr5I4SgEVV2cs1Es/jwnGmQyvQ4I4N4coTAKOiKsXB4xnzZlS8vws
OZBdXUsHYInwi7uVEAo+NT8ArpsYstuQ6IIKlDilySZ3R51GCg0Yw2UG+5AjL/ILzUemXUAZ8XXH
68PK7e25ZinxN41Xis2OttTYwucWeKB+BsRD0nHGG/SQrZuLJOpIsLxHaXRFYhasubdc5oTShJdA
R4Pa8teCMLAL2bPBVjTFFahR4rZcvVa8YLGEPcsCK0ZA1pnIoplL09Rjb/2LpJRVTSzbgATNZ9o5
41em/OEPKbVMVdb5IXN14H2jXgB7I83rH/vEj9QVrBSiIgGx8J1KR+nnle4mOEvuHtcbhDhMGpMR
mWTO9fA3YYLRdIDi9t2AvE+06vudRPHGZq0/DffoRgYy41VCN+a6mlk9b7xva1OzM8e9vs7/svAk
6EjrDfAU4DAFYa8FlOCfr6AqA8WuWsSp6tzRN0BQWfb5zdd98t3TSQhGDZXxUcgPLV9UXhJpFBsc
VVCJ9N9OI+D7aYHgU93DfPlS0PJiUMTbIgIP42JpGm9kSx/nBuJkto6qnbhvKVox4/pK16WwlEbm
/0ZQbZZTTmmj3oYuI99GsTbDCtqGQ7ysWXIcpi5/kMppscwrZJ7wF3Hs2EXiY2HcN2mZxKNQiRd3
E2MoYYmFos3JtDharyENSJKask8jsLLf9yBu8ZcLIA4xjXQgjNvKfdhKluqIb3q2cf2l0ffGPwR1
1okrmIMk65Db7VuBcdAcgb5ogSPGnKGlx0oMeq1TqudOd3ocrJ3lN8IkAelt8WHyDrD7A53qPR9y
UHtCUQTr/L0CFg+tNuI/51DV9DAdNoOX3wazn2kcgav7rs8RSs+nzQSdTYYEnypW5wT73HASybxr
L5fW6VLbt/xH1KLZxEu1/Zt1xIW1sFwJUgPI2QGmAqQxR6W6/CIjjYcVdjiKFo5S2vgvSnHC7DU0
BzfbfGnrdYpSZKbfE5ljHTKS7uScWAxbxqWtr0+pAqQWljKndwv1FwA31lsl51UEgiY9Qo7ZFyPn
IfvX4MkZYMlY6SM1OR9ktysyhK6Y3/f310KEo3dQ4MLKwGSN+PoAyrraNG3ckSJDYDVLRqhoccEs
9cAcu3o8SwSwhotgjPDW+ixaX2BGCmZUg4CKAj4A2UNMC4HNL0o9sLsPZeKaob1pzr7dyj8UsfYH
5m6tOMOVh1IVXWQJhwwm8ZnuJCYHafDgt8JjkrRqj71jXI9Ywvvm0qhCxtUwQBUnkDYLkDyLzRIV
h5r+WJNNYWFwuPrpM3flqTAikH7LuJy9YDaFzpP+HE6U1nOsLHtyD7GomhXMJNH41h2RmMaXfATB
DKfA59ZsnZ0LtZxZ6IY1TfXGLgOpPMqICw2fVtXEsQbHubZsXi52UO/BJj+qWs8rN8xvzNS2b44d
bZ6GrJ9sE2xBvcKduLLgNrRyzYnDHokooTNRnISK0Xb13DzlBwLk5kQE74IhlSnH77dRVx4Tg0mZ
nka1hIPYFvbbaX0o3C3g+lIWAjKNVzeYh/fJpuEVwfODTJdIS23zadOxia5lLTEHsO8+GU66qYp2
1Ba+DnFy2nPoekfwNqUCz/v+kjCW0WS05auh2XJcrQlM57XixxKhP6gQL6lVeM/XhwNStINFLTNI
wCnlWpkK0HcFvTfvgNgLbUJV+Pm0j9Zw99jhSxcjp0CLyubauHMeDt+cLzjnlqfRzMi5YIg6eBEU
fNpLBJAbhosyH+hQEqJ7whlKFV4Mt33Apmv18XyLzXgW3VlG3ZW2I6BMrxLyv36GgTWkPBpf0apd
NYFWuqBYRa/Jcw8JbuIj/07weADXAi1VP+4fIHZFMzR3bGugEdEqaQPzxifVXzS164slopA/yqIj
u1Zn7IUShzt1MLKyySSrpGXfIlR4MXM6Uq8SFDbUz3YjiYoayxonqtg8LoiWEeB7JehOXP7q8Vib
G9SVbDnfqXTcsIYamk9Z0bYddYicrZ77iPGw8CfupmDqZikh63/gY7IPtKY/uwuyvluysvEahgI4
nxRfC1rPOU35aCqoB04/XoB1pNZuZfxMLa7bbe3zrXk1eTBYU6aotVWGQLk1Z3UlCNDplAhSLYZ8
f6luPVN/arNUprs1iHzuDglTNWn9yZVX8OZq6G0BWZR4SfGcOLPZ9/fkmnoS6PC/KcgdMVe9PMPs
muLvdjqbq13AUopOzIn1SkSfy3E5PC+zxApa5JTdPXw8n9x3DDoX8E8vn3bYpDKVw/en84AhS/Nk
iy3mRsqPStmJxrR3RdjRCBBvvB5EYmDoWP5nSaamtxSzswFRbwnrZ5YCn1evmQ0abc/lDUkvBbMs
VlDtUBoXE0+eXFGygHevaayOFucq2W8WQbqNGD4nCdCoxZFoD53+Q9xV6ifzPAmowsaLjp3LszYT
OjmwYFkdKXy0wxCFov3kIJoxNgmeULgGELJRiHLWfms0qXIYcyrQto4AODwK3bm/M0Hv/ieR5ohT
a5Lehk2xIzaL7kBOTY7v4oGhqnEXggYGRfnJZa1bulk/UjsUek1KGO9/MrPg2AGj4DX9eliwXkM3
KcQ2gpbtvorK8lTk/U+0Z3Qe11FJsssouVXfXeLgAzefYVSsZeQcJ1Awp3GWq4HAg1NTRmr5ZfXD
HcZenazCjL/4AzqvUMlCq9e2w3xDgUwATASpvV+rKhG0g4Az/aKFJChU70HWiGoUuNBOrrx1rR/0
baMLnmTzsWgkjppo1jSVGdHuSYXIFacZ6gbIgXNAVhJafCKX97S+TunVjSOtR9BMULG2GS/kYjZw
nNnWdwAAn3CIDMAqkF5U+yVtIi1crDrs3F4YfhDVS6BAGVePnp8KKpa0GTmK/uXh49FvIoDU4hnV
X/7gfPNNdAYQYdCQC8uyy0DlCKgjABrT2kBureNmrTvS/v2W3kfOK556Nepbz/NDyq1grcqjRGkx
JUQf7S/+1DjfEw50Hkpfx/wXiDQ5dz9y8vWrI5bnYwsb1JsxtrbNlJfXBGygi/uTlrXat1n8YG4q
jr1c3ltKWzHcUdwCSL7rBpDaawwbC4XrZqVS92FIj683XHUhQeX8Sm7dN/tyzNZ1Fc2ZBW3Aexzo
Y79WiIpfi2BKrjBNNMP7D2wnIsBU6O1PCto3LfrARTXNs/EQfq/GKbF/u1PQGenhv6gwKVN58T7P
W7qjDwz8kW7ZX9Tqe2mWgqH71GVLROWotd9L7bxwbZXYoZjh4xkdDBhw7CvpsY8/DBlaOcNqp5ds
zhQbcCz6LWgepbcA8xPBSyof1jk5NyAfjMc7LCqc2/HBo1IjYmXyitij78UUieoea6xAuR/W0Wbk
Hobjyuh+LsoOzzzfTpv33VrzzQJvmuQDIHcnELOYRsVcxkB2dUS1fU5wPQhmBIG+Dq4uRD4M1FoS
tQDpJz+XERj8QxgbDglWA1jWksY9vDBwHnV0J1WsoCZffHXeTGzi58dmfukuzNJPaw2KbDZF03LM
bmld/N4z/sLRkdJIfS7MhjovRggvozg4ZUkqN8NYdavhZh++XYN5iqlL9hQg0VNTyrrGP4hE5d6H
wZ4n/q3yJ/TahK/mdBwB7uIPEDdJHqmxKSULhI3WIBtBZqNG/CSXIX2LGySnQxH/TrFVEQwMGUaL
ET+hDJriZyh85yc/x+PU8y5b81/BrtsRcEzWS6rfwoHtXV5gt3Bx6uS1dO0tXFtLf4M0Y+cv9yb1
AbvQB3/aklw6kzmSHO1b2yIuvDeZIXYLgu8cjg56xR1VsXmfaxsO+DtclUKx/sHoMmfE/jq1fc1f
d+oLF7tsIPLmU7Tng/t5S7zEBFrNTHIZYiUwX8888gjQI1cvHQl/4241nfkqAEdkN/XmxT3CQXKo
TkdCsja6iwyPT4CDH+HjQVFLiz+E70NBzeF1J9Y0vahNWc6ylo1TztdLN5D0puW+I0E5JmD6rUpJ
uAlm1wxMEKKvg/wXw/dZgYHS2h2Aa7oToqwUW2LuZ6rCq1SF76njCfiFdLMOzkfMc8n57CzXVimd
X6nCWePkRPZicvmwgeVYhvbZuHZ9Kk3+4olCt+22utHnuKjZEXvtWY1PfeG4SKLF5wVmdoJvkaQA
edwD8X+VAJu+f2uAmppUdB6QxtpA/H7Cit27D9EWrgY6cK8Afj6tOhmtMP6DYelog7wxV73p0PMU
CZjaoa3N7aQu8hcyYZ+V9FhCCZYKpGgAZX4Db85RWPxewzMfZRDzZpDAcA5o6EclwnrNU8uqMk90
4kGgVndSi4kud8KZfwP4mH9k0MwiDe3lCI8E7iUSpFid/pEJU9qoZKSqO7B2ubMlzSM2MJ/NXIiq
rfprmTM11nO1Clfb8NwNvTt2IWtpvwK7a38vhvRGGCdIuZmxRARDqWCuXvQO4koiC/KXW2pvObyo
absuQVd2fmpWfH0CPjIDSSCiSSVhHcVX0hs5k/jFZTG6RXSrEpb6cSeKWTyCU15llAwIk8OciE+Y
uJadNr0kK8/AEM5bqnqWtlIUCKJjYYNIgcJdvCWP/2eQIQpefpBzUDhci1OKwpHiJE6v4vDzuKtL
aQJ9aEBMtu5ZtNALc6YJrW1t3BtodR9CWYIiKRLFuTA74hnwq8G/0XPyFsqzAkuWPl20c+zZinhP
OiVZYEVyXOXveZ3B9kmXnmotnn76VCdZ2dwwqfgnadQrwllU35lPtQVTYKaIamk1AgK/zgn+qT28
EFixCPrflEhheIyAGdKpRGaDGkWvtPR5WYDCE9Gjom0dS1wbAg9j8upAyFyXHmSINT2kD4CsHo1o
kowM3rbVnEVvA6k4sZI49ST1yrVNNd55DnIPKtS+To1rNNT2RQc17GO+OHwzFHmMjGozj9+Oxw3g
46pvQDmLxpMZYqSDit1WNmC1tNFto4R86anWsEcgvhqh6ruHE2S82YSFQNRWUQZfV+Z2r55N9nAk
9QKAc2Y9Dk/dl/v/FTTDpUnqJs1yaF6JqTSMpIJooX9T+8O8JmG2UCp5NbJVZot2SQDGb893vE2T
I+AJkAqKcI5tvR/WwgBrfZ09y2VquA1eKSQmHsK6PUGwk2re8HSpHCJGvjPRAFsXr1cvzY8olgPO
CGSKFWXQ11lFDYM6mpsweIAEh0eaTUSQaolmIdeG2wJ9qBytJKMgbkbZ+1bW7BJ3ecLbEp/2lz4A
Ly5AWzgEODcZ9IfoEi/7VYiODKv490dg2Z5oTi5VKtY+GenriJwYwUlLPpGVtilgtycDjiHksyoY
QGV4K4cbZV44j0InVj6qLGoMKYWWE2m0rknrVw3W8IykiyprMKAnJzfZPG5+9RqZLIE0xTHKelgh
COoSutjtrRf6o7rFeCfPqg7dZXOyezEX8nNPqsVsR69zLYHRGRxz/QFYFKyFIkcvGLtvG1lLpO63
QBkWmVJSR3jJcAkP1dwT4GORr3rplU9UVyiqqvFPUJIoUAUNQrZm8IAVzdFn+L8XeXefSE0Ul39P
z7q7k9dF1f2RYNgjr5tf/Bli5cthvjPcesGTGFB9G24ahSV3RCZt0CYa+4VAeEm2SSuSGTQDCNck
fIzZ4V/GGOuN/pV7MX569UUGnzpZf6bdBgwSOhwAmNEEWPMcl5R2GfBQCPcnucwsBxj2KDdb5mgc
nd57XB4nfDNWSXpRu/PmF2UOPD+TxtAD12qzLU0kp5cRoZ6y+q+DtmUR5e1sSZoZ/nttA34MMVvk
3WwQreAhUbIRiviK0UxKokZG6CQE3DZfZJOEQov6Se8sBVvQhTb1Zz2sPbPax9R9prVd4dsneyWs
fj3wCjnRXwm7UMsvjuaotv2/Co9bGhVqZniEvjnFkLoXFwhp3MmK3Yb/UAlRHY4mFWs51GJWydCC
nUkfhqRc40Pd+rhwrofvsQs6YEwPPnHbd+0aWiIJbRD3jmxX8gcx/Q0HmIbKKTWJk2QV/iom+4CB
lTEMGkUFavCXvTAJYW99dRpJzR3MSDvVi/n8kj0nZrKvjLkCudwX9992IZfZbu+WUq67fKWOy4XJ
CRzpw/rtGaGzKXvQoCls3pO/ZEEBhIvcOqSZub7e5+NHsd7reV7KfTzaXIyt6aIw9YcJCOXVdRTs
VIqzaxhKqPcSoasdi65oUB3nUxvTCqBig956Z3ucLKzfLDZZ71s7FapSwHi+fzRU5HAA2s8jnIkj
ATPNxen+saUpzcmOfC/AMeeGh6YOXECeuX1MhJCYoi8DuFH0M1Zkv6eaVmKRveNwvQEjKFHDUUl7
piLIsXqXMLq7coOBNP0PU5XA5F9uIk9YMXDGd6++/D9dJasPCn6d0YyhyobxeN6+LDi9bbm8oEO7
iMwT9cOHWC5el2/OjD6AFip3//yDjGVHZ+bBBtEHpjH/lwUCS2LwQa+P5XEcpknsGc8AN/VvGOw4
ZXkFlMguazWix34/z6npiEE1UAYqT9Jusp+kV0FhtjAM8hAXyrGBsiP1dBVGfwf2gltJilVGf01I
iDFZYzc/oB4kILnyMwqLY/jzHhR/Ij7+oC2Ddh4lzaU+7xZjCoOenpbEd830vyjwUFec75+XD8Yx
5g6AOp0J1UhGTxdnPrU3utmARQYIbo8j8crLVLNa1ew3Qs5POh94RNE7WFJLRTxFy1ur5W37d4pT
ZpGjINvLE6o16rzxhvR3ZshRVTidnvrGwkuN96KRXiDJHFHcdfbiweN8EPfGEbH4v7p4kX6NHi4h
e8kvm1QjJDmjsJy1t1ScUXv6bMtpnK1y1ytRhW4aRr+MrrQyRmFNxJpsJvqG46Th2CzSeSQ6YNxy
E00mpHH/6erO6cHiQeXjKWVgiQT34IgJJ/0xRP6ZYPzc6WyEEdVDqgpX9P3eyBrlVQZ4qRLfhOrK
HJjhgvUEaR55jVxGH/o23HxQ846TCpv/O39CTDI2ssYxfm657M/IEQauE98eCv6imSX+aGmQTbAu
mzdCiOg4PwosnLtO02JEhIXWEqtCXHwWzEdxK9wX556kf2KkM4tiSdKjJ5ZA75JsIdxEqZhseAGF
olVkhq0IsOR+aZXUY83S58uaSL2P169AGIJJi54vSXIA1fX9K+sdN+sKuDQX3SoHUkcgd56l8U90
SyJRZYkZ6deHllyRLI5pOJKCKMFrbd7Vu067XGVADADZQ65G/sx7WvmiVnmL3cyO3Ix/X7MilCc6
VBeDvv9HFu8ZGTtpmimoP2gGm1TPMjb4yvmR0MqCg+DjRTBXbsUcZjPAKRkk0z24GVMpLfX/r3FD
9TRWxsMXQD5wNl5Yjxfllql30KUgolsQqkoG2cCkCGbh8KbHdN11VMVq2Vwcb2pYaV1XTQvnVXvM
r8hjDWQ68jV4qfTX6Jd/vjASClpeNELY2Y/RApX17jvORTkKUG1UqAELAqSyQeqHEFchGM3bLE/x
oUZgMeaHR2CEfnN87e7kJfiWfzB7+gTkM5NaFwYnush7CqoAlwsachBHwKw0Oq9tdH9U8v/ozkZK
8ugyePhCb/bQK7L7h4DKH2OQ3GNusWR9M9ExsIvpx+5IvccTRZKKRhLZL8qRE9WkCNH+pQPM+CLs
X7PoUydz3LbNo9PeXTbGlYT3SWmgJUVPwdzcCbGbg42CEFozYfc/2WZDuzTHrpNJiENGuWLvu7Y6
X92N3DhlyoW90ryrhFn6ZYOPrlKOUZFQkzDRZroTfLDG7B1lCsPfoh1+huxQkiAZvTkiXMP3Ua7v
Gx0R6wDUgRSI0KRtWHJ+3eRMU56m/c5yIGw4sBI/jxeORwMFoguzLvyS205umVJTypsG5THzWYNN
025uK+sLHODWupmVDjNJOGVZD8ln+ZfsfMn2XBVNIaKNmNGb11IKHbwo3GmbHgbrXDtVb4mxoVs1
yS6jBpSTPPsR1x+Y3W7DDic+mWdfbK/yzaFUSekvaJL08T1amRWsR+bsvG1g2vg4Jg9pAtut3Yu4
qIR8BQjCk/aH8l/86Hnq8X1I1paW4U4w5ojbXpm7TczaH7cgCm/h2b5QwclB6CCm4UTTVMpa64Km
IBtW1tOJC8X+IDcg2lfioB7obp+YzYdDAofr2GcUE74rqHOCbk77Ot6GjeqExZyOY9QtjWRwDcRH
Pl67YO1KFHSVfzDSCBnKCFDmHnnYztT8/k9gUK4lZgVzn2VmMcTl3RzXLCcm/cXsCUfX7O5tX7IX
nBkFUSyUfGbfwRJxK0z+HtnR74UT7XGIGPo+jLQKhp+v3hkeB+aHKc3vDkcDttdn6MjjzWUVECIk
7cGcsn1HP2qACtD/gAGuXB6R/0s1g08/FECK+ZTCEG9ohICvLViJH0twjxOQD4ipqsPqNdfDVlvG
zGJohV8v8ZqtV0PQsUEvGQoOtWXnm4yAW6jc1Ir0t+PBs6JvF6/bZCFnxsem3zF9x9XZ5Ue9GbOg
OW+zroqBjJ2K9u+UyZc7r1LrFp6h0RiTt02SRBD/Q7BSJu4eXrpTbNH3D9JMhsePsJO5LvuchOY6
o+9PXs7u6I9iG9R1+SlBFrEgEcThfOE+chXixfP6kpJ7pfmUP76IajwkUFQxtibMZn1SDZF77dJy
uYuXiFg02kXxzS8v9NN3X2MZwRIXGHH8Oaik5ZXjsfaC6EhOFL84Kj7t4L+UWJK22lISPVZQo2kT
LYC6Hg3W/ex1Bp2O1CiYD3tY0yl0qpW4ZHRqLuInu7syU9bdpX/Qtt3Xlg3UVNzgPJrr4/leijaw
R4pYi5znbrW7JNS8UhfmOqOckuxWq/18UwT4ZiXp4/YEXgUUZOe1w1S2bWZXSGYXOkvVlzgdFmQj
YE7RzU7JDXi+b8ke/87qAE0+jOp3vZlTQumaVAOxHb5uY+9zfqlxqZ7SHBMNMrtPRqPoSUJit4qB
e/XmGfuMhXc3I4JvgHaJ6km2s827NoId5o/JSehXXCi+SzS8c+JOnlKzofK/PVbIqI6AA++rzJc5
031tLoTnYQyynnRdg1obtVrvOE5tAMcRsgHLtzEQnqSYXHPI7xQ2ooMI1Qt4MkB9kCZxz+Q57Jow
HAQam2H9+Qfxkfvd3k5BOqLmNU6bgU+R0Ss9KvN+kxY9Wpx6Qx8+//FH6+MueZbxzt2E8/9t4YKc
kHyaqfYfUJX8u4uucm4EK/2yvY6bd/5WMYOoqEEKA2jHfhCv8h+WhfQvdCKAbyp6aPJxHoaFXPEB
aJyaI5iRE/UeYLU5mm8Mr0iAsMvbGcdFE3Q4da9yxLi7ESTG9UG9P2OvJIMEyvciD/mSNfwu7639
JtIwnkAtRt2ZKDcmDjmW0uWuzTkE2ySlnCsP/OE9jHaObSjf1uKMc5cl1J/lzQbV0g/mhNwBrKFI
dVO6z3WA3Ksk1yTvJKZsL8B6OMoAkoXYxNFdPI+QnCiMzxC1oJTeGGhtJrLJGUGPOgdlZ2NN2ot0
RU60D9KYkPeJdUaTq9t2WXVqlrAwKwb2gAHbDOTdX3VeM6sXRLZUElwXO4s3syksp4cpRLXo5N5V
Sh9bc/JEGEF8mD8Y80sSDc7EE5vJskzRw4Lq03HzLPVu3a2t9xCBe04Iw3HEYrkB/3latXgL7cyO
qqm0ikltXoPtG1za3iUnZosxQWmmRi+7Z8twXh+jvEtvpDQOvneBUz/haulGEcIJfrjH0plVJofB
45c+u/hIQtblIpEVM0UzBBDGYBXfTNAk1/1NMgqJ69FSTFHmi+GTBn9pSqAXAZr7quvGrwalI+Qq
TMDkpPWQhJgBNSBiFnnOmLkBLOEe/2kAyBvF/1M+DMONyB4ITT15izE7Y2of/1sRLGCJE6EFI4tS
oBTPkSKbQlSuVYtzia6EltG5M9LKQgWQvhdOz8fM/7ARTbRzREdkLBUWT4riam0wf8KdaEoJObQn
kW9kEDSLoUAL2dKJp6yJ9Mo05beem5yKbusmx+JcECsTpol0WCP4YFWGn/6N1tOvZq6V+PBJpw5Y
a1OpJ7SbpnuDuGJqfyFJPEOXVwS4qgalI1Pt1u+52z95feBZcI5iudvHBiApIOGsC5XCsxmoJwLp
VaChx/qxXDNu70RZF+Qg4Gw0cq5DnQ6+8pzDjOBFqbcYOqdSO2L46jPcu+lxenZPBYydDiVTk46h
WHCn2hSkUj8TPoaHNZFLpsnYReLW2TrUtHrA7YTfcc9cNoFhitmq54uFFB9DO0qBQqpBiPE3xwIP
DoLG2Bab/4JYVei1AjwLqeSSH13KgnmH8cuFX7L4ou58yeI0W/9Dth7p2gFdbvoTc46BRRAcViIs
qD7zPEdoyTS3vSTg+ntwscme3wDmTGxUUsGEFhtIB9alZyzAFyvPATYcQuywAjXrKBPEHmPjw7i1
cYK1UCN37E1Ss3z/XOiTHRVB4Pa/eq7EVjSPL7rWGOy23yh/WS2LMUWOncybPWIrcxXNGCse9Ucf
VUXgbBrA3daTL37BCnRNnRSBrq1PI9mTaYB3PHL+5gkZIrHA8qrBpBHJuRl/kXSZ1XtljhyXyMYb
BNQFQziTIJQ4gnuYD9Yn08iCDB34BfZlX7HMKv3Ev67V5rHYMk+0v5XzI5OYSSU79a9FadtoLwoh
R0e35q4xgP+CyzBxweMZedq079FkZtpTztvFAGbI3FyBr+aH/Eu+8AtEbRnQe0HcdJlYaNON8TpY
Wdwyq+qdBEebeHiDuB3pkfkzmfNUxPRImtKF1KypB79wfxm/c2iaQktPEFmgSG/iSh9IlH9mzhZW
w+aH1EpHg6UN1tDxys6M0kg52Jsihu45EfTwie4XLSjiAgq9jOHXxO2pDv/4hx4YkrbLpftqBUJ1
1fMZAZuEkMZG2tvmpNyUmopGB2n6YE0BRX/Ct/bKOqVOTVCShOsIxavI054aDq+eb5E+lDLc3FfX
PMUUo7Qx2ehBN8fjJmy8i27mEwUQKG6i6KovAboJuZS5yfR8/S9W1aZT7cWm5W7BSVJdU3ev6veF
0IJhDslZNel46C9s6PfniPO+0ciQCGRBgh3uIIGzCGP1WRgI7wpcrXrsaBQLj+7ZafZP0Xpt6q1G
edATeyoleTfXPRcnNCwN+IFIUjbgFFSjyG1YKtZRdIKi7UpwCmCyaPTZctLUgXWSv/SSdSBX5hl8
2lpegpRnyYasGVTWuVi6ZDUjqDz0A7UxzJoqAix0fiksMIPuuQy1cIfl2o5cQt725WKVfi62PPlD
KgK6RNxDJbjRkVfuhBWaFbOQmKbZaXeTjjIC38xQJaJxQaHp0/Eve407yHT7zpULxU+WfM4zTWI4
l76QisVEiOcLngARmaAuxzTG4o/fhyxr9vYtephRpUTOJkClMhhZo0SXQ8cDptD8PSzODvnWVjlr
2YuO/X+yv71BXY2RF9H0/24mAPF13DNQqLibkRvPOHX37FKsUt4eqJeJQtcuVlECeCTVCeoah3EF
g6SBqmMsZ8QgjG1XVZKkR5Md645g35wfWzaveB1BbZJtJSbG5kXG/k6SNy/1fjnVLgTfrbt+pu0o
rk2EXwE4iUyqAQ+NfBC5xULipjIn/mG/SOOXzEzyJjZ0fVxfFCeVl0kBamkKM4aOA4HyNkJWxEvB
OevNVuvVKVGpSN9nYyTSoIpi0B23r//NOgu2u7BbZZntV15Lfi6NT+4A417u8Qkeu+tqOfxQxbDV
g4QIn6b6qH8aslSMGzzHBQk36NlbU9MAllUMJvssdp2sINrpEDQI+A3i8pyYJ/ivw2WfWH5fPB4c
hofnR3pOdu43y1ak7I8BSreZcC3aQkCi+fBRBiqXoCVLuxdIdlginxeC4y3VE02GIXgbLe8T7mBn
RBn2WkpnsXyRFHhTRJwVRwnhM6HPCdDHybtnlQeEPV4jBDbdTno8oI4Jy1G5k3EGdTDdt0dyv2bH
LLKyQijIzE/LVw9DLgXJMB7DE0Vnf8salUxkltr8JokSeu02mauCRGos/FPcYN4I0B1B/QGUJgAj
BtUgUnQ1AuLcYHIIYT2Vtf1hS+YFgkwfNrZvymZKEmyL12XkFrHkrOY5v5F1fEqvc/7npUkowH6S
n1nh7kWyAOxMMOtRc5S+LdWa8oqYsDE36dKNr0rwa9TPRO3QAijwZqAHP2xVgIxKTW/JqQH74Dj6
szflFpm7F3Wun51BtTTm7dKzJ1ZfhIxUuGEP5xGMEdV4fKlJWHqFfwDr3n+LOUCPllHapGokSgvz
Ec/4HELSmcDTdqB1wQqyNDBfTXNvNJdcdoJvfXsuxVTX89p6VoMQrUdgp5Et3vXj8oTuXKE/1vlw
+nUDsep5Z1330b7CfuGo6GjaeOiqsUi/F9JYSIFZvllEoQnheaQARNMJ3vAaUBNcRHslGPzOcaAt
VF1aFoHu+Yg1UWOTWqTpiKKLH2Wywk6/Xbt6sQWq1h47ZXO1Zu5kqSN/RjLSRWsyr+LGJOJCe7Xx
WkTTNiwgjMtgmI6wQbPBdETD/1+lBwwHAdQhI4eXW1xhHpxNpgjmNvrThQk+eyPDJaMR4PYdGyCO
ssW0TA0qNIU2qlnyn3D3MRVdWWNqLTFMV7fo4cqPQnLX+nAMEG4ub9+/vIohB3PlKQOFzsSqWn5o
1W5P+jKbPoJ/cnHnGd6nqhSTlFEpcao/UY2IjckpfVN4pf32U2n2QkFQq3Mwt2DoWhkNA6M11hN5
2W9URxcDKPnTWj5ZmluOqX4C5HJ2e8+/St0d3dffeZ3h3H7mWMALqqU3gKWWOxGBkhxnuJEvFSQ1
OpnlnEazcyU6HyCDAxQ6KZzWfH11Srn5cfDGlA4Wnzb2fqHlqzD/VcZp1RUIfdxxiJ4Rpr9bwV8q
OIYI/9ADmoUMdbGuclenFqlYeK6oGV/uul/xurQHfgmyVYRfsxuJfLGnUEYBrFbX7IFjyvr4wHDm
KY4IvRwKXqPZiEL0aEykSwZBT79vWN+qjB5GoN9LzOfgRbKCYG7GD1ouDgbXhUJV61ljiTEcIiY+
fQfFSoVC7ZdE7hU2DQQ7+IbqRWmmLr9iNQyMfa8AmGyUDrHcF/xcr3o2JHbmVsMUcn0o4S++CbHE
bVjpm7srF81sytG9Famzm/zJZkHhH0KV5nvieM9/o83nq+jEaDOJOLx/dte3PGSD/EU9QtrO4uLR
8pS6sg8csKIxwUdtYYlFVzz40idXoIgDxawgTN+Q6ssntphjFuCKHkHX9RNkBfq4U471mMj8oWfj
tNKmY4iRc0pKkKzGpfetWEOJGkeak1K5lNxh6kPE1H6c7DM5JPsqTWT7ibiCEcHX2soPCniTpKl0
pxsLEMZjKdLI98x3kGZJ2i8+jXIlYKWmPnZzHTOLSa3Mg1c0xtdbT1h5C0Ex1oOlUOcAPMS1BsUJ
j/MkU3rWQhJHZaadt2fHwZNDN7gc3MBJ8kgcyeiBqL0m57ttfk5kWwb8AyPzVkETlw+yzNY+8fT6
gIMdPrUIxwLBZcrNL3VFBVE58rMCwNjc1ZcXiwf4RDxbaxtFuLs+a4ImfmGiLThOoJxY0sqnaWMW
+/R9gLC1AH6XEitBzzRRt0gw5YV/DHl7riKdpFVXRuYV/irc6qAu+29GTt3PXLNv/OSdUvC7VKnT
/m0z6EnOt0cMjNRou7JglDmLANAajIlCWlb1uf6l0psVdtsSF3KOy2oD/zrjHUQEQR/xgD0oz05f
7wqv3Z2hjBiHkx97rEEAujp2cNL9jpUa8yJKlv/y7f8Abk3WUjl8gKAfPAJky8AAAo0cc9nu7Lwx
QXn00JJoJUTgjIWQ7Z2JxlGxj3pDVFkhWz8BIZfbQrZq26mP6kb7DSgqxwJO2IUffniNNiklRGOG
bVkz4kGSVXZnT00HVkjGC0F4xLqgnbMI5oX1utnNfZtznNLGZK8qWZkuIZb3cNW8jpMOMZ4iQFOW
3puftgjSKHS638BwJTQ/xaZ5tKyFOzyrQGGlhlXGHHXjxS/E1jGQc/1icQEnzgJI1v7eUyfE0n+s
7dbQJKW01jrgUCS3e1ddkr1rKU3eNxmbIcIY6sjxoZOaVkWq4EOjRVFm61aEuEAkfuZZzFEgdtgg
2dillghvwmGN56xTlTaGP/7gvUZfFKffnDNsb+ehFelCqQpb+Ge/eS417Sa55rsDe6usWLXy1ONZ
p+VLSFxvtlLQ18zAur2c98uFL8Hv4IWul66eNX98Ee3bSI33mmG4rDTD9n6ojjt1vsaU7+j++raj
rztPjuR0liZxq0NK8X/7ugzsnkwalozp6izeuzNk7yYjvFg/CG5xuPnTk4snLWUXqvzMpQkoTQVV
oJVUdR2r7uPYxNInRq4hO6Bm4YRcHeyg+qG+rka32YTav5egGHGuz5Vi+DshR+PxONrBGFC8o15B
HhFIc8OKq+9uXGflSaGE+/AhPKS0zx+6ohSxgi+C5rUc1IreDIhYwPyd36Vy1EHQYJcEc69fveUx
Iudeaz9ThUSGG9Ft2KC8fDYPp0CVYf0pEq0wqaeQIA4L0c/NMgXj4T+ss8qNLKkQeMYbE3JfCErO
HIypF8qQYUF5JuCwjLIQYWL6w9LICrEwQcZHML+WXpmD03H27W4UsnRtlyg8Apdgw/Gb+Wjvct/L
pI6Pwj9V7RHgHjsorra90JXik2zFIK5oi4N7Qk4QX3CwT2mb9fyi6vtdUvbu3r3nQbXnDduHbS1P
AqETh0fhk3tXbr7okzz6ZnFKYWkP7kEGRlDCgB18aYUzrJ1AqsaR+8eV5/BCFTz4PDylxBjJ7Mlg
6xmrrB0OJHNoaI566Vjs63oV+5eziAkDUl3XwbMq63Q1kVyPgwrpLPKsVMeqMiJmVbXshERuxr6S
2goNj1dQH+T6lgYVIDPwTpYYf6kXxfZjudDuEmv1IwT9LtwlPnuWSORGYCiNGXe7pd22A6xJyRHb
drc7Ob9a7aEdLF/zykxI/R1i9XX3xESLzi0tFCfhnMjgyDuU80n2uUasvjfNXRh4IL4KPI+Di8xr
kmmfSKfEUDedrg6NSD+wcmbIWsJfaMEl+v+tdCfkHLSwSdio5VOned1lBzShrBpTwBLz6QjOQaNy
t/gGjHUVwonhlo+SKVBIq1YqmQdRSYdzWSbYyBczKwLYRhUWAply0dtJFIbl2vGwuP6Ipjd5EdAY
G6rS0A4DZoikVn/dNR7ezLJ2nn3jGmgxnwqn3uE9uwYjcWZd08+mCJxwEbK0DKB10hvRUEY/dJa2
Ml2WZEYTtJmMK/4Q7vglZAOyESGsqTWh13/dTotWCS1Yqe3w8REwGKLAGrn5hpzKHkrzXHGaxL7n
WlxuXDzG4ptbMHWhcmaAr0EJLBs5VN1s64dI4BPhueVnE6nERdnkpgkA4ssa9nt2icLyNgvc30LS
/S2quILceonkLBUvIGsdgjBu/h+LcIIKoi/5Nt4yH09xYSuil67T/KEqmSql/jPc1VMaLdGSkhwi
izE+JVqhmjzKmll0a2FydNcx2UoCk6cuvZeo0DiYdqwHwHe0xet1NJ5v3g2GQFWnQYtuW5eQ5Nz4
/eSaVPEX/3EqDxMYodtlSa7WbkcepfJg7Y2RxTMUlCV0Qo7JQGqUbEX8Yh0Nz4g92bs3JhpOtCtA
6pHD9zr5riIwSXbK4DNzJNfevMIIqRVun9QYgmuNZ7d5gX4SAY6oOPEjKArT6JKPSy7I/E1uuZhy
j1IiyDE06Q33TyKDcPe3xsOL8BWrZ/CpQGbPz9A5mQmuPy2Y2TdKKDUXt91rTBTKJxIc34GTIsvD
XPP+FBvOE4Y7QCIPcB+tcTztIH8X0PFgaLQ07+uKafWxTEq5NFxdbbAgOLjhXcxgRbg9NEuunIpC
SQ9n6xSCPopmRy7j2w+C0c0YXmdox27Re/F4m/OX5ufV3aw8edYOmT+QnL6RqGByPhnQahmiZjVK
TopkBzqLDMi8Wj8oRQoBc1hVbhcy0gLDlMJIHIEMb6VwqEQn7/x+O6VH+Ppmi4DVeotLaFiSsI/1
lgmdDD45kEeOBREwjXYUGkQpYxNcGOY3VVcK+ajo2WftrUI1fwtEmBDsDCLwVmYejQmsnSm4tQK6
6r5GeQB8IrvOD10Lm1F4seDbzsvBXEkRZreETw92uPFkz9Lsy/U2ahxXwlYiBlQtUsCCyo8zCI5U
NXf4LF7N91gfOrHFE9CypNlK6RcT47xqjg7au5/PBZvqD4Wmvm6RpcPPvoQZwrLhJFOe2Gs+Iv0X
Mwky/XAMfqAg0mGLoIlAZcXl+b8JKgBaXGhsuUSTBr/InFtM1kyBK/RVW3fjTYx/A6812171A2M6
XHl+PbUenJFz0iDJ313B5IlGckJEipEkWsPJQvwfkMuks14NOS6CfzPNhKyd4gf0T9C7CeIK6ZCT
v4YXBcuYopL2cu2geep3GeR3QFInhOoTHzSF49TT6CK8LLI9uYVFpA6C3EPO4aLCfLAjd5liy/6M
fffQDTQbZHWk3veySBhy4odzKE6U5jicsnZLQ8l73JW9tYTzxx2PdIoW9DBXXhWFstacJsYghlD8
PJk0aLswxwGAHggucAoyosbwr8C0r1M8RDGSr2d/5CzsXDG29YjOIaKEbmY/Mojqt823rxSIWp3p
C0lm7IA70NluileY52WFIaTK/ml5EwETOsvKo+meEiWuhAllmPQZsxgkKE/8bjBxPAZmAFuBYw6V
zqdHWTrtZoWKezeKboPDQlT4E4ObyFK4rm6P9Zm72gQUYfnIDSdGcnzmCnIRTAdxoKSsvGcxU+sG
bdtK9P9IL0Ga+l/4dPTZGz/w1KTQJfHntfPFh58R/20jPh8OUd2DqXwdbop5dg9omPY60anC7Xrh
LmL0Ra3961r3nkDDZp9HF4bXY+zK1RA9QdI83oJN1lkzayvNkx3q+rUASlYilf0/2QLkpQ4fys9d
pBkos6SyBh9Vmke0b/JuRbn3/r7WaEGHsRH1DYdsekvRofOeBtvfdI9FNmTnG6ocesAGnB0p7ZXW
FKx9f+31I9KJKv4mc+qTo+Z20HsARx83oxuTxibnWeSi1HEA6Q2djeMZVayupeqAaMPJk1zN1hdN
hh7reEMxhHV4vV5zmly/oklle4hKqg/HH/qHX1O53LVfN7sTJwwDdJPlc7lnmcSqbrzYNc4QC04M
Aq/mZhB2d1kf0U86yBSJPvQV26zcYWEN3MDgemPRCYikxpc6R7JweeyKX316I8SiDjllq0dIrveS
YxFj1TaXTN1NT7hbeFFMFtKjH5lJQnCu+sX53JcnIY2PiQ+f1d3/Dvt0WY9y+cyLBotTIv1dt8Ys
WRaRHLuQGRvt+SnXjT269f+3vE6Yx9xvHWBj/2S/8+coFHigkvSF6PdBNbFbWWiIRypHMa9Q0+WV
qG6pvAIdsLPHcIymGMd16vaZw3IaUlor7s7iulmfgg+66yA8EMxRiR8XAMJYtYozwfWn9KLH/E9M
+cE+OskwTOCKQ4QSqDWrVo0yIXElDFJJAetNekh2DtusvWGldb4ShxrRpM47ETyHHYrkzxH+VMEU
/cJpRfpaQkjqPo1p22S1VPvPvrgWXnRf68rYtAwEoixrGmT/4eEO4H3hTDuVPUbyhburz0YTbeYn
B5dNCmeEQlZ4qHtnnJEdthTKBavrULGhACejYULQr9pfTAJ5E54SOm6No6eWIEJTMhCfBtejhA32
rZgVr528CEJ4K7nRxaNgttD+fPxm7doZxQUk5wV3/d5P8PzrG0KYRAY2YpHr+4iuMkMtKqf40HY5
gL5ChkBeYC1ZnQ8rdTKcDDEBIUEv8RKa4qpXb/iYx8luP1M6Eawpuvulgk2FWju/XvesPc3XP9LY
tXjmwNvI2Gb1OnqhMYPuLYUdTyChkmKTIDpv4DgKBieHn++c/BvPcra5Ps1MN1dSw+bLMd6JXVnE
NYVz9eiuYtTsRIqTyRgiGGgT3ubk8hYcZclgZM4xBaZTdCa1Sc0kjsdQXo3eI/5drCVSftk8Xt7X
FHCIUVf2hZ0JUcZDoxWaTpKIyF5mHw3t9PCsTKuf1b8v4SQk0rqFGg1ipIFOcTKUar+w78CF3JiJ
AQJeNuPqZ+AxX6qAPc3oThRqnhtFnjNiDWrRRlKQ5JUo7cIS5J8WFnlaHuwfpd6tt1v8Algk6rU+
jcIFgrNu3VAHd1oBBszMa+iNs4luutLXj/Z3dSTpTa2qFMXup/EN9hvoSHn7AAYNsUXWOcDjDqiJ
zWV1ZKLKtf52sd4jFYrRuxR4qmp+bxchVC7LOZKQaACdlgUhCPeVZLvI5JZLNH63DhCEi2tRDXd1
37mNWIHYEqnraldilGqmsxZmyStrZzh8m9JzxEvuFfKSfKbxmhUf22m7niCfxFgjVz+1ni/fPWj8
sBZ+SAWSXGgicUJGo2y2ME/Gf6ncJERK9idiOHkIQmU8WCPIHXKHsqw0Q3JErnar3HwRV9a7GJOe
5Yh5Zy5ezZ8HHaWAaW9CgOHz1gx5YU8LOuEqQyPWG+My402dYoA7d0jSCnMCSpnIQRg6LSK8D20s
nbbRTH855XLF2882vhQolukfYVgx/7cy8vYLJYv7Dfxm7Co5/Afd6uka5204d8BIj5uUN6vWge/o
Owtkb/ryYzLDqTMql1+/nbElsOeM3EgAMrmCQFddBpyek9UWGj88fzyxTKYyQmrsb6G4Jxy9MSfU
15+V35kat3TzUWFnhcO0FIwoSAgHY5U5FJgkcJWQFeIpwy+PbHZAk1H+vTDG4C8y4xpwgMCjIygy
gpF+dkRjPXwbOqfWAyo7xCSGvHvUqdbxGYCsb2ww7lHapzJ3SMLZGEaTsz7wKamKvqqnXFC1Ct38
HhAoKX3s0QYMx6VW7RLh1YBgBwxil5zrOUbzNLhblljs0vIEGOPKklHZ285wkk2FrEwgBa4kQ11G
u2IzcEf8y89z37Z6UvIVIe/sgvIXY1ON9rofP6UyQBNheYWmzIW1HOLYjWhOJDD7IpSEvSMX20+k
i0W94Jqw67rP0ryjagoICzn4jOPLOPpfDs1RZBOMwx3THcM0mutm/xbgO2zX9TJPzr0BwztxB8TS
XO6BZC6FKWPv+4l03bqd+z6Ai/cTbxy9nFVldpwFlDWLQs+eLUdXmQ8/cbHDRi/coW3GqUTYNJ/W
8Ua6kjN74Hd4wHj3K9kgvWagnScvfUzbPhAeTMZeWKdI6jn3/0zg+fjPgpk0Ls/B60dCwn9s5ERl
ENHWnY1RUbnC9TxgQp7FcQvNNagwNdJ/Qt93YzE/goHRMC7R5zW3OYW9RFMtwqOVmx/TJezj9ZWb
AGCmYks995Tg1CieqkJhU5KY7SP21dFxBe1WX7WLNzBQ4TvGbPzzq85Ru95LocMa/d3/VgM8mmcb
pJvdKL2QUy9r9dYxXo5cYgrhH4vKFRuoY5zD14U/wZfj7ZTVqpkZ3ybp0WRsjWE7uDEh0gITIl9U
g+u1G+cZn9SVzuCtm+t5tkaVWJrFlHQ2p4kiBcbZ6Yzkt9IPgDGedOm0XDE54ORVa3ECCADpYP0w
Ty5GXNwz9Lom/I4aTqpGZmwwJ9YaNYIxMyFndS2vUBUAFzFW1B3S4smK2luO2m+RAXotqyWJfPzy
dctnE7h4WqYFbtzXq91XHmGCN6bTKR4D+2YOsxYIxsO87v0HS0WxIq8qNHpt+iZAPhKCive863c7
Iv7OxzPXh/wv1j2Ba3WY+OWzXBgH1D1ClGqGIIHH8l0GEhPdKoOxglPdx6hzLcgnzXSwpBKFdldT
F0HrEXBj8fCyTCWiYxZTiDmUqnLZa85Qf+XEjY5Buz4ss5qbrQbwkZw/oWTXcMlW+b4ICCEEGheV
AZjsLk9NPaVAJxopnvZzupzPdngjSwjKPirS7NJQp2bmXyDUpQrl3kaRLlF98XTo3QyhS1z9sBRd
plLLw66pvBFMlThe7YQwTKuIfXn0ElxhVJmNCezdRhbq+Ujgs/z7pdW5u2tpj8qFff1VWir/mG8l
oollvobx/+NjnR2znpe6polP1Kk8fWT/ViuBPYRHy7ZnyPHtXlPqah0l2vw6e+aN3w5YM3zdoS9f
Du26rPh8ZwcPQ2v24AxA0Z1curGrX8KFZyKmDnG0TtjCLbYmsyU2q5m4dieJHQSQFKE1b8cDd61Z
gMpuuJVMEGhyB0t8WVR6A7cVnQ/hqrInd6ZkCgG8RXEMKLC1feRN9VwF81SpDqUDodVe7eoBb5l5
WgDccv1pH7RzkP1OnETPm1XjPMjP06D7V2sERV7JGoO4yu7ZNL64WRDyq9ctG789FFxueQ2XgFuz
MjdEIkjif0sNoYWSEQdaoh7MNPDCemwzwxobHaAuBT2cE/j43EASKzORgOW2jl5huVvGKnLKMXul
aYJlg8CQNO9+RKnamcqWmq2WaoexWd69B3JsJJ8DleRUETUMLVUq+CcPRHgZtA2a34LQB7VRuqbB
uSxeyQ9bt/JqsofkMv6jGWyXzScn5h2F994H82Rcs6pbebeQHgTflpw82iUfy3eryS1Gb7adzcET
1TQ7MRDDoRZuHRaKwHWX3lRo/MTzBZOVs4B45XHfDVkiaD++ll9uzUAf9ptZnPYwuxW2iZok4PDX
dzkyrBPoCvIEgSiyW3TpqlCdgHA8dYtBS6e2LD/87R8wukMNxAQdTfPeAMKDt37iWtdEAvkA4iKC
0BmU1iFXp99xjS/oVySO4fEtb/ZQObN6pzvwAS3oKNwNrc7XCKVzcNNs+c7hosN/50lHQJYrTpxH
RHefc7VttQ4JVAZdeaQQixX2RPHp752A0Ze8MeDacre9UnkanvAdgWXzFQU/Kb45EictYfy6edwQ
JAnhmQEmV/bB9c0gXWet8hHoE4m2fR4Maw1HJ7MvrzWNwZxpSlUEaUYz9S7TwHEYCU6SlzHyIZdA
nPW7HeRAAVZ13tuR+erev3i8rRgNSddrXFFeF/hrieCmu6YjqfPhbMCRxum3xI9y9xyBTFP8gmZ2
AHmMroMm1WAsvgvm02HwapFwXWZvK+xsvKOmxDHl+0fRqNKIxVihGhqpCX9++LzPBMy3vbzLetpG
PGP18bvRYslyGb2mXzxi7lf32JAyfD2dredRX+GWkjacFQSaMNBJalXqiQEAWWA9rEw1HXjqwqmv
g8AqSSJPMsKf23Au5Fn3/2iljcXKeyxcjVErVczf+EO9vuC/GNO2MVLoU/AAfWl1dEYgkJx5W39+
PR0wXTNdUuIYdzV/WaRNG9qhZtFX0CtdE5o4SKm7iGnU3dXL9SmNUwizQaf3rQl/JxY5JiRFbjt9
g88NpJNHjXj5Ji+3zppXNHDqdJD8/NxvorqRgMXvIsa7k5dOCgL4Jb2sYrIfs0T9VSGTyNgAxw49
xj5QDWAZMZwin+0oNN93X05AR579LLlTxHzwWcPkswJ9jC/UPK6K5FVEXY3NtVy4u3cHSBTPWyr+
bpKeatf7jog0+2H0444jhsEdXdiim1TuKATXSlbfzOr0wLGE9GHNLhnMtCcDB6jb79CIj/NDLUY6
u0Jiq00lawXnfr/Nle+arQ3KfZ46yoxmBvTvjU74D73Mz1IUAFRt3gzcD5Kp5dLmkuKpdZ89X6Od
fnWerxRpHdRyII61vP5r7eI2vH7vZsl3h/6Bbo8oQhjihXZCNm2f+PT0R8LLQ+fJnPHM3YdxdmHq
d9N9xFgN0JtJnDLlJV4wfsmKRieCv1NiqcUnBYYdNjTCqqB2OXTO7I8ItLiNiXzZzGjGdsyS8Imw
POmTjIa9OEZhOVLmxyK1zVRFNc1j6hj6AKxNc9GBbbqIF7GZ3n+Kw9BQIOjqRg/djtxsp2X2d/5+
H2nxp4e7buX9kY2QA4Znsl6aKpYsRxxLPwxvvOxeHcBTiGKb5HulKLr/XZW0EsD3zE+vpdbqf2SP
gdxNAuZJatcYKJ7yOFvQyh4sKZeQxnSpbqA/f4zlXEB2tvpKmAsomjzo3IUnvwQzHxSv9blf9Lto
fMIaxw6tmMLwuFnOv+VKkVE7Lo63SEcQ1s4ygBAOblDU2UPw4pto3WrvLmzjs/yEk+xaOu/n30Rp
g5Jgx2KrkRHsQgTsOnlNeImXMgusS0CYSH8oDXxB2pDYlQBA8fhmoNsG8WJTpVDFFs3IwmpwDDVX
n5WMatrEljGgQWkFBIWyCnaZ0FsFXz5ofhZxseP2o6kQjV1MugC04tKNEiq+2uP8yykjulJeo3gs
wQO8jHw64mCUIYRROCTgnAeRcS7JVoxMTWskp621V6qa/E6nbxDab9GnzMuuH75yOE8DwadokQwQ
hARWumL9AGE0uShI5JIthla+rvWeBxOxGevblxYjFVQdZ8dESh2Nsyt8myr5WpFaX6LCQwD2Ztd4
j5JYrZUZMaJ1s7nYYQVcnv8HfQUIBTob8QvgfMHz1a7ObL00Cmy5z7pRbduQmABxD0asqkvC3VE6
2g8D4d312pgrCe8ryinS/lDoZQwpx7gMAiwwl5L3eDJGNHZN+2MESmp+CIU3xDfEcgdqpF6CtSOc
6t/g4gPSeGUUzST1ZdUThby6uzjdlMf7Oo6CVfzQiTao5BmFNvT4CrxRbENQ9tXBgF/Sf4EuhRKB
eonzIZXLSrROFXpagKMBw43nYbSs9pfcCB+TWRRetgVLk+RdDtZkwiw178FJIPFZ3nYM1NpwTIOy
ji7C7gN52HYG4CVtlFoV8Jyf3W6UoNwPuni5JGjKhdYy2d4/dvcnij6dWqxoJ3Fk2xx9tmrsfNAR
fw4milAhpMjN++7x0zZ7FNL5oiA91zax5xa0vvFUH1Up3AZME3WUbglTsjIaUevnni+FaIUfu2TG
2S8MFBBrHsxPTaog52dXB0UmdDoMlWeYuV/x/GOyaU5bKVMgt9sEaNjmG6mngOgdBbR1hIZnVYZE
PRwLKrPR6Brnal8GUDICyUdN0UwELStcx24shn8aLmkn7/QBsniECbT5ZsKaDTPg0ww7BShwO8Xr
+P2EKO1s7SwwRs8lkCNm/k58JD+W82bdWklRnSS7MmP4P8HSg2BjZtxtxnQbTEDEhnEi4jZZZjrZ
BkUW9XmzevxCadadpXG5J2weyUyuBY4tM8REKS5qCShM9aheKHD5TreF4oMka5llGwd09XmOZasY
nAu+XiCMpCzkwaGwQe/T49eHEdBnU9Edkb3YHsFjIOZQJlbE4X9TtoxopXmZTL8Ld0INH6EPd+yx
lEHXinuX1CZ6+//LbjoHspkC9Znaemgo4+/AfSwjgIgZ4s6WcL1zHhkkTdAjS/hq0kREORdR+jQk
AcEI3Fqzq7okIpRvHgUXli5y7JgG5dUV3ryYQfSyZWQaGk2sgChGuDRDxMDWrApjRj9Eioc/C8oF
iFMj3Xa3BAF3q8oFfy0szb9OEQpSaizhDY3M/iQkrK31hYe8wEwNU//TOBGJyoGeVGc1lr4tn2Lq
nj5nI7f55hqAtbg5OhDr+DBIGnihLR3iZhUCQIZtCBzNJAWHB9XCjYaTiTCxtF8SYqDwcCBMLaiA
as+UK5aaswWtDI0nDXjO6weziMv7sVc8X8fW+tBhkJuPksihTOSOKNz8Dei+kBv6u7pz4eeligE8
t2xI9RnvXPuKSzJPwNC12DIeNu5lax5/7O/I+PPTCtKb9iNqbyUNl1R4ALWLmGtlzbznnLLC6jAA
x1E33IYyjV7p1akfxrfCjkkcPAIzKzbxUMsjtU6Mp3n52ln7j1oqEeITGU5clf/QhZKOSAHldpUV
NWj1kB+8lhrIcj6tBw+sqwFmvJoEFxjQ+aKJvk7d1vCFggGTY/AqSM/r8jwNgWwIkJ6H/3Zig4YF
oMArlPFa8c2yJsttLBZZxajWg+ywO/2RpabxnFqm+rdRIS2z0mEi4V5UOX1oUuLQ2AgPjK402MDR
rKIHLunsHb+ttRdWJP9rNdFrv2m5vLjPizaacxlqdMm9jZ3A3xiUcvio7020Qp+1C+nbEqbpp3HD
9u3NuDFjxzaQcerY16bMmbzzHn+K2OCl9mvuhUWK/iw8t7wCQmDslALcy4KYyT/Vr5glaAFkVooQ
Viqj2sN+WLtvkvQ1ZdwX2TBrpytIe8LgyasJKo65qi+zZDU39NWewQLPgj0Bm6WMIgZ5V9Woiqlh
P2k0sECIYXPn2/699gqkMm9Go2XlE8E7h9Poxcr0yXql2Q712wo2fvsqGCmhv92oS7b3FCAkYb8z
Zl8dxnPefwnM9OWJ5Hs5jmmlTV8Rrf61o0o7JMt1EZDUzSOWYyVxvsg89g46dURtncZbI5lEGknX
MYaR4zdYllbC27MgUv5kuCfJNYtH00skdKMIUuxWP1tF03dsIshEnvcK1deG8Stx6SLsBqpvmX9H
vooKozy65jOki/fOK9D2gdQiBv4hIttMiiyNl6Om3ttKkeQnvvdBw4MiMZgpzz2KdefvraSJtzvl
KuFF5RmM/PuiXWuuXNkPwpc+PEVb4usfr765b2awanEej+EZQ9kAY30yrMoEpI4zFT6ubOXhD43H
K98wu494uCAIHbDLbxfjW6pImB0D50vZP8znq53V2OPx8XEgRGKOSft1E7WRzInoE4W1RVXwtd/i
kagLhOxEgBoN5VSc7sMFzcplfisnRJ8k9FImyL76ia9HoWArYyRi6keTcWwzHg73T2DoLrCwMPcE
eRZAkcQDL9r82qfA5DbdAq/MjOBnCZSNQm2XD4hMBu8tQMcemv7htJ4c9Xh4wWZh/IPgS8aY4W9h
GsDNcbRbTEGW5mdUNBN5w0enBaHPvrD2n7A92dLdnjGw0+6tABD1Dg7pSS1R+p96ynZiO+od+Byr
Qu5KAqerkbtJUUtNW2rG1cUtCEchhPOXIbp/Q4BymTBvKKbAhoqNa5Eu+Q4ML+GBmicFAKkfgLnn
WHuX6WA9OMoV+rNVsVw6THj4Lu7GcgmGG1P5Vnp+r2nPhdjpldwkgDMiKHbP9rSZYB+lR68alm/p
Rrh9+UESYctFXHNeX2rPQTSy61OjsgM9ehGU5X0Pme+ucJiJBJ0fsjdjhpxVWOn9whSC8HjlC47f
d4qWZuGy9SgQVQkBIgN3oLTQLjSHbQL0TYg544XFCQJrK8BAdpDw5/AGWr3kipu0VPXqJAGYRFD+
fMPproeFiDH39/yaGFJybjbbYGmdmU9nYvwBm7uG65EFLcT+caZ5SNqRtNuzUnwekKuwHAy8K6I2
SDvmHJ7CgmqMYt0yRNnlgPfxgydpOwfVexJH2Z9L1DiPyvwjq9vI1rO3IrKykDYaUeogkPEOi5h8
Udup3xcYnijEh0BYRrfsoip9ZvOKNMDiqPjW3HhOgh/da+jHSJJDLcfM/9W/6PCn6LpDRVmv3/GB
txBqZuEQYBSXtd5IT63bXzJiBIZibn1IZfCMX06kPcmzdkBn7aG3T9ZA0BPpeSRJKajEMEcYjhFF
Y9slY7DmBrxmzsU9slJg8oypnMHgbz15sR1Hm6i6XSJPmradfNHKY5B6w8Bb7r6Wzb1CcHhkxHgU
MbBUx9e7+FrAXG12/DUNkqYjiqnTj8krYEknxoJOgfM4iBUqegZ60FApMl0sAex+xjoZBRbZ/Pz1
+6cnWnPXLEjrUvwjejyvhsRBMRvXruuit+ckMtDyax7JOkhkfaDWMW1+bKawxi14WF5B4QVpExfT
yaAuigxCc4X9HgC6idqqyZdutpF70eTVR7shaK/XY8m5N7ENhPn6sLbufQAumrRDsZKiZ5FQSSeg
CwaI2JKKnUQkkvnspTBE31bSOxHqQ5yAY8e2dZ0BXgNCCqtW09x8MVXHJxIQrdnkbszQAqEQWY+q
eFggF4aggM6b7yWisC5P7sN018SWEjuAQMqIN3vvIL22CCUxGj/SHuDW/KUaLOKyyszLRj2YD7xn
3H5SxZ9lJUZVn9FguTVvNv1u39QnbMZINBBSmtoNPKoR6GDR2tP6co9Knx1blQvpGfo+o9qhfL9W
6pv9bkLlxsTJWcUfalDZeQAktIYSWqcmsS033E+0AZ4WX9/Gv2Bi1X0FIVlB0jS1Ng+IQ3YJkX9m
c2Wx+/UYMCX9b5FumjI18jn3PuPGDi+X78Aj5SV3FNRHxuGVq1eSLrTJmjuUS7fPytQG71ilwa+I
DJ3zDZUCHbCcW9GDm9DH3ohgEx7h4Qb48ndjr1f5BXSUUAh27lFfVpFcYTAmSaRJ6oQUbaR7KX35
1Qycv3yj0twx9UDEwKNr/tJfg96naWSJI3msfTYysoAng3+ZTB3O1LO/U+rwMU5ytYKrouAJGnju
hMeIrhFJjyZ/1wI0rG89KOuX/L0RFxb/I57WlifO28qhRS2xZvnf6x/YZF0MwyBaJ3T3FGSb/j5s
+Q8lV2L7+fy0ppA6IR/PCJhO7FNNgFaG9L1H2lXKNO4YegBo9JSq+IiXoBDUd9zQO+NiFpYOYaoB
fBuh2R2R49FR39H9DaZDuB88hMQBgZZtdWEs+AxA1p1I10ec2e0vwXmq6ukdDRanoVF2rWTeSjwT
IHgM5xofPCaD5Mv0TExPCMegSONU+GDWTLaKC85hYDMYzNm4BVgRfKhYl5G1hnM1jbeiCD5DI771
zthfOFMxj0RVVRn4Y2WvCXT4gnmR2Q42OyrartA0G0l2ZO+1ZNc7yrz+z88fLYag1b+KJ8gPRkzw
5O2OrWpCgFT/M8MMqDxTc8YCDbv8YU1qaytorZelk6UM403pgwdpcR8Wu5aZYd2ms3jzGtx+i8rM
X1bV2qV5iRjgq1D53kwZRN3wqme4kalDDBPkFuJShPC6AgE/X6abgPxAQIzHAsfUq9J7BmwGOvUu
O6br86XWWGecDwOFmccUnCytiDP9mcM+g/vYw6nRPuwrMZ5u9158yIWRdXmSlSFJm6bInI3/uR0N
Bj3/ya4A4doUE9QvlptVeh5BfzyBm39ACFFyfWcIwftwj9wQKDb/qVeeufw7MCZYI1hqfMOHk8wk
cvjAgKVdIW5f7SW5X/lcaQ6mQ5A/RAng1jzC62F/H4yRpBkQLAswZER+rUkq+WmDFSgHWjHNfRN2
PHLdsMWTVSfqaMyLQWV9k4j9bVn6/EThh511DU8qLMILNLxtcTVFFV2iAm6fVFtKGrjnpmNeK3mp
YdJxmuaHFaimH1m9DyEU2Ah8qD06bN/d6Eyzj0pCRwa0bNQl6dPkEUd7LjDkl5BTpOZDSJ0SNmak
OEYlhdOG/0t4E8NAgHa3C6WtRAh2uPGrX2PAgb8eF7siOSTW6zeVMewBKYHM8p1Q7s/Qmggfps3s
MVpIEckiBSVMhS96XVX3avXitII/qCs1pNPjvFRBIk+swKXR9bCfLFhUjYSUHmoImDdjfuLaZ7hI
fCKBLYiIv63y7t9XWRB75MFgRcLLEV4fbNSYzkfJYD1Gk2VMcjIRagWeZBAQnryzSjetRC5g1VPJ
uTTlIJx03bcxCLKiVz3V6QRptekf8ynz4jMKCwE/XICnTo4+OTKekhmTCkpdleLhuv99rhz/aPRy
yQbgRevZxptMiVbebgQS1FcStOZuB+26ylOsY7HzsPTeIKl7OvqXCb/KwBKFmaxvyAR24LeU72/s
8FuT52BrZe5TrBZO3lhn5oax9r9UG0ia0UCUuiaZ4Mcl+yRuRDxYqGx+KIbrkIg26Xeaz8tjOY+9
L3noFmpl4GRbhM53uUQGG68+gZhNJVwcQ3vOcEpdmuzuxV788it6zm+ZXhpB0mFpG6QIgV6kZe2X
wJl2j2xar1gYm0b2kxqr29eXXsHPBnTNbiIoohVfOqv/mASkBmzZMcmoyk99ug+SSxIWEaHvbosx
mBf7BL5655PfSIZM3R69jjhtEZe/MmpwCSLPrUeKZyoVYtmT97Dd5i9C4m2KNxE1MX3fssF6AEgw
uVworpoJ58l9hwcatSouXYrtODjL3lm5CP2oArpCv/e10Il2PL5kiJGEVYNb8U10/He6JEIs4Wu4
/wqR2OGe2vjKFCClpM1HgvZNs26it5wu1MNhZBC17MC3OTv5r8wPNwSjp/xuPNG0StdQpLsn9MgM
EiiS71grR4mSEj2ObqwkNV1VyRQn345hlp4N3IOlS7YbncRsv9H7DhGbntMYVWVdHDRsxhZMb7T7
q8a73Mj/oKiYsEnTimrFE9Y6TboOZiluWcL9SPYQcsnixkn6WXluCtbsEmOXnr6rmIbI1zIaa5dG
qmkaksPrkTXr6yJNv+qsqHtIZXNdCZv5JWBjS6PsZn9OZ0TaXtW4ehOrzWirfl/z5LwZuUvo4rwv
lk8t0X2o8rtaiLtLJ3JHCCYFz2ctUtAzSs8F3oR/8usJZ9ILIoLdhcS+RfJ3T7HV6IMFnh6mPpls
r35q9tLY5Vj/YGY6tOfPLW6i4tMGtmOSeuyIWaYmeK3NJWA+Sv4SyX6OzDBmtPaS8upAZpN9IQIG
s2AjjwlimU7XZTLffMiwSSwCSupFWH4KibA9adISREuzcsvlg6oV1LzOgmR9EmV6zq890ruQQ7y2
RCtZetFG9sVrJUKhMclJF+6TvOi7f5U/tvP5GrE4oE92IJbpVuLMq4wuTjKV0guVPYNN5WWs3Hg4
lfsKzl9/M1YALPFLpbUWm1oTn7GLqCUIlqBuPJPjanjfekG9MZXJLEcE+8pFA8Q/jxr4VB6LGnDM
QYeBDOOX8yX0Q3zDPFPG4V6O85Q+F9slPyhWE9MfKdnI/z3IqSPU54gjXOAuO4Md72/KJLTGGGoR
SQNKWMY6Ld7sw9tg9V0UzmOlRMmmAtJ9xoxm+tJG6XiCfecx/3Q5Rw+aeiYmoosYjFWkio8r9OPO
yLxqyfEUj0uG6PUOsKMPZ6Bd0tjIdDQ0QmY12Ta1dMop0ldJz4OvfEekLlAZd3qDryf9zYxE4kCq
LDK4U9Qb9sCttHzr3eZNc61hh22DtEXGT+L7ciGFEbkqU8x+azTiZBHKup0Ljr1VcYqUbOdzNbVX
YW4RtvhCIhbJehHBoapbq/D2iaW6WuGmKg2RQXnyPmBVdeRj3knkjIrh1ecnWpo9yvPHs3hAqqVn
TJGzhtG1yDyvp7YBRFRnnX4n25Aq7tGuvQFnXgAYQjRdXruZE588t7CMX4kdoXQAmix00TXhMxsl
59I/27oYQkYLHLtc3cGoHCvDCauyBkzl4yHwe/H4stJJG6caodVwsaBbFEKgSPHBoKRetwylue0q
ebMjFbqs7bbgvYaarUxMY7xPKJhpm6xgo5NqpBCGkI0QhPV05b7sUbzV1YmysUqmbztCLwac4Ao2
Vmhp5wWGO9gh/jm5RSoqgl42A0NB3ts14PgfI1uGN2ZVJblzL0HJio78lNNIPnq7ebzEMZGTA/vC
MM3fcMisjEw5+Y9lXTVIq7hf3RLx3tLVW+69CT0TSS+WI0zhvpS6EHoltiGJjMv5EcXs4XFebrUA
BEHnEkpr/ynPOIGds4tMguXlGjCi+/w2m/S/VZRI5OHBEHWtQr5Ul4QdrghqUcdSNw63dTsQvbMt
Zk12vQIAx2qNODibGmSIFWbJePTMOISgYg7j5q6H3ZKmoUkTGya05JH2iQraMGEQxzWCRI89HAUA
pyiybbRQ8xiA5Hn5UozKU9uhcCOREpgWRA+jkX2xhQ/dsmpJShMUSCsUrzg4uj6kSycWrwMOiRv9
2rEGZdSTJNHas0gz6OLmoaF8qgcyanyIdgQ53pMMj8GSNzzHfw9Ec9Umb/xkGaYq6UZ3x5Sy4EnO
kWU880uMWkRt5UyRD85bmB4giIN1SIS3PVM1047bwZbmKxbWq3mdKQWSfDN00g9EsMvWQoHtQFnj
hmMNEvpBXrIqlDx9LUcRjA44hx7S5xKVJDJHMATvpHWGphnnUqIlhqz6aY0+Jmwa3JmXPmqcU0OS
qZ6ipvFUjCCucmFv6e1/92vLt2mKzeRPcJLKVq55k/+S4+dVufnbycjJezbdLP2iRRUkTc/w3FLi
hZuZyS1zOG6psjbmU0P1eR/BmwcTxOG9pihYBYFHpod+jL2I5OemYZ9e4bqJdvIlMTOQbjudhCyb
ldpvBclfrQ8VidGkwzMgaFwrZUkI7Uv/azks4FReUM8KhtkcgY4kMLeyyCSRDH59vpndGzky9+x6
nJpXGXfIV5C+gjiswpEa/s7NmXjrNrOzM4yYSXAlL1mVEL3ecLY6GCXenPT64XWQE4Vh53vjiY9E
7hBaB5CHBYsGdWmfMpJQU47oTBvZYnD34x58Y/JCO3BoSMvLTtkIL9eM747blfUxkXxy65avT08H
lFAif/tKHqlKPo9QV86coF8F9jwymReIXe4RBt1SF7mx4kfcRckKFj0W5HUnEKyvSzhaWvW1N0zm
hzrhiW40yNp/TsMujB36jcm4IkjYUBpEcanRNsj2Bm8TBWVWhpauqssv23OYnrKp7ye5a7MUcsAX
yRydXyYSxeFsirUuTvgGBaEV8XAiUDd09nL6+Wi26Q4fM3YwXsgdctDnyrb47wWs9a4gtXFIlOEE
PLYqnt2nwECsUlHpQkJ+bv1+YtvB2ikl2+1G01vn3UFyciUO85NobcxQy1f12+z8vkrs5IDrNJd6
nEJQQ9hrOzgeaKmfvyTsuVexG4JfivOzphVJ4xyN0OYnVOn55il/r7PKHzo6VNFnQxB0daMyEOCI
EK0LJuIPivlZVEhxLZWk1hloXeH16BmH2WV6Sp8NpYC4Fv/BtgXzYR+tf/3VEVvNuc4CeyfCdE/S
A3ENNJ/63LcI+ZOlxQdg/YGtSZiLKw9wgeYHmPc+FVkbNpxLbxM2GPM2fiqH328YqVCxS7y9zNm9
neUAiy5U+avMXQB6OjF3kvqhKhdUqhEOMZfcMVQZRYrEFlzbzsWX90vNpTUOpB1DNLsx2a20ZZsN
/zw3AKO9TBHfAwxNvGiRyLv+ee67626cyMc9nJrMU7tyPn5LKeOspJxp+jokj/Cur6XMH6ZYJ/IT
NBP1o6Wa5Na9t41fq95Mzjm5VwpFZLiMjhMF5QHVBu2/e9fjSQzbCBvkEPaLX9z/i/brX71CLeuk
UEGPP5tkttX29hIUn++MOZAwKQI8BLyrjHiiParmM64niPcYthsFBDJVUM1OWP6xtxgkbrMGWbxE
+/NMKXAuPJfQs5nYZQhdbZmJQHcvBm31WRhTnGz/STsvaswp1zCBYq/rHkgg9b3qiG2f2y6Qv35w
6YokB3btnCodZAgcCNB5VU3iTW3++974yxCvTkaLuzmds9VmfHhSvqtUHeP83qWJ/NLhdP/0gLAO
CBuTB/LP0IGaGhX2C/tycIIFifvuy8WuuoGxexmXasaGTm1pjO0PosmHDAnAyHLuUiVG26ZHs32p
TjsDIcnOGdhzF8qrsyVWsSv76GT8atlKVs6ZC7EA/0d57bN51lrqt0CgNAPskl+XYjZ/lc1PQWBX
4TliJA8Kma2+65m8su7jY4B2aoT3QKTRhezrzv9vqA3PYdsx/eVr8x1aLKdGAdP4FbXGzFhJyc3n
FlSeUwomGXUJKmEuUn2TS9qS8Acg4DmHSES8u3kSYm/NXAExON1+PXPuElM1n+2htXgGSuE3JIwa
s/GjUYceHDqtFPS3a7qdR63ug1PQ4BjK2SuXUHZOl5WlkJwJKCIeq4qUuqzjm2A9SclfrPW971/A
g/CLA5h5ZfvYcl/t6ColCGGAgcf7l7tw2RHmXsV48xYV7Y5h/R7TZ7v1Nwfr8TontzVcAAVF92bo
ZyTX93Mcx/ycRHJyAwlYFP9rBzbDRjgBQ9QPklJxnIlyBgJGYi2hHxIPNY6VuPaK/DAR23w5kQcT
2d+9DxPikQaqbco3v1DUqgE+v9RJTGgncVhem9KHEq2FMQisp9/ft5atljhC7wFlsw5RYJ2niZxG
yJ/YngS4RzkIi5EmqlycJYbqZCsYdn8JCrozluVdIE655j1yybcAcJgkVC/HdCyXNuv/UYemiqIY
hvKvl69owI2zJTPtn/6odnyEfKIzGr6TxhB5DgIc7IxDdvXuOnpqhEaXfye3tpyNrOhIQB/P6Nmm
GGuSKYlb8xvYjHhIFLQp2yu6XSwhPUJ/OKf1mT2eznZBfB4bOsy4tb07G42K57cb58fUZU6qzLwO
/BiDomGONnTOK4NiKm1jZsJO1XaBrKPGzmP2cqnAE8WSUlSbj9RLnVsN3HiLCDguJgx5ZZU8ICuo
4KBxQgfCYTUplOiVPlzUTo+URUyRqZp0Srkwk7W9ERtYIsjdG2gpPXHV0AvRiUfBHqt0wfqa1SEl
HkLPMB0Yg3bJP1wfvyfy89Nhng6UpNJFEzpogeE73D6vup4t6GB4iaCj1Cy+IgrcoYOqjpXprknt
Dh4O1VjL3EwRv6hDciyAeXP1IdbRfNCRevLbLtELJhsZo+4o/mPs95Tog1togbQamND8TN+vzvWZ
1AXCrlUJYReUE88+6qQ/xMOmb1RmMnpmKFXwMUcsqcec2YMwiEeaLj7th942BkbcF6TSlBghiFpP
mgK90lBHXu7EfasG4UmXfF4hw1mZW16qmM4pZbNFlpfuP9a7xPwl6KtnkFRoJ0Dc4zeo7yVWV8ZI
g9UD3/vx7wSi2nz6QWUfMwBQoxIDYjOfmHk5Vb0g5jLoUtReQ6oxHL4nvsuGsEXRFjKeJUN7NG4t
it6fpwhyywzgKUrg/agOWuAHEP6F5CE0/8zDklLEk9bG5GEmkGXCnuO8LwhxwlZ2YRgk1yMWbd94
h1cAmRbetpd1vP8Si+PUAE8Coq9CvsNrh3LbLrh3RCIkL0K+WnZT09bT6IrLlS5WhB8uO0STo1fS
MXHNF0+VYbICJalrqrY/mL2yqZ01Io+5VfxASQQ+BD82L9vVs06LI9NLDQw2BG1O/g+h1BwAnV66
/a1OrdAy4N0JYkEdyO8Ukv/oa5s5B/tsPHxYgLIw9qmRM15LZyU9kRk1PdGxESF0oSLxaRS+FrHW
MiCRz2HcrpS99LEAwmIyMryI8rQUj44zcCDqi2K7Zhe7TpFxSH7eIb/I1QUEURYnzAsg0mSzYPKr
bO4ZmOi5W4RNWbDEXRaOtt6zK28NQxNB2g31V5PddHjOQhcopIS0KK+vOVRvz/lv25gPwYneucj1
Dj0FB7FO8vPek+fbFWMKFi4QPVA935RCVT9zTwabWYr8/5ifKk7UFLODnMKaINbnBU9tjYVxC0BN
ukTEDjqfQC4J/CxAq02prEVrWLdr4NNr8J57h1qVmQeJ6gq3gG7ne3zNCpvKD612ErztJMll/+NO
McHok0zBVObqtppRxPBQyMWqDMwiaoE1QwcNVwrKemcO/ui0I2arpPFBMXVPw2pcA/qYrNKDRUQ9
rBX2zUDjodcTwjzOn1Oj/68l8BbMtaeesovn5fojsYx+Y1UchYTi/ttjkgBV+tNLUbyN1lhJQnuK
EJ8L2f8Db/9T10Sj7qNknSoTSQEb54OniK1vy0TCe/VJtWAAJfdzJCsFhBNwtJOXMq7NQoTQ5Xl8
eF/Yn8wcfayx16W6q/CMSuItet6tMpEnlm604x31eUVeGMiB+8jL77tvf2AH3o5lBGceOGuokujk
omE7ee48FdiBKnK+kH/UPAbliXeSl1UA74AXA/WvdxJsA61402jn1xsXBS6vWPoNB20xKzkckRHf
G0QpA74p1L0E9Im5PESukHke+Vg5hgSK+MkN+D4vd/BwgM6n2TYgypca0FDT07Dw/ETlo4FlqR/g
3rP+bnPlg/DpOCeshiNXbnVKo75wgizO5uHjXKVKMe/5sZkVXpXt0DK0WrKm7cXSlWuWuOloKo/S
44ZIYC/pqMtypQx3Yj77HfzilTQ5LXh5dLG7MCYvDUY09Qt3jJS5PMKcJNlGpt55ABw6bzpgetne
cPJRua8+li5ugrBtQ/ls5qA1kYgbhz0I+9lXrUVR9ZWiUTrFOpGsRkJTzkosqekqImAxrGmJvdVt
vGC/bxaJpcX0EHevBV7vGwTH2h4pIqCn9TF6Ntj9/dM4Eb3hlCEDofQ66YeuH5U/p/Kjl5BXof/Q
oyHfKcusGUHXw/nFTxItWMrL4tz6EVzqhBloCHBQKXk4bhZfbHe6PXUdhQ8DmIjiFNQgtWQyP7f8
W3moPQ2cbv2m4L+HW4DiuEdJedZvup29vV84d4j9ArbFTaLUZRRSoQiWX5V6q+rjbDu8rrv0cC5B
ULoExIxv6c9clpsuybZfLcXeiKeDJ1iTfnHgNF/Rv8bUQGZgCZ51yW9ouW0kdyZeJijvnnDMWe0T
sjksoXMlHGgZ76TGMXk2dsgnJMm7b6jY4xj5Tyjv9h9MbhQZpsgsbl+E7KxLHdnOuFjKoIRM2rcy
LyqcEvufd15/hiXNsUHH7JlHF5/JwMlYzJ6za76NjEyxVJJCg1PT5rMiV19hqBCk0umhB3RXobZ/
FTcThA7lCM7SUbZ/klYxkbad55bKi+GyNCZdQUYpiGwhnO0oZ/jeMUnCADgMzF74aTxYQKN4PdPr
h/mVirYhKMazPVhyEIi1YrvFqX2i1Xt06VrGLQi7qOz0GRgk1sDVfpME8u0pfeENL3StyRvGwccM
3PiIMdmKN4ai6tl+hv0hH7HJJw8/5BoxxLivIuQ5QkrL73yf3YhL1QIH+SGqCAyo+j+mHm+HoS5x
jTRnR2cpOwOxlTW3DdYz1wnTPPlZbUiSkqnfcJF3ZhTpOv0r76cRga1IVBYQ0uL8+nE+DyvBBmJJ
5GaBaMF3Rc/hHpMR5EYHoVcCFuHP7BLYvXDk7cynqViCh3M+LHuvyU7gpB5LqGLX5tezTdOHn0bA
nJVlf+q5AdsIzPMcoahGHAcSMscuLxR1IsNR3D6OSsChcxufSAVTZRS2flfySEpFaXLqaloBzS1T
c3qEF2a6maMsw8TAExsj9ugvoO/tNTXjdXGRVOlaG1SrUx6n+fHDJUQ7sI16MLVyBsPdSN78Xm31
HsDwsiqpiLTD5K2OWEx22PZ7GcxDWB5wuVIdXOqN0VDSoyYzxiW+1IzbSGb+0witdh773ntXixdb
T5VU4k2PdW48ZWQUOacB59xvzAKmxVpKhrz/v4V2PSvn4qRBqbqhYuWxRyNji9Wk/PuMCxWXzV+E
jjX/Ipo2n9aTZzsjrhD4IdAWVsE/wXw2P1MLk3fum5KUfnkcX5h0K7d6X7rHkraD2M3QW28BcUCn
ra97GNlrJ8WT3LfGltLCDrHYjP7O+sOHzjinZ7JDA5sQVQrnBJ8e7i+5FRD9wcfuD9ERXV2XHjUf
WIlcH5sHxoCZPj4na+OHEtQWJNiffDMAb1ustLXNab87yfwDSMzm8jN9av9LPupfn9IjKBIKwAJU
GgUO4Z1wmcSyoiPepdqP6kuMzBjIR12FfwNKTDQ60bMAtGNsUbWbBQhjorHe95FSzW20SXv3Sj7D
SUYmTIDJtNuLLIsw+tplUJ+9MLc+Ban59m79QXaS/ZPdHxqAYSdreF5KK9pNUlATLTMvDVt/cneF
ukkL8NzWKxumXa0OAchttx5pbTAVvxhvheli2tJJDI1djzS0I6gml4T1YtFTQeoN+7wM2FJlP3Ij
bngML78sVXS6IXt5sUwS+sgn57X3ei3BcTaunR6dWf/pgT0rlxadt4vOg94VPegtmouccsl1iQ3a
P10eLy8FPzDFxb/7RrgGJ3/AI3zUc+3RRmeFtDVE2CJg/gRoDv9Ipfn4WAYumMiRuJPB47U/31/a
z1bUFSvkqhksiG8MEzp7mwFguA2aMwaJJfn3ik/eUlLXMhCNO2SCIgr0gsMQDwwcIhKLSy/vAjmr
QTjNCDu4ivdbasyJ7yj0Sj+fzPjCiVYeeGZ4oJs8gnVAcPJQcdBYJY+gCnYnLroxIfeyy8hZbJBY
VTHQSRjdoZzTHw2oWZ7DWd2gZzCa77l0RkyMT07MHcpLqtKFuLQ8/ryqVWglExPIlbY14T3+wMZl
M/E3JlpFWVOAFarMsBc33zeHAr9DWmbT5+86A2uOh+iwKrRYeWbkpAMZMICJiR963xJRW/jLzsoh
0OPsGmInPC37ad5L3N8lHjJ774P3gV+0pZOxeRtWYS9uoidShL6YZLKxZ6EvQEgee/y8m12odU91
gDRo7KWNH/AcG6cLPJQoDd2m3gkWMW+aJt8AH6sWCt0ZnCW+43BWEvRX61VCmM0YDpqb/6X98z8L
zlFPLJe1uYRe9tiaY/voSJ01zN5JhzamxsDInzZJPcTc6KJ14BTCOPxzDyWF+NStdXWlhGkZAZ1R
jOU6qDjFaWOXLldXuq8UkulE0oQl7zKTeRYX0mKJVi3OYRuBhNRXS09YH3Id6BzbEcNSV7wMaID9
mrgzryrJb/1QM6D2t+2qfekhUs+pAnM+naLcp3Kgy37ZDkcwB53bA9Jm317umpKad1A00Ii6rXFA
iDAl9AwBzExfywhFFRspV5cSisaEylmCe6amFl+wALYpKRjAXK+F4M7k/uspL+SaRBc2W++Iz85M
kd7CZsZub2EFJJ41DWArB8tSVgs7lRow/gLxpiQQ9qQCsAsUIZnlWLHguyX215JAX/fudsBWWWG/
IMRaiIWTqXRTZyWp4VtCMRo6gBasiF/dR4QrhBR1JPlkUFCccR1OEtbOyxEeDUCsKWmWmoMu5TZR
mi4gL9+U3i7eUNqP7JdT2SaI/ZRv9y94hIAY7G3Y7GfWdH2zOQDvR6REzJpw1AYZ1d7WCaidaSQY
mNkA2CxvrUmMwhfVFgEBywYVzAGSHJYNorstkGsWvLvkpYEp803hrSIBQRqjzj6/faI1FOgXG/KS
OeDDuQYghOoxWAMli4V8PHs1tzPBLjDah7BMiDjM64yuF/plc2F24AUCQ5B0U1YkPc7T829ANB/L
+k3fYl1U/MJP0JG57/P/ECWhS/hJ6pQnmb5PrBE7Ue9kgPrvcAgWB4dZSKqqYks2qI1gE9n1KYvg
l5YwQR8dXtw9jTJ53+pRhrxOQB1OQhymdgpH31I2Vcj87Jeaviho9V1BM0Hc5CyGC57f1R2/ZFM0
QeBIHfvmFMRGILrupLUJpDyC1zT+duJqDERVIhs3i3ny7eeSoD8Tw9BepKrYCOmpG4hoDIFp6Hcs
iBcuOdcNVmz8efeXIXzvqY4FIKpcyYScrD1OKEd/rwVFuaLMnhLItEMZo+JFNpkMF066X+EDyncw
0qSkaElJW5/vrthxrdTE02ecTzeQEL9yewJER5PgnovGTQv2s1cjwJA+ZZwtnoMg8DVPeBr5aCpN
2zEzOtBbJYcwNwCw7rufb4/jcsy3AOB05iWDHTdRAJpU9PCd9bu9IhEGxRtEV3bquIR5sPdL+VvA
R6GnNkP27xkjmaZS0z/CfYXBYvPJo+FKQoVn0ODhD4BJF24hL7Gmte6+d+fTZIYzmak6MhBqn0DP
oBf2C8IfhCRVoMcdcsYnZKKV7eSiiOvcqm/2Tg1zziGzbK3YjyfZEDJ61iH4nq/6kYHze310XoZC
pOnpEnohlVwA/MjE7Q/s6ZT0ZZcRT1MIUCkuoEPniO0JJAvMLO9++cnGUelR1z+YzE5wIQ7GtRax
xb8EQLFPBm99Ag8HyVbdjpcpoTrlkqrHeMtwKpEUxpyZ+YjR7fa8GkZuNR3U6FwjZFkwctiEfbWE
xPMVcOr5THN2H5pp/sI3puQ8a1oCiHBAkP+Ew2nzsZdL+Hw8gcRdl7vDheXD9inbvNng9N6icZAw
3CUNfu01iADdWaj330TqiB9aJJUoxI1bR1dawShrfW4Ez115fQBsrmH7rtRea3r/5pn7rd6ykgPt
q8MCPHvPAB1T7JQi8j70AesVnuV8Jl27DgslxtAJyA0/uPE/g/XJNrkskX8VZOgiM1mIAD9vcDFo
mwAd6jUrN+uHF5KrFFBlSUB54sAZQ/1kzAEo/MbluC/SjOR4uYtDu3pY8Nbg8mJaN9z4awdqB1qn
CvsyaSETVl2Q9ZJwWy7e/tfirLe8QD5ecQbO5fwVtVVgQPWvkcXAd5BAQileT8g2ROiQRAeSa5Cv
M4JS9Z7Q25p8s8QT5q3ezdxQXbPNmET1PSac4kpZd/FreEeMlEE5ixkg33PikHi8K7i2fUEdDhoJ
Nfyrwmqq0JD+4WU1phubVqfCkZJo2NlglOXCPgxcX8PJJnb34y4VUm4CrLnh50RmXsMuXI09wZUY
MXgkxqtHonb9poBrCp634Xej25jyNOLPXLBWf0RNmJalfmoR58/p/zCYMkmdQOHU6oF1bWHIZ+kR
V0JrNMVH3sXH9591r46Bo+64Ou5o95sql1YeHy6I+PRHb9va25dPhiSprSdkyW0Ezedg3gF9I0HJ
bmpXRCPt9ep5PsGPdCphhQ+f9z4d3qd5ONnxeTEM2aq7+hKv2SAaVNjMgGXvPBfIZ+wciJ31twj/
xUJ4kauC7/k+IHjN3Bjjujzsy7FvcjERGbEb5FuVgdAgxcpWJtyqpc1og2qnEDkGe2UQgW34sHfs
5FDjoI3/umLvdsntThgFm/Zjict1sEIm8rsnIv154wuooQOGaRlyFZPAYfu7y6k11jOzj3oNKqwz
cPgA1QdKYtwH6qV1+DdLZVupZYmQcwy3ZYJm8iEofv26ltetGIgDZv80MMZgN5rox809Q3Ed6eDO
K9U1oUQD8tUjFChND7saPzYm/J2It/fSJDlIVtJ45cC4RY5CtiqaXPaNsoHWBmGmdU2/5rjVV0WI
Wdw5I/Mp61GEEr5Y1YkIqk2l+H7lvZXpgChBSMHYITTamzuCmZG68zgdokcEuVS2p9ueE67ZTD/D
auXgSpOoS4q1QZFYqJqMM658YWUjI1TbgA/3TV5StmlRJtbP0pBZ0QA1USo8cQy9LQ0tz0V5rPQU
vXVKrO6042DuZdhOfHJiwTxZ8y6rXPAHF9NQCbgZcRyQi4GmRU13fKEiM4bROQjFrsYTY4ogC/sY
cPnwrdPUq9h9SlCrDe28OVbd+SXSOqTsdMVAqAXbHQGoPVKbsHy0o7oiMB/cqNheFsv+htYx7Tvs
u9W7KFVIWTGsDklTuPArIgtGnqDGhrsKQuRgQBiBMc/PJDg7lDk3HuZdUBdnEP2CaoZHpzfwFMyE
1sgXK1X5JxsrDhZdxXOETl9jihSj2+iN4wY1UWPIktspgjiI7JwwPaePGqS11rVj2Mraznl2CUIK
QYksbn4Bg3ZhyzxfoqcZCN/Ww5CclfUMoVzX8HRXU6lE6uECaUvmEE3rcrGgQCUp/+dc6GnomKOL
8JWTnnnL3SPvyc1K7ufp8+J6d5Kqf12TIJRy5u8g3IMOITa1y+Or/HYCOnWiAk3wOm3XLZHMxTZN
zT422rmrrstLWpcMokMj/pbW562/CQWF+t0qth5TfALLL6bH1kloqSdotJr1lRrmU3gHaJbIgCIV
yUfIOQixpwOyMp/ODQN5J1GSbE1MruY0CHVCxUX64HNciesPEICOfTn5iHQwlhz4wUfg81OFcR2P
6A2LUCnoTHpHzn/G0C93xRhO6GnhiN5Hw6mdt/deI8Jk2mgeJ1dVxwh/nCyGUSjQZXcwAOHh4Se6
6Fct45glp5p6H91HBTJ2+0XELKamlDiX/Ar9pwfyGV8waEQ/NRayHDVMdV3nhMu/SUl77L5cBpFG
pB0FxtaNsPBcSzD3t8qEqem1ANbsMi33F0x/Tao1ifBBTAKBXxoK23AzvjD/6hS+v5GXtvJSqQja
gnAT4m2ZZdsjnBMH+a2emqd7E0pxNzzuXops9WPz6tYu9xDJKLm2OEm1pzSpwWYpspC8ugCZUCJr
yvU9n/K5Vq+e+X80R1Ub5jP3/I4hNZqF8ZqClsZd22nRUCxn8AmiSzX4MFmvq4kqVEUF8tZGAMgj
+TtOIaWtqpVfXQ/Zf7QIVUqhdGpekgsp83vTEfd1Z9xPi+t9gOgStIToqYILpJmxcBvS88JY0+LZ
560zIk65sQm550bKJcBKW9P8oom86Gg4cpPPFre7JW35VDlFhdKJ8SihA5TrZUM8IRZ1wpgxMRi3
+FIpeOmIQu/EwkD/W4LVm89D9XCB2HdxnyBnagy1TC6/1NFrVsX75va7hZ3zKGJxilG5NUsuPoMt
qg+Xxi+tu268Rbq94/2zmV2JN806pl+Qnq5+f3xrw1QwhbcNlQqWw0khXxkdodQ6/fFkniEIOM+v
AY7xkHlyvpyBrVEPrYutUF9rPMkM704NGdRc+E08BOuk6OfLTqrHtSb+svnNRfL6hpQXoAjqYIHv
fi1fwzQMnncCL9Paeg5SFcWthZGJzOKN0oG3FapVwlyqYDeXRecU+KnILXQghbgJdTFpuRbyy11Q
io8c60qtCeXpfUOSDJ7gzdmLFJ48ScwNlvW+JiAndvcgUa0oSWuo9vP6o7wagBTjmAqEDpVkXNOY
SvXrsvnTfu2jkBsw0uAhflvse39dQqxsVS5fKgax+keTceS6gwheGxfLutG3eIad+IWeEfgQZbxj
RsqVBUeF2ywLW/FFYm9rU2qne3FiV2hOR8Ufp4rZV1dMAYNPsOuBrnkN9qfsQ805iAe2WT/4Slcx
vNPamNDvJ5CzrhZzzHzhe3Eq3cFKFfm64FWqa0z1x3RExHilvxQXndsoPdoc8Ybt/cyBA2tmgfO4
exMdkYKJhLsK9nL24rZ3+suJMBtoMEXXgbmGRe+mFbrh8JbXFvHNUG5sTZP0no1GKj/JniXCMbF2
G6RqjN8yIRh4vWYfjVBgvhLbePjiXnyRc54b7BGYizc6NRgPYj/Y+U6HpymWR/j3OzwqoWatZoUA
z8E5FV16sOEiLwgraOKj2HFBOL4mqMFAOIjgJ/shobfCw+jK61QXbVM31tfBoBe+LDUBR86i+jYA
KgbknYsln3T4cDQ2ShlMrPUDMrSqlfZKTaMDWVf9Pf38rStcVC/s2TnuM0b9ZI21pNU1gvNBPiwb
z7XVZ7bA20Cxm8MI2gh51xbLy9WjDYd/UittMAXPqwc3kKznCYLqOSii3dB4UUp7kh4mxwOPX0DN
dth4l9R9jt/pFsXfIgvQ4hz0Py8E6hrS8rXem4P2PAYGihmMhic1bnbN/XjCXOYojqcOj+kvJD9U
muWIcVI5ovZV0ATS01qzcP456621aqQE6ai+PJPC09yUoDs4nrfOUTT6dFmXZUUqF/FAoSuPhj7H
iH4wvRebPKzszfDuSt8nGLEhbE6xxzpCYOcmWySwcpdIXw86DULuylu/bwKdJvsfRQAjZjiASSVQ
suk4FNVrzF3hgTVSd3ade2ThIr8cadEfpUnqVrGo2mxVvR8Sx54aeko8qYvz81YApIIdaEe4LLyy
xZsxPrDycak5TFyVe4k8EZSiWGvKp8VTpJbwaFdJcgSx6dgJS+7dX3zF+iuo7SVa15pwQr/9q01T
wwdoimfsk+JssO0zz3GoOUDOYMUy8/hALvRNfYDQyle18W6C8BoZ0448+mB/9UY4Vn7n53L+jBTV
zgxXRJg/Ue5bX5bR/xhSHtK1fx3vLuPd2ilziODhJnco9A+KhQo84xMls9OoRxZ6QMZumnyYKzR8
MoFsiPqOp9nBDPzyG3RZgXnx3xFugOAMiCSOmU1V2QTTgGN9lLPdxmrTAClH/rCYnXNOKbG3uKta
C9z8RzrZM2RNkqij3LxbmOE2Rk3yOjgHmF1/FmURyWI+aYVusLsNdp+ywAk+B6kBmnJudIvc9R/V
3l/N3lECHw5N8eWs8YGDb3WZGyH+Xt/2lOTf2/5joYYWcx93b2LM4YQccRCqPs6iWQ3kAPAys9T3
7H7ID3R1vuVTDHneXSyNA5dcCC9CthO0m++jhaITBDV6noET7tRITJrFwBRd8VYFiaMI6qJnGhjL
7kaeWiaml4EF2bgOqt9znDglyTM+mdHYEV0oOP7fROJKXqwIZx49rTGD1Tb6dLfnCkXiUYcRWhr0
ccXfkm3mZlZA/WCpii7NQzNioz8v7n1p/U6ZqV/AePGXs33qtGUmaOlLjeFf7MSrKUYsfrZftSCd
F5ScRfScK4EhzEosuJnmrEzl1+JqIkeykgK0hB7Uou+xXuElCD1Rcm6uDLyKuTUp9+Lr5FuNiihM
zUIoWnsix/SV9n2SGTUxVULA3UI/qEJpGrV/awgFsflKo3k8UHNMZksr+s8yB7rPC19ZCrRDnq9i
QnDNKaCeEEYgLwt0bgykAJbbS8AR5t5S5ZukfDVVA5oXliEvJ6WYn5ycIBhGEKsqfXvEn/Fqn/ri
veDcDsdfJiw7QEjYBMEbP+7+Tcz/c8Ih7fotqajZ9pgU/fNrdE7vqmHnkN53gkvPZyOPupawz9ha
w4t1FTY/qfdJKm62Tp9DSa2M+ibFaLWuRrp4Nksg/gbVjZcJRclooW0j5HSEehBF+AUHIEdzDL96
EPPrZFOuJ1rihasVbkIO1GvviiETvX3rpTD/zKZU64qyKJdk/2b1RjDA5ExusSz/m/ht6i6JRd1y
As/dnQcM3gl7CB5DaZ2Zq47+058C17sh+mcuHEHEdr66C3VcWePCLEQ0pBb1GZ/ZA22fOr2f3SQu
F9CsViSEvOEIvcd/9wJ715w2cRkYAzBBSvh+smniVKSWpzoz5ebYPRW1Xz9eZc4EMLMcFEVAw8EI
6IXP+QBlvDKN4DzAiAjT/FEWaaW16x7KEyMJzZ36TB/MzquLKf11zrLl1hhh5qKNxOUzUdVYmwR7
8VvLxpWuXyv4Yc9SDi1GLaEy5RkTHXeJoCQQd2PyMQHQDI54FEdPhmYZjVdKtWdCkJT4ohNXOBHy
o6078TfxlyZwmYhxI2TqHScpW5v4Lt8wDuJXx3hiqBuv/LnaegPPiM+RN7JVO7Sd3BhBeRQFn+gG
sdenMmAia2XMuWQ21flXRC4yX6Y0R98gl1M+nDUSJQ9oYqHR3i2MB12G9t3gAOB4qHiGtM9FdfIF
q/y8x3ezw3rEOEESEKfy74085vlt3kmrFaS5081pcJlEfD36B9nXDa0fZe9qdo6zVrKqzRk/2C3T
4Zb7/yidjhFJqONH4AfEjuJ7p5zDNJcmT7FmLef8qeItwX9uz+BmmddeHTcTOotyMLBpWoo6Kmxd
fCNbqYMrvJHbnJQcRsgvJOEdA9zuLVne+SH4w7VqkF1trL9bORNflr3nhJA98jRPPt/5j1peY/ws
TjTVu8YEa5o8o4YVp8T17g9AZHtzU6PyTwU2Y5mivhdsJJ2xW3A0HYKVyFszyzVKJyKzPZrlcUI9
czcHliF0+cf/cvyhQiW2V3U8xExvv99L1ALmlu9ujTjNr1ll6EcSo1SOUCo/2AxsXCZ9Z4voJy0N
Gb+axMBULYnoEd7iRzt7YFj+aHShaYaTjJl04kyxVA7p7LnL7wcRHunTadm/6t3N9+EN1kpvgYtD
Y9u0Rw+q4TaJUiDOBX3nebr6MByVOD2xbaIlbfbnzCPVluJtaMEI6EPm3Ag1syGb8Uju5Q+UC8Ct
3wyEvSpbPQ9fHFIt+jhrDDpyeHZVDRZjF336/XQXbK3BA1DHPz2V3pbUF7G7u6J+MrBTVwhXovFd
mHsZ+oJVje7dPBS0L8c3n7++UvDN25q2nUGziiOaZ5MKyng0B4IEv+83i03OeUSucKjCkgecJbSy
TUFbO1ZVuBeX7ZDYSCeiAdWbdu/268tZwrwQz/kp88sMsl6J0lmNBhCmA/VBfIPgG854R8IMxRU6
HcagFBuLCdYeQZ5isct1pfEAVUoBFY0wvwXdbdcbZE5tWl3i9o2udAUOKcCdbASnK3KcodY1eEGT
MN1X8vzbqCq/HMusD1JdafyQQpkx9/y2rBQ1Nl/C5sFz3SbwrZ80bBT69pDtAwRTUGTTSfAKHsPH
aWAQyCHugedrv3i9Jb+o/XC6LGLpe3r1vSo4ZJGgNbrN/7sEE+4VGnelLSOALRR8qTcK5mLHfIH2
WnT/hfqWG+3Qhsc4cbbu8Oogx86QmU4rrQlByAGll4MIDv5S2aUoDy+8qhlBSPlAUFgHxfsua/WN
aS1y2koadY2lJy3TptN70IP6n+0ovdQAvoXr5lnczxa8zJUFzpi4aUCgaGyZIzKTb3e5Xn27ZpRe
9QJSbrJQyJKbabGqQGH7Y+Uh3tMhkptJSZExgD/a1gL2+8Ghhm0ovM8zao9nNOZnCTg2S5dhWhgW
7DB5i9hQN6w5/X996PX3EjPiwqHCVTqSPsK2IDWDCL7qL6uwUPrPLcEQlENOEnU7B+oplFJU7dF3
7zaggFaInpWK7JVSgMXsHk0WqcP/X8BGOi3OCkB5y/5vLDiTF9UBTKKWpdqbFM8WK6X0lYjzjIAt
7WGwIojdCflXjI7vhVZcMDcwTWhSvLbLs3ZUxWyWzST5kXgSWCDYqYrVbRcFZmbOyjtuuqmb5HWF
yk9JUfR3at8Cl3H0phe3tpjN1t3RpEej+2FndQt3KX00OZh09fDWUeM3duPrzwWTBKFzxFqjxYrT
n6caY8VmH5EW3MRGWw+uQmVrdZMFbGav/SvIKmnHMYVlhzvwHxXBfNbuBv5W3IeSWjW4E/8YmPpw
3sPoXF7hnnouNIyIQgHdKcnKwEUk0SbcOxQQjF8Y0PFzM4Uf7pzgTnrk/3eZoDQEU/MN9P66LLVH
qaeq+i9ylST+PWy+4d5FofuQNzU8yQZcUoZxalJEPCoW8jDq/CVwYQTzTiViG1RlSbdNM5eozqzR
BM85QcLThsjI6wzjOUvcN8V7H/D1hlOl7FNoDZiGGKGcxkhJdPWasNLg0gCoCWxPLHe9DVtgEraC
c+sR9eQ3vty77+r3ycwg5jdJ3eAmW4JcZZG3wxlGktZU2iGKlBvKdlj4ic8JrowclWkVy9X8+0Pw
5+FEFd+MgSwIs9zMhgjrYcMReAVmDRSZrHITpbhWYG59VCSxgnbp8BUZ9NlMWxErVkuW79Sow1AG
IAd70whyvnS8UJi2uWvcqAJjkuMVdG+ch/jVPPipaiU5OvvZ7V0LfCIBWcxVT9MqYsUmBQLIZqXY
yybaC/+bhnRoB9C13fNhJIV0TjF1zDvcXjccrG3XJnVBNTTXSvn+TdhQZ0lOgJCeZeo5eVMpKfaX
DDBDrIhRxLnuevzzCh3XQWKFbCWvusvijP1Akncbq2OCsH/lpyEwVi6Os0cO5C75tp2zWMEzvZVb
ciSyqfv642pC88SnXYmAbjtS0o4XkvcuPZ6NGYZn2ZV5XQBuclyKuqRcovkeFZyfUDca5yD2Vtsq
KLPIOt6nL5ZBXyaoLVoH7SUa1Oz8/ygOS7cnYNu0vDP4/SwnDa6g1Py6QNNuceVLGlWMl/2xoh6I
4zDZfcY0Q3FLqVX0bKJqpGw31v+DXT+UhutRum9pvVWIsfxsvAKRKighXRzxPcYaO8a1c7f2f9cj
c5xMNEWq0VnIEyZQkz1dz/MA8qsE12B2qWxv+wMsf6CJg3pJU3NRPdaCmNjbdnirb2IY/2wdrNmG
dQJL3GQgPB9LfpNsCeKH6hyC+6eHf/aWoOb1C/2TATVet7qqSccfnk9p3bc6qb3grYHn1j/cZPNV
OwZesdSa0MNOO4euFInpUBRweNsaxtembgBJvOMil3swGgnv5XDGQw9WZTNtdpNdm8R3llB/pUhD
U0GSZmnGFpIRlxwOL3+iRC4ZPXbR5uTXyZ2f5H5/zcYJ9TBHGtxRevMvGCBAdIyKriqyrCots4gj
GjVvBgI2M+R0E3lkMXwXnNqhIHFe4Lsf8Xqr4VeYLo7rydfKDSZ66p6vQ1H1uYbkksiPq1XvLjgB
63qwef4ZEBlawET3oHu2r2dSIS45zQ0d5HtE2idbMZjYKVPDhFKuKWNRS6XHWhUSK25ctG8FQwSP
WqJcjlAeoti3NjvROUtItzjCGa3vPu3RBoKRvo+Zbv+Ok6ls2tD+c5BBwNmRK2gZ+eAgaajvS5lL
JczwPEwQZaXYFEDEwtw+RrxVz7UVcYCy0GQtg0GOCV0iDlBXyFccwQpPVLMge526XsDThttHg+gS
HrIeLlv6RWNKXp1jzB/U16qhVUJ1IhorA7ErTrKUG6dMkaZY+3Mi67ep3r3hnLLMOY3a38hj/PvY
4JbO3mhaATMEcD/ZHUztVe9nVNQ99c1wiuTBIwYu4jyTA6j51/ZyKC3+ldbGj3ORu/QPzq/Z0D5L
0D2PbMCpRIZDlLkA+rqNcgIEgbQVfM3VUWveMC2/HUYqVTm+ek6IYXrJ2yKSlG6SGhMu+aEsX/p6
Rm9RQE5R8kqzwDSlOmlzb8dxyVVtPgRbLUZmDm6tG4S9k+tZkitOkpyHzHrXiA0Xpy77lS533M9W
3fE0rV66RXIBX7jja1TOLpQmm8C8I561h+X1nkd7lMUqKj2j0MxHYA+5k17AYMPYFNzMO1kSnwvr
zus6BzPD7vH78L3fRYOFrKHphUoE8/bxcNcVXQW/z7JR1H+qeAvufKExMHFM3KY+F92oDrppjLz6
AaOQ2p4+ZOBiqCc8mLQuWT/VVT77OhhbcM6eEBbl6rivXF2MnWe3/eYmhhKQrFzkKBoTblg0XG3P
sPXZJmvCOJXAVrMGHnnsq20E8BVrgKPTC4W1rADht97sb2s03UnpQocrTP7rYGrIIrAUv0AX1/yn
WdTqv33XECoTOa4wPZ+HoXJTyr+tYAwwjVtIASOB0Q9MQaBfWPRt3OshHrIY5M4O1d+gQE+XWUtK
PvKhgVbhpjXNRkk3WAiqOWm8JPUGwp1hZZYhkOn1FGW5Gdg+ktheFsTJyw6Lv3WA63akXkEREh85
h0h6LbMSSDtrJj5nPzHXm00zj9LyIizgXTmigAlCnZmTqQFhIuWrUxdW7h+PfQ7Jl6GnuQ6lWwWA
aHNZjnflC2dgWY+FKsF6ADO3XL9wGXc1+0HIMWiGVvvx2TWy2vWzSugQqmzv4GZnvZQavZFL6y4j
HIeJ/vvpa7OCkMmIFDgSsyPL84DPP6j1HmZq8i4jQYHE4Leui67hxhR4Wv98dV9UtgbYO4FrC0um
dTeknczixIMlEdRTP0FP59wzssdKhpyrRMDixrbhybTBT8SViMr+i1dmDfzYSCUec26u4Epntsvr
Yi2QFD8BHwL+gyQ8veFf1yasZbD+4lHLdpNDRN60WpZPD9WDUlehbehQWPNraNasJ5zyxj5MEOlT
Us0qyL+t4bL0R8DrKDUR1gxymciMRfHL/gVnBGwPH50MMg/w6XaZSxGwfcDXkxgyqe24fF3j8W55
vey2RyH+klMRf/LvBsfzzWQ5VMYLA/C6P23y+Zc0vsFjfJmunGLR3btmTLKVNIpCQuALtPjg0sEt
vhoqdnLOIanuaK/K+qKxkWoFiNHcNVCaZcLohSGblUKD5WTW1TvJ34EpuHogf0aETAwgrbwxtfm6
azlrIzph7zENWSB0E/DRsxEIh58jIBOBHUOO557yH50NhRE5hJZP8ckqwYCUyAIVkC94VCxFoyBy
axgG2w4zsXAn6IlnBeLiFnkvVWeZIGsjJ4kqULZCdmOarkEpmVNGM1mghshZd+lYUcYF//X1pFHc
hKVfSuDRBdDlZAf/cuJDdvuS+h0TNJZ+8B+zkJgeMqiLCAeE7SyVzibFhQ4bSvhP3NVZqQ3alH4t
soFmRLq/Gp6djngIMmOqGosO3MtBYX3bfgSLWq4uES1JOLMuIywgkLnp8lQlcZPJas37SEmcNbNY
9Ka7OWNo634YPHmSFFkBUC+5wtUKb4E7STfvWPkO65h5KjLUeAKOxR+qkd7JCfOG+qBZcigS86Kf
yBimA8uOUv+cSU6dK3zCaWLoJ139AroY5J6KXUWXdT1ER3okKLMHlAdwLQt3TvV61A5JdrEUo2QT
oeuXW4Vav4CHOM4kR0GlUAwumRL0XS3OpEOUqIzYTVupPQzVKl+Q//+mWVqBAriZbr+Vh1c9MwKH
rhCIv/WNfQugoRe+4vTTH5Hk9IU7NsdLpczrxNXJGoBgDxVLrCUROsWo6ZHR6Nt1e+/8qD+AEExu
TlXU6qM8t2yS4pVwIw+4S6682R6CFiMoOVBDxb3GGMu0Lg9e6QipOSSlAz+ozx51ezu0thMTrU2c
4Tcm4h7FG0e00CkVS3TmWYFdAIAdeugU5EOKljRBLeGeqKW3yhIi0I3vzUtsFkM1afF27S/NvBHQ
0ciW0WtDt1sKFXHCmff04cgT1Az1i3+tYpfwKk8Xe9qJtmOSjEvGKp6HFTBH5GVid6X3wKs2rCeS
siuwMMrdc/VnyZp6MShT58ksjWAvbEG7nDGcbdZxg7SkwM5lZLkcYM3QRBApq063m9ZXF0F6icz6
PfOajYoN2VXtA8QUXL0NHnz8gozy2xeQwB4D/Vs9LJu9n8q5lAjBet8hUfnU80ETnZT9dqp91pIv
kwI9I/hzC5EEmP+Tq7w7lO2agOwkS+x+gPD1LXvnUD/Rcws1WXSWOllkCwkNWKrZwryQcVxWl6uj
LVmDL6ezOBLmD4rMEF3PSoZXF5dtWpPW2R9GBfxf3hnNExE/nQQB14hGU7bF2Av9UxjzW8QxZ3jr
YaQnD4YQyqZnLk4HZbRIN01ZS0+3YjIaZVV3TZbzAm/lP17pzTpZ1PwCGvsBk8Pn+VcUIhzwQOoz
Ry+adAVGYprmSHvTH+hfT/U4wt4Rgs5UQz+Kb1uDHQ3+NN6SoRPpgDrvl1iR/zptDu5m3sIzYkEj
j9iutZ4lb36Sg2mmU5KuI9o3N4csTO0xb+EHsxUYdmtOng9M6m+NdZxRLR2TbruMzkDGoBdJoPwu
3yNcTD/ryWWQUbro3QD72gGmiB4j4LMfyt9QaQGh9K/8peH5vaX4xrj6nBIZC2QR7maZydPXma+9
MjV/YOudzmmOKZzdWnUw0sDzydlyVYgwQOmrlr1J7sr2jOuU/zxqlSqAn1gUdNNnGFZgkQ4CnVKG
VLvJ0oX6j6WulgQEfrJtSIs9z7u+aHcMKYTvAjWLfWVLcVJxohk1XuT9mP+IwQvwY4ScmbKRYmza
ZcAvWe3IEaP6HBR5hj7POosTrQxPv+3F/JrcX3xdH3KJBxGzXxHMjxoakz2g87blhTEQmUdLijni
SXdb0G46Qz9v1vx3LxAophMFMK2sVENHfryXiacGPj1rQK8woAtbp5yA4TBA71MtpSgb5lVmJO8y
aAbj9lXYdHje4ryUF3YI7m+TuJ2uvhuvCvC1njZrAisEAzOyNcHCJ+jcrnNM1k+h5I0mTXh07CDd
GPpUt5RiC2Ja+I3Dx8c+7deNhowqVqiEcsstKtDcNnozxwV3dL82t5JXP0ee1IiPYnY2kjtIEAg5
knUpJ/Q/zfgzaLsR8TUuvqtC1R1/zslib53h6VIVAAuR/D6eH1eXY6Z6tsNfQkowfs/l+3UBFj1+
ObziY8ayhM5nLbdI7cf3RhZ3+mJBzmLLXYAdPxtR+zBJqUyVC9LcWGgypQ7qGq+tvY1tryY5IH+a
dKzzYS72yzBHkrOJA0dqL0MODUp6E67dO5bkOduaTUeDCLruLX8/BAmoksgFy6ER877i8TidELpo
7zOlm60oshLSMgiPJi4OphwGwG6iK2K6DFOSBI1uO+62rFqTQnw6ANZllFRL8oC9FoggnSSWkau5
4lrG89JH3i88vb4Funnpqo5a7YocYbwOMSV7c92A87cKekxp0uz7yVv54knozDzKQzUSbG3S1ulV
opopG9x4mtpsRGkuH+zO/BfCfoneWbYbd+EXmxjK9imF5OlhHFZ/DRCu0eOg4XhgwcTllpyJI0UX
uBSr4N0swLHiuWp23TOuO6WeaXrxW1J+T6qe+IRjllBieiWwCpE0lEmmSPlkydybKSvcE55FdmUK
/eWGZyosHMF07qpgoXD5ogL6hMtVUOcIyKKoAb47EzetwC7Q4cE4N+ef8FIbn7CPFDBkkX7IUs0l
p6Jr+15vlXDAZQiqd97ysNnJR/2jxjoLleStLK51GFsZw5ESmWR6QQggO2stjE8Gn0DswxrVDnYv
Tgk2KVGgLCPMfQEsCclxQoWb011PNF+w99XipMKcpDD6Chsc6uoWBBUrfLFVKpCWWA70jVmXaV/U
UDoGa1FyFogWwkxTbejSqiEHGmk3IR5imu8RhGE+N1YVu+qA2iFwL9ZrC/RPGMPzrjlELFkHGQAl
H6nQ9A/ASaFzhfQGRobfZcLWoGvKRhQEBaSXaduVFA5XgHWe0LEcPsUotVxN6KO52irMHC5PK11l
kGGY82SHuLSZYNCm7g66/LJJtnYxOLJ+4rJ9DwWobz+ZJ6KY0sg7cXrsXNYJaehv6+5Pz1EbFc5B
HMGHhf4PLIdiUuBcPRZOWuDoTGnNWgRqkQzS0af3jgrks+i1qlO8uM1i3ubIsGeaEQA9e929QiKK
s+X07InqtjQhNSm8hYYLKX7YE+W5i3xXXNEUsjnznJv4W2252mXwQEpRGbyZWU6+4U/ejeGYz9rA
yq+dtXOgByNZrTE1WvpIzP9hzQ+VkmmveEkssT9pDaVFYbW7aqWaJMnvd8+Hx6sfCny8UJ2ei+s2
Apwl6RNODtCRyu8hBdBcBEysc5itNkKpGDOTZot3f73TeoBGxuOa6XVJhMhUKOYMGvsN6hrPzKnI
YJVgOZVkdf+sSricNMHDO9WMIWWGICNEHi9MFP/Reiy1Y0a+B1fdad7JlSdSBAZJwPy/Fj3Hghq5
3lTtyuBbCtmZRezXgPMrhImnsMj62hNWpm/obhQT0d2YU6O/4exlZ1mX71xcJ+XePPHHYhcQ+lGT
Nrza9Jlh4nmxiDw6bx7tJL1I+4jANx+0UvJAw3bgP0aENZIQVnzoPddiJopGd8c1o9x7UHi9XpJS
351Tc7tFRstCbJDDMynA7MlmA1aHjBnGfc4a1Xi+Utql0T31KhvEDPJDjoj9/9GBwrO5H03VYeis
9g/6eL6yZLoY1NZADg0KqIFn8STNlZkdKFYvOeFoakJ9OojzsSiU61q3L6Ey7Dfeol/QGjmX+iID
bNIbBt7XAzT/YhbPejf0RDJYrbS3ezF6ftenoRrDQbdwtas/3MlG/rrdlKye8/iYoUfco0hf4x/J
VGpy12dJKPmNx3wUwBO9FlVBc8l6b6pg2AX6tkKr8LbGON2zOG6MAOayzTtuPH808tr+pSriarh8
R+Tx6CoUDDRy1ffDE5EBrgYaTaJ0eHkSG1W5ejM8cCtFJrSiTuaToPpGM0G9g7nwyhC07v5KVul+
WTucGDHWicpBvuanyZ36qMyH08GNKq2uldjDClsbRZhXqt2uE+EQ3CNILQn6pxCmW6VfFfnuhEvK
ojYdeA7pXL7GStdpD3wHOxSU/IcXG8lP2+34tQTRK3guRRQiWq/oLh31y/6oaKHkzbEGwr3N5uos
NEJRjK+t5dpiV7Obi4oS647+w0TiWo2XGcHqK2/SE5o+Hbz8d6OeSzsAzwFv/t4kn1FCfUJapkwf
Fq9ikOYo9bZMOUxuJK86y97P7IUvxxVmMrFhGZhJY6K8MSc+B3T8AbCEcWdi7cfAwchVMfb70uwi
7XIxGo9ZbXHUEbol/dmJETuZ8L042F1XWFoVJKt0Sy0xD5PoZFeR4+6Szoxk/k8sCXB8gtVCVW6J
hHAZmgdowry+6i0choYHRApRH7ELcmjmlqBFt2TtfJ1MxS086SeTwyQN3hxwVTQHzdL7Miuz06ur
iHKGJ3n1cYZX07vWWb9nYMXz6Jtn5W5z7w/8zzueNFmO8nw3IpTOKcKx3b+ngYR8l9Lh2qF5lgh5
ziuX8ReISr1pm99v5ZqxCYHRdbwO7H1kIlbLrdD/A7/8Ak7VXO/+q9yJ1mCfiLUUePDL+nmGC7TY
PRsrSykFd0s60p0D+VoUXe5rNau19yKaukp3rzZdzoarB/xRlS9ZITwgNvWHfKtZyAQebwaMa1jK
IWrDI7GgDaM8OaUf9J3HLb/2kRDGvn8RSweRhrrLlfhQzfxgCVyNYajRuzbiejeZ6GsvJxEqLfhc
59AAOA5Iq3uzgfqyvwp/JxdZwJCiAymnJkWFhzQ/Q6l3QvgWReCmaAyExhKT+/GXrsFocMs0uYRd
e1B7I6i0vdWbWdoTPpVVnjqcCSRh4okbT3kHEjFpp23cwL2b3cyHXx8ToAk3o4Cc49rbtMQfU5P9
s5iV9tDPbgu8NA16zKHrzBcBv5vyzVTnWbqS8xBAvZ2yLsjetD3Ry3w8P4DVikt+RXlmk3F5XW2y
NgN0VysWFtoYc5QvolNOpFCVYgR0MQkks4qRvwgM4mcKW6hfV+POVQf3+33iHuDnRyLEuBgrtXC8
u76b6X0Nla7lsNuBCa+FUjxC69RSEIPjVz1UhC/OBydzaoG8/TOVUYGBVfAz5TTHy/ZqPPh28T7h
tTobfh3WJygX09n1Oc/qSTlw565N9/96M9XwU5CTIQp1qRDF48F9D7Uhl9IKH/PHwlMStsHvxdKl
3fSUH4mRkYv7rUf2+lZL+Q6JY/qWFSLhwJaNRY4/sF+R4z4jEgyDjbWjeXiPHCo+oJfDwqGbOIOY
oY64ufHYEngtPEqC7woUEh33gwmPLe4nLN5k9mc79vOcuLobTyoPJ3JHa/xhVYud574qLDjRGTBB
r/oZ/AEIWaKFlDZxZhHV/VUj5U0uv15Coef8IdIGSv8/1hj3sSmqpE/Uyqo3AvccvgctHqgcyPXz
d/r15JWLLOlh2KBTC0iLxo5rE43q7kHSFH+suB/K9C8zKHI+RJIdpOLo36BtgThgJKywVha9E7wp
iP5CFQAbTgpnAIeB099ja2cDw9Soko0+XByaQT9GdjK9YM2EZ+Ol3xQ8cwHdefq8kFAnsgyI+qHS
1a2HIBVTEFhJ8hWOZUMvlUSQxY3yNyBZsMkQ3rMTJkZrajiHqKHeeYVFPeSTEc65TGF9FtUXMqLz
U2NNLq5gRYBv1YUfcJIHJL5vRLIy6Ati9RB1BmNLJrdo3bwzV32FB2ch4Q0bxHvYexqfWZeSmzue
Zvfmqr7KgRIo6weks7rFYJ6pDpLbqZMMyM1J6dLJtneMaep9Ye1c2BOLJnVSHg2nzAJKtd+cgBC5
qFUqsg3fJI2+XJnsWmlJ8mZRsE7h1Xb2ZVv5XQDx/hloYNwWlWI+WcOWoRKPmpM3ugbIBBMq/Tjo
drv2m0cBc2LV5uZmOB2HV8wzZgoxeSV+dbJaPdyWNQMAbA/HjIC1dAwwzhce3atAwjKshAIZY95M
Taz9yTn4//QvClVHfVoZF7ZGODXFaAVau6hSugQPzmh7vJwbUDA0QiIg+C0IcUR6PUtlx4QkGIST
Igvkz/PidN1nsWZVDfZzvzQjUpsu6ugfO9/XgXcngP9kRXT0H6ofY4XQTeUjWSTnja/9lg+s5coP
nSyVkHp+L11mLvgrRqIkUPHp1G7ebYMMDlwHbwiO3HHh+q/E1EHThkLWirXPtZOvMmCErZwcrT2e
pPcCzcIAb3ISCjqWcONLwdqDFWIDWSE/t1wcox6dV5p1IfaWYgVOzH4UWlvbFNVWLcSGdXl/rDVG
mcE8/C9dRBMdU1plst1U39I6b9sPnWxZby5nHuNFQavhmwA1JJFektlRF6AMBJfA+yCK0gMFhH4n
qtcrKd7Grq4KliKh10DsA8n6DEBRTzKdAkZ3orkS+TW5BlJEJ6N5XIuheF+fCH/RS2q76Xln6xy1
fSEX9CWdEEEL6kxkLsN1mnIR/wvcsZn8HTERNYdcbTjUKcy4uMGf2ki4wbrbYqcWpzuz9aBMiIDJ
i8prexHN56IReTB1vOAt5DDBtUaGZzV/kXizrsk+amMAjddWOm9rAVBPJlwQyw381Z+Ppl85E+vz
9r1ZiqQbCY1rIpkcbwvrst2SVSdWQ67cI0ZTxvn50A/z0UxS0gBqtEKkre+UusxC/W43n6xTEMGq
LQ0Mj/mpAtKX/Imgk8Jyn+IzPMqE/QuJCP2vEEcJgMqgllHBcDxCqVJYxGnRbcumTuA0EUUI0aAQ
OGKPCZtW+HXtKLrucM5c+bGFffsvnimwpYU9wVJsjNSTX9p61sRaYNmikLHMOVOI5ohiVEVPkIIP
xP3mFcwc8HREPo0txJmHhEa6VZjk7EkXyrFae08rPG61LN2hbuBcwI6vWwcxksJ0DrT++Yosxmq2
+WKuyG7cr3zARLaC3/P/LrKV0l5B71biS0tVcmHBgygPBrlUJ7UQgtUTM4AdoVgTaV5JJUrmSoVC
7DYOlETHCM0iFneuKSvExb1GHpa0i5e22htMT6CONCQacMaH4vKSKa+WZErGdVaO7c/IN7LcgXn/
8ZzjbaKZrQ/CObkTTChN/Jo8/97h9xO512aFE0RtRf8r3f9MuirpxWmA6nka1Crf05BsezNLCHzW
xvG8cKVSJ1Rw9jRg8UB8G9O/vWQJ0RpT+1/VobfnI/F9Ks11OAucFoda0+7mOPe2l8E/jvSRfuYm
ee29eTrSIRuDDf/lwwD9jj25bbSAvKH4MM7RUnWPhGFgMxv0+CbYj8pRUOgnxvA28QpBwjGzvkMK
Yl/rUpuRlEtKOAjGqRM9Utvo3aDTQ+okxWRuKyfsAAtLAffFt71JB+u88yvTvH6JcEves5i7aH76
4D74/h8LEEWaLtEB/QF2J+pg+IroQkhPbJZFPH8FMeaMj+pgjqHY2jOJAG3yRMVdonTL8g5eoHJt
fhawPbEo8Vkj6MtUzzLbpo4nYaLxa2by8Zq1heT2546SubZHqOqSckGb6R8p95a69C7HNPyEjBtP
WwSX+tyGxQcTFJ+oAW6tm+3k+UQs0qALd58JxmrIZ2QB4vGfRwXBnO04ItBzHKjyHJewT7ukLgyZ
OwN8oHgA0wZxHiKKhmUOIU+iYUyE69YAtsZLjuic327QK/yQxlxC5IbFwfcNsJEpdPPt/bR2Mr/F
ftqx3OlkJqUh7NBpWvjbtAe2N73PAufqbC5Js89SfNB4pVzb4Aw0acPa7ZLmva1fOVcc1YkB4ZLm
NZ1D85DkW4A6q2FJnQ/NzrVmHBNyE3oxhHKa6yE1ZT/qCmtWQvK7YdFyKLxs819U67ao63SoW2fj
M6XZxBnALWsqrCaOVlG41ZvJ6L22Y+uS6fx7WubafQaqRBSRTAjT1S/jcCKJlJhQ2Yn/WN7HVca4
kUDv4XHrnpCdTbWlgYDzhjKEP8DAa5HIillDh4NpXjD+4Bpgxy6XzW+KuX+GmlUGo4pzS7zDSqTd
GkKwvM/WK2C+mCeOTk07Onq+dSu8iGcvM5NmPAyJfqOh/FvsmxlouO700aniCtWpg63AYL89SKOo
NlUCXCNtHMq9+vH2/bUaWTUVVkNzRYKJ04c9JFbcrASp71qILYf4BjPsnnHiXd5x9gdmzGjHa9oQ
Fq8GQ1AIkwEitrIIiIkKqtHTDCHUUNlExfgxDFrtJHNYUGNFtirR40fvCA6EQ44IV3HAUZTjgf06
W3Pw6gYsHjKMioBjDPwNB0NXATT1L50TFZTQP7/8RL8jvkwWppNElrGtVuCiz9HpCCGrBujrXlzN
v7WQq+oIcCxTBlhashwqhDHOzhsvsAPZu3oVftM+YcZEId/PNC6/abwlB9ka/YelsoGJ4P8wRUcP
ncgQ9l3Hn7/tZX2WshczzkOoAsB7M8Nklh0x4ELX0GwxBvZX3EBGtZHNQCaI6Lrv+01Em/mAv8Wf
vs5GkSwbPYH3IE5tfkLGJB2LosBdZNGeWsbge7K2+pc+cy7vLWPUMK7etpBC6ykIHS59OccThkTc
7f7/aWTPtV5xKSCWjhaeRKMJjv7Ax8N1kTra++hpHYHkWlbbaTGalu/ZOy6LQJ/A1SpOfI5CQDjW
6Qqi3wnyaOSDEjuPBrtHxugNq+LILjwHwmnEP/Gi2jATQIcmsel1sGiZA6BeHATnkI/EG7m6v5wa
2MfRRJBgBxjPJWzNx5e9KPhV/S31CB96lWz/e7HYoR9k6itzrCC30Q5miQWu7fmCaDKOPJGFZiMl
oeONcmSGobhcrf/XfuJQb6zdU05c2ZodRNWU5VTZf2qMq+JeI5T/4KJ1LCpUpFVurP4RCRr4l7OJ
9+C0kVM7baeRjebmnfqilrh5xP+mHaRiha7uo4xOmeK0g57SPyHK4UVy6ieVxCRqgfmeMjBfFU/m
Y8NtbvbgcxGOFpfJb7WzK9CkuzRQri4sZzJ1v117+bn/h5j1tu/I0ITtSpQy4I7R4jL+HmHDg3TB
AFlQhYXX5rMGr2icNVdKtHF1U59gnCjYNXIWaGhjwGLx4fAvES3NZZW0iJhxsIPe56repWJVw1av
GIc8loqWkyP0uA7pdZwgPn1FgqwFSJlYjuIAIF5QpH+jPsJsUyZ4U9WXNxnCwVgGi4cbHg9Pt761
JFLgloSH22QvIpx6zT6cbuWj7LMCAeqWK3rNhpzaVyTZJYaeVIMzXRgZxc4Lgi3tbp3UkKRc7+1n
PH0HZsBYX6S7m2wNo1uMxgeVtwn6WbWqRoOdfydWtronmpxQur19EVgsFHbXbknVngVVej8gK3LX
TrGWUAGwfkeWkIZw2kB7TP2so6jDeqZYnP9sMk3G6aBydffaq6hygffmMX2+kUh9/YksGeU5HOWo
IjHGlRskjLN3OSv0MBN4XJhF04eYgynDL7KGoHwupOE74emPxdTi8tviWwDhYC9/8b1+m/WWKHzB
EZCKvZ1Q/UHmpLOKZP5yMM0np/YQ96SEdl84yXP5PZJaT4c7dhbtzLkPeIaAkfHuCN3buY4y81Az
mPLGsdDnahCi72auj1kBFngLikFcfWOvIhvSu9EAV5qNe19lJIrPHTsnqwtwCRMfQEw8DvJIjO2i
NF8PE977t4u17EZJbCYHnZ1UneDWKp1FQKh5JK1XwOJjs+fm7YK64HcqPFMnt2a6beQxehiqjpZd
SD6jwXexzq8eEaPTf/2d8Bduqg7243HQZ1QWidHwdvyGKf39a4LEi5Q4eHZ7NNNuavgWZGDDa7HY
/RYoILUB/zasjY7qpEC0HZmt1anm/xoHpXvmKaaeELULiT09+uuePxdutuQFprs03Nr7EVAODlz4
Wfg4rtkMVjAOluOCPcLct6T7fNrJ3qmvMlBXT0nmiBP8G/edWo0KGVwSuGtkMrRda6UniCheYGc2
EXDMe1ZgAewsUQgua2fg0x0afQge5GA3rRluNwlf7FQIPURCvle7JdKmWFC9J23R81GZATP1RPc1
NGJsLBaDpZVVIdlCa5/vzjYBmsqSP4btxZ9wNIbaWyUcspp04NBfZuOvVijUBRkqBN6mn2/GxIsR
bFYTpitMFmC77BD3Ut/IVhHcC42Gym0lasXBvtX6ft0vXuDQYode2uUrknYG0mTDa3qlIb5D+T2r
5YcIsbajMrQrggHaJx4BD4ePTZVqcYnO+YMsGSd7Vjw7mUU8VhKDbEjioT8h0afp1HNz69Q2kybA
D7+HxhOBjyctx9fL81/MSRlRMt7GfjcgHAWFlhmxJXqDIQxttBRAX9VSLGfVHn8fByiV5HIkNVaW
3OsgIs5eOTEEM48i5M63a/qEdS++OVzC5rkxMharoYch6+zGdLsGsTJyrLqGOgah5xbI7ak/LSFO
GS7o9R2UzooAOwQhOdNNGAb2bcr1z1+xIhxPw6eMxUBMuSOvFeKV2xNBBKz6wy+djn2bOF+sJlYh
4vJbSuLlH8BwEf3TeDdBYfN+LM8Mj75Wt7YsrWZpqvj1JLcLpvOTPrGlo+X0/DOAIFLqJ5mF3YPM
+BWmS71rvRz21RtS2VB+EC6BW4M1PxhnudgsSyl7ZpRPbuqEVqWihtafcOHl0yK+zyuSs1LY8BjX
+ywN5ffKwRZ0yMQj9Al2i3buhHgV30FErOkvNpdRRb0WNwIdRSqfOEYOGxzV3yS19diJE+jEZ+f2
qn+xwJOz18OiY7XHLq88yMClzW6s8OdC9/pZDamXyobfhl0ZRDSeqXaNa2eVLHJYSdeSYbPaH3DK
mC2O821BYZdVXPw7tEL7iXYuiwwwcovO8IC5zrUUuNbWX9vmN19hqISOYum5yeQ/S4r4h4e+TBIP
syEnZMhDRmkyaRunrvVrlUma2xZnvQK8qu8ZZzofHD9rJ5mnMP6x2/0zvnDFcdcrs9knma9AhwM2
iVOl31sPmh4cMbInnleoBpvmVcUwiTrKUXvVC4YMkJGWAFvecckcwdUadGSOoRpnA8ZdgukEpsF2
Vi4+m6uWRLDrGNSaErcp9pbm/WzwdY1KbZa/mSLQXEvvx5xkSJXAWmR/TWkUFLkY3RjpS/86jlnn
B3ZwJWXOFOTG9eTSp0P9CUV8YAmlFXGU5kxyUSdadyu2I0Nb5s4uAc6aIAU3qBKU+M2T3kJAuFWm
VAsdaE7PFRjBFe5VOTSFJamtVHeM1ecbTFDn8KS8fMC7Jy+DW3vwCjl7JSHXT7Pl93jsc8i/gSzQ
OkKIQfnujPbL54ugbWO9aXufLSwapyiXpZqMxTQjN5gqfBT8vVEF9X14njFPmERNCIInkv1G2kYd
f9kwGm7dkJ7LzgjExJ7Qod2B0I1mtzNZExjMg9tLHOU1M1bUiP0YsJYMogt9A3z33MWr50/8e1dg
D0QltgbpYTgujPzKL55JZLIzA2BbKnio+U8ZwH3CsOw5ZYf15g4elB22LqjuT8iU39XmSs7b6cQO
wpxt7W9GAUcIBWC1Ge5mGzqCL6tPfAnCQm+iDpGO7yYN4NqlbDIuos8o9bG5f6oguDIgS/dxFiOD
ev8V4Ezucx4AqUH2WX1SbIry/rwieq25+2MzndxuGMrRF+l5RsiP2iLXthbJTOFEAtC0Y1pLMMmZ
kWE8f/oaEcbhR6620H5WxDmuLmQTsag5QOiAsHxK6J9T1QkIjIgSVxqECcjoHhWXsuLZiDWn8VfD
G6jDn2p5xfer2a0idal13Veq8vZBze3jf45LDzb40UBZILEjYav4KWQ6yUcnMHQrcNu8+PkMryJj
UciKJtW6qf4lREYpmmPk3umdJMzlZeot2wkB2Sh1EnYRfRVFKAuurCk/YDIvsH6GMl7nFBrQWuFS
773cnZvsplbDsTsb2HdhYSgMGr/SKGbtwhFCz54TasBam5wFfRhBRQhh5CP9gEPPkAdVlJ6paNTV
vTyoJFZaPs/7MVHOB1wncpPIav3TBFWe4RkQpTjFlaSPCrNzWMbh1Mz6A346+eVHdVtA4CWB2u9M
jaU2Z8OSPHuzSdeP6sozHgrUcTSJNK1vVjMtwc9LZkf6EAlS7vGKvygEKhFq3apfJQohh6kNnLb3
egKyqocWFoso12CqIFu0+QOvdihe266eA+K+TEt3nLQ6G3fRxnR/Cjj3MSe0OcW8UU4rg5Z6Fky+
njOLVGedtWRUOjr1IWOS54LKcYHu85LF5Kthu/pBn8j0mINfGfAgpqO1wRPpJ+zycr7GaNAiEcD1
in7mGL86kceCrt2rFj/sKz568yPKDfPza8UBU+QlIXAIsLIWqvpVjaXE+jgcwNNz8Lt7czApL7MI
2WzAiFA0au28DGYsEUUWHxkBufQgTcVR0jHHzLPm2PDHC+HFpH9tsmYoI2ib+oS9Xz6K5hhZCROx
i5qBqlXaJSnDivHzuZ/lgzF2gTGWBg28DY9Wuuxrzy4PP7kruLIIDIT8Y531bdn06T4Blr/dXmjQ
p2Rt6mbKefiSgxhu6oK2afHknpIcE1hijlAHQsvXHQlbIN3oGka0kLyc9f4skYUnDWDQ7Xo2xfZs
0QqENLErsUdmk5qunK0+sveXKwoultbZqS9uBN51pkKhUYdjO38bJUe08nODj7zQuuaCRUHtRsjD
DoN181SAkCCtvKYsmL/kSvgKrHQE/BswfyeGkG7pQg0Jr2DPiapukIrknYvRegr7ZbY58K+s1fT8
c3Xhiivhb4f9/u810QmJb2Lcc8KfH2oY+1QpQoCdD20cMTqfUMbEYIUQ2+PBhSW+zvllZB8BLNQu
v/S9+JZ5graJj3FcotGb04SmUaBnMBLuEWIFGysFdH1MjoqZdeIb9vWJ1d0BBWxpqwKM0A1Kxy1Z
kaf0Gh4rbXR2DKO8o5DVPa1kwJnb6Us3o2k8++Bsw/91/XFB5TQA/k7GO7kRQvlWLMJJacBvDYB8
Ik3xhm9FleF4YxD43wwnUKTX27Wlz5KTQt/h6RQaoY1ffu13bQEaY1d71s0Nrrt1Wmu4ZVZEUE/W
WCrNS5TFWzkJgsy5vehpvxERUpwBhZtwHQaGf1UIct4fK63xGtpjqFIkgfBQ0DhTrBwGoRwLuIh9
C6fS1l/kZI4120QSz+42B+yhDgW8eroCMve5kdcZGanlvK8ZsvR4G98dRRLb46UjP+7UuKg1nxGB
3ERTLPiRw2I/cszJ7vTXNOy72PxXRsUGQ5mRIL1GIu9vRbxL3ygqr2kTPq4zz3DtcOQy6vCDV3Cq
7ZtgFsZFI9YP3ZUe2eHVikyps/au0wQOhGolOk+gHP8VCaulB4p56hm1mSbE3Mmc5wJZh3uG9b1J
DQM3qaDAiThaue4c8QyohZM92LEKB50SYbFLQnnjPYBfdckCUQy5PpjEuD9ROnRtEQY9qFN/qHxp
vYr+naoiELv9cGLOC26U8ZRnH+IDesIY94zQ/gJoydbJta8s6p4u+H32mYukvAvkd95Uq/Xmwp7W
7E6WAnZyN5jaUc7VKMBTzuNqjlkX/0HxP2JUlZPykLKcd1AF53iM+H6r0oeB7aFCiEkwqYqt3dQP
pZ1F2Ud3oAPp2CET7QR9aAPKmwMXWKokGfXsmQfJkIZBWXXoEu4oTXTAeGr6jntROsi7i0/1Q3B1
l3+ysNVpi0QvGT2uzBu0cz6Jk1N3IvZGGJ7irBS8VyhBEJmL2ax1WKNSqGcy9v0FqIY0spdXTXVM
MFqysTrbePEl2NH0wKTFiUgMtplJ/KH+N2VtPzUh+vgVX9Up5VemHD+vpdAlc9OLdfpHqtJOTTM3
v5JLBc0TncYcQZtOTzhEBf4OT46hoWJv95Zk5ISyLwtyXTb43HkioODyzMXeOkD9PW8BA1JTEpuT
3S4j7LnPFuaC/QPcuRmxQlWoVSUl9XGTCymF77ieCy1DmloK+DyLqqJdZj4eOWdmtpwHCo9gKSdK
sNS0YHS8N4jNVfEMbGfnMUM+bv1ka/jDwL0U+hbd6+5HMFpmUKKjZnfiKkcPLBezXQgjj2IxWf7s
4A5Sm7zn4TM7s4CGv5J3q3t0xD6kl9Mou3iezoUXpTG6NjrtFECyQqmRmTFwO19vJ+Mj7Y2mIC13
/snBErzKkBlFx1Z+l7o2m3o40a2L4h2UUr5rouWtFbeCQqhF386lussttFyISJ7BOINFBjNfg6RD
Cfsjgicdn74mlr6t3i5R6ANTj0vY/2s1BY5DEIAVesYzWgDYfz/YYr94n1Bwv9Svt0UfLjwQlSYE
BjnBFR+qqAaGxxoLZNMpsE4J9wEUsTSxKOTe0eYjCVodfbivTlLK/ShICG/kWOS7/ejNPcGuMQh0
XQvq1U0skMPsp9hriizKGgbUUBMx8R5ZfvsRME5zewbhZ8YdN1AM7SnAkRXtkiSAb8aUSApcNqov
Ck4YU7Lvl4bL//EO/DYiz9LXEvcI4UGtd3R79VvMmJtf7hy64IEYu00HG5/8ICFFshLe8WztGhZn
Eqqy5f2+BXU/XPMgefkeJbnZAwAChQC01dP20ToeiCsBB0+eRew0g6tmN6pu9DZm9yjFJoPfLN+j
YYiq5BMzzl35wMIP9LG8sZ4v6x+pZoLuE92Cq1iK1QB7ZzmuIuJU1vE/ocG2sGWMM47sDK6h5+YW
qdLCPQ1SCYQd7Azz4ZdAYX85ZSucx0iLG/8ZmVAZpQ4b4lAaqKdPViL5/fSjRuB5iwek2xNMwsJY
QuUcYrGQegLr/bElYJipxtHhV0rsWUsTqPWfE2DO5QCvsc9FU6nqdAtTzBnWSZbzsqGw26sPMNVP
S5yIl6KAm0VANva3KlvvGMx6WlxEEudD4TfmFaHogPpR6ahPhrGXr+Gzzz1GD9AeXafyqxICN9U6
cJospGM2sgVCc3ZMshg+VG4uP/yj/8kB8kKA4yvbyXL9nvfU3nVkA2tvAlYJUjPzUbcuSyWLWErm
XSUyZlNzWBPGYGDIF9vEqfdRKifStmKx07/45n2t75qkcFCKpLCUXu3qiG/gds27Zt2Ycx+hUDJo
p1tYsHv0/iD/xlHUcBpKXfPju+QGhu5fR4gcGEuI5r0eCK5FDglnK0l2GxkUv8ufoqsXsgkAp2is
Gnb0/ct2yiVPyVrbFHTxmqLW9aIGEAuxVd+WyXfHaX+l0tpUOBufGhLsb4UCcnT4NHDsmSfkkoem
zSw25AgJuXOTGdC0j/KAtQ7bkvydB1MCcRbU03k3Yy46/SX3nX8+SfirzouwjrR1mTcVfltd15Fg
C5bDIKB3Bl5JdPMGxYTs5k3kF3bQf5dvL6piYdnHfGUeYYM37tbLl2shc3p7KcybICa1oheNKgNh
xsPEFKS7mv4ZcPhOvX1wLoXGPpbEo12j+PEJpHT9ggTqC8MTJg8q+cISOXtnqic7wpDmixJrzQFg
9OUXnZ1qHp/KzKDvWynNT+knSADebxcX+jeySZoBo6b8Kbk7VlhZ3lhvLt+Zx5V/0tjRKUm/Jb2P
E0IBfPSDwwf4nZaqYLF1Oz8TAbHAdtCmfI+VBa8JT1Nq8h9e8JSWMT+b1NT0OfxFUJRyuP1S0E8f
HhRpAwMRNRlCchPpUbeQBeN8Nt4jd+qvtXK17Om82QkN4VMNLrNzf/Siq9ONl2s6Jfw8JBdQa/k5
QE7+yBjcj8xp+hjp8UK+IC/muuxq1/vYMc2pVn3pZpgwwMWx/Ym88qk2geFAME/ouqKfwJH0mdhM
evjbNOJ8C/oH6TomvxxG8/K5FkF/hQ3FMjG40s3l6aS+foPSiKVztYXq3Em2QmlIwhcmVmv/a7n7
WyB8pyF8wzwWK4AxFGu7HGav4a8Iv95S+Rdg70PHoiI9ODOGrhk7V9XPtScyhhimNP8WRQrjGWwO
4+siksQLfjhyJ6x1Ko/IRMXHbZ+inCtsct3AVWSZG5MebmKkXaDEW+35tBbCLpRFJOki6F/9yhB/
/InSmMvEmRgMhR5ErFHTmRk7ONX4DNDF9qOVBDpHoqM+RVK9Ib1hZ1voJTB5NIrABaCPcTl3vEh8
r9svDvZo5h1PCWvsd8Yb0pFb/pKNRn4VapBiWnACJ1FD3VCg5tTJ0GNymQAb0aBGIVEZFoLRkDiO
tc9mQSGnLEhv5B9FT5Oq0+hMOaQBW6+Cv9HnOhGb+rXBfgLL3P/7l7Gzc86X+mo8+N0d3TC9P0k3
xDyleF1L2rAZgeQlR/A43CJy5ofwMzZq0qqJ7NXs2zPHP5eypXso8qHDk9ORIGNoDWSUcJ5fol0R
lXWZJeOhr/y2nhKD6xQAU6tUKpowhpNo+Zlm9mO1CM9vtfrTuDcfwygPLT2rioDBOu7zPML26a9w
BcAtxMZFlw9WmpIX3CSblMOu90GtudyvyqSVTebCDjihX1GI/E9cWw18Sb+q01EypwVwtRIKbL0m
RhsZvDi2ftHC5d9WVn+JAIdOGdWI9VAjpXcdKYMkA8U8taeB5HNqtwaRPwX2zUb/B8PwdlfbAFq4
hvxp797TqH/+rVnxQyN/wC6h6tI28+NjDJEnhemioa5j7Zix1s9Tp2gpgsgZf+EtAYxidPco0FOz
4Aa9PDipP7feMJu1Mtm97JcMhPCnlmTIAph2rL9PpSvRpFrZhJComqaoHpQXEFQl+787RKaOOZu9
mKmEA577KppnX1Zpur8wkQzslmxzMoOCwfbr8aWPwv5r/j8bdBT+9JigT9hEgd7FfHWaFA394biW
vryoF8qyVSZdFJTJ+LxeKSCd5EZpQUHHvhmWif4+oi8EoaVNHkVRSJMFuJF19y0vIkmRhWYlkpN/
Sbtnf32603dsjmhFB7Yxm16BQo568fUb9+ouOOTSOKIvupS3Mrxhb7l0KJeBryYvWsIG+UF0qn60
Ovy+rHI32eXaHh0Vg8vDwvYJ4n0ORT1XzKM8n9ZbQ3SWtU55zcD0fpo5qpwyGrrcJGNUVrM/GVwO
L87aWcZcoGOTDvdcW0muXtQjp3sGaQKmIfVLLpONH1kQelRTnS/erzRWqQklecKfmuOdkAUshZt4
/m7ZN5IIOZfXUwsgorZbw7AY+SVI4e4aQ9IxcSna4YvES8dJHuGC+XRAxciqSh/6QOimZBekW7Rw
X8j7ufUNdFQeJSq17wXAj5BJyZxa5/E5RUEGXGKElJSV+NjzJ5KqRQW8KoIDJU59Dqp9W0wHFHcl
POj+L+hjORShjeoxjeLoePL8/CLJsDDsq4YfrkyxwwYYNSa83Tkqm+Z1eiYgNP/kHdugr4dBrGdC
MMsJlb8ynRDp127t098DfXiBZdV0NqdY3XHzeJD9Fa/WVTiwHWXB6jWVooaIGmKQXpA11/4KWpGP
forxW94GD+ZqnIc6vIYWeWDdGqx74tJjMJlASBwa2rvXqaXX/9MDmh2CFjx7pXgara5ceC9VfoaU
3UP1lbqgs0W9GvRFXIUdMFRsJytnuovy1WTl9q9CJnoytTSHuw3Y/HfcaL7RGgAb73v2cOT3i3Jg
O12nhWfzIEyCuepjjBzKHCg705B+nTlrcadpDx4GKrIGqVLgM0sjB33qzo99S/xKFM4PU+wJJq9d
RtXJzB7ocjK7FuFzaViUVMQcMb+rZQo4avL6b93WVLqIKiQNVz3WVx5frUi0uY3LBRoVLEBRyjDg
+WmEi48aTSWeyJEWUimVMo+gQvIP+ZyJ/WOB/GloLwntx+/rJxwAAW7QPA4zW92bmmtqHrtagcLf
5RDfyx9V9bDaz2ra3rQ42qoM6ZneACcZjuVl3px/jlFTsMokn/Tu65iaeNdn9KBU7RWZNIdIdSak
txNEFwD3yJTVogHR1nxF0Ra8X/lqXnXoVJxg0t6XGB3aPY53cNhdzq/3afMKSPx9RoB85PVyV+Vl
S+VDpjNX0tmOhu59n2nij8WrI8LDgeUtkQ8zemDeJQ9gIi7Qdz7ktwWU+YZROQr3Y7iSMat8Qxl7
hGSeJvxLqEZS5fBRjgp3mKjupEz9UQZyhcNL8ndSg7xKfh4WK/29Cp46ppBFjDMOUYWRJPF9tARW
s4+BV1FfgrFdBuXu/9tTYdZ/Opp7p9Hgroj+taGwOVvfqSC1jJ39bU9sJDw+5otrLRerTvGMX6R/
pPgqKrThV5CHejRC5piOTBnJVmdU66hZUp/D75npMeAKByKt0kDmN7hJtMbj2ytm0GMwMFgmr0pf
LCUDUBRqUGYAbY44mt05NF/s68s1OMjHgifltJqfkQHI4RXYlmhQRHO0N6KArBjEsv+IYqwisKdm
zYf3/bUPU8U/Szfn1S9vkOtH6P8zy9ahtRru9lR/9O/hHe1uYSS65RX7WXDohbGrg/0suGrW8rhO
eyvO9C+Nbz55imkk7rdMNur3ggJf9897rzQKo7sxZc5Ccm9Etryin507znPLDUmQt4jz+AcABxYg
AjPZ8glmsbA/aNEMmoT6mTiuwX7lVUtpDtEMGrwii9Ppc8qBinoQWCGA9lKTw156wDbyuTqPyasx
Rj3v8LR6sNUkMV6ZS7LIbKV3OOHgXTlsCD+B33Vg8Ue3ZFn2bnjRVKHi0/5Q087iMOLNjnTjm8Pu
QqQeqX2/KFfx3DrxX532m/OPiuxdPo+eOtUeZXZM6elfFqNtOLkGouIGJJthPayUpgAOFxpxJiSU
B/S6eq2bKiTx6X2XsWv/oJG6DbuotNruJoYKNzec+DnluQilXXbq6f/Z+a3Z24+6iTGF7UZi2Tc7
s2WILaY7Do48W2m9YPoQPSygKCcunLKFH59S3Z1uCHFrALtprIX281vxjhp42LPqrXtkYqveJgol
N0XiV8SH0jL6adAX9Jz5ZM37sJouor7dd3QXD1laADY1IZtG/RdquFFx5E4yIP3ZfUFefamtLiYa
mIMUX3O8no9UQWpkRVl2DvvqxctOSB1vMXZCcQ1PdbZgwz0Dvfx/8iOVqydqlwMVSDS5er2yPrjo
LcRp42BU69oNI/5CgtJlSftvBmVoODR0PhaYdhaN7ULSoGsv05S79A8Eh6yI/1bVc7J60ZNQqWm2
Biw8Xd5FDvK3XUqAv9Q5Qza9WyWBc8eNvyfTKc1/t01Ttaq5C8eYBfHssPFPh4U6kHNaY6BQG45b
zwrbTKruXleyjq+FHMV+yikYZQ9BnO8Vy9nAJ6GfQvNSMJ8fur14kDpN8ZVaxHlJnBHAWX5wu4Qd
SSheFPTdpEXuLwHjY0wTZPKudXvw0NSthH+MiJCkzuC61edLo3UFqGVwI0ecWZQeMjwsGjqafh3m
9p3HvQQdWvZ8gQO05WHvgbV/YWJawPe7wzR+YAfuMk9sr8PaY2uh/EWvv0jPH7CnFRp3hX5ic3Za
qFw4sm81ONhdWZbv8K0DXo78JtzK6a+/PRQxuIL/pJyhDCKs9tNLgBZNzYlzZYXhguZGhVjkFtvb
tQZ5h9j9DpRegRPeKRG9p5I7lybcyOEgVUkUuoZDaN47/xZsLixlqHBo6JvezsrY1EpHEEeXdqAS
4NjiQNUEe0/x2WViPnYHEPeodQ7iaBAkFhIcu3pnpMvUZtEiJj8QFv87+Ef+c5JQFR4NdKcou8aC
e3SLRtSyFryGxy6HeGoWlwLgppoGTAgjrwV0PSna49WqWRkAcSW65kK8t5CW9xspBklaS3THeEwo
IYbUBS+Px1WbqZwyWOulC66eQNuPBnOOl5BGqwn/XdnF+u0ix8OdeQiLTuOJItSsvVJc5R7ybv/k
67PyAdMPPi7zvzjJH5+8c0pHM+6BpuCasY02K4Cc5Kf1VcHwZyLmHXxGoQBjiRHC4rO0YZDp3518
rbjVajndURHq3YAZDZl8vzt1oFmWkDvwP3BGAHz2fSNfNFUGqlMtFKnPt3pSCokPGBgbhNO5JgHs
y54/ShHoE0ovQs4EgGIqorIxHAEOBX37YXRhaOR846jV3SvlFCys0vY06gZwq03BzSiiBDj7g+kG
hrHi+Jt+v3gN7tYNZKy0Kme0DwMNU7UuE1qT/tSZPkHbeeMquK+nGlNDNK239woL++LI1y5krP8V
hA0URHGn40J0PTpuVbKVJxmZEmwHSzc6zknltoa6z4iaq/WBKQ9Upx8EyaleWNsCML5RTZqmljce
nhrnyWJr04wFPoMfJ2UeqXmKenGPibemomn6Eg+2xBANmPusJY44z5TBjTujklYUPVCgbVPS0UOW
sDA9Mm6C+OCYjLBmjCb8Bp8FJJAKtYABElnK63UgMPz/4pg2rYX6BqvNasRqi+ClsQ7mIkA/snp8
aaEic1WIUuOSMjlgonGJzIvc6XeU0pwz2Ob6HktECMrTHRvc1VxphVc+MF2ukM5c8OZNz78rjOUh
RhYLdWczTbSbE40ndrIagZhPiyVZBab29BzanuxfHYs0rhFRaHSo0b4ATv34XvVcpevmMXzrVrIw
O/3pDJ2gHMdwrcyT0cxPmqjMd040MXRUne7zyy9J/PWvgSykYCapd5cRwpJPl8YZhGp1sNyLcF7a
5hH+b8IOb0m2bqWF6lSEhxMH2yqKDOPdz1uC8qxD7UnNrhX16KyeVhoXMxgBqO+KpbVgIuww4T/e
YLDdI9lYwggp9FkIsVsFRzEV2SvHe7t7GwRF0rMTsRaDmsO2lucDGd3m9FJLsT91ZNdeePVqDInz
VysO+7HXwZeVmErBX10IdX/KilWslp+K6lYRGM8mguaDumIcwMJjrcPTeyhrYKSl7D3BJooh5gID
67AVlGuIL+YnBKk3S7Cfo/I4TIfzJnFHE77TXALK7QS7DTkzCccuZGQopBjobPF9MTdrwU7M4/wb
YjbSQQ+HAcy8h2Tq4znoW3ITbXqK3MKX4WIS0aiiBAKfxBfkJ9ZQUAV5sQ/ySYY4ztYJq4yzf/QM
CoKo4k6stURFj6uICFgO3xwLQRWm1SMebTtc5zJPXJBY+BE1K4dO67McyxTIjpKcw/QmzMGgUO1w
Hza8Mlil72I7uccaS6VQfGektBCjheXMsNdUuepnHQDO00x2HI3ZYKL/EcxC4HYlT2dazdrSebSa
hHYxA5i+5xo+RSOcPUdBja5W7FwRvUz/YcVWrJM8XWT+FaD3nIusBMFrt04FgV34H2nul63njrpd
BiabG1IG3ki/Qh/XdARGJ1Cd5GhQLFtH8SM8haf5lk/SKE38aQR2ukXffSzFEv320kQKQzuP4FVI
PWa+IumfRJaVpNzrMCj2G6DiHrt+J0vr1cj98DqZmKl399SwY3nfPW3OgsPzGIeC3kHr5HwIL2Xv
GQOQiQzliKT0qd/HjLNoE3eH3Hh4irvbEhkUOEwOrUXshhzbNFGLe5m26fR26WYZ6GUckEVuKlsw
drgs7eNi1K7FdMISld+Kl39gmxQ7foCCTnmd3Z9Hsyha8RXh90uQmitkN4FrPgliC94oDVWVtl5H
ED5GYD0LvaYs8DqMqrQLNG1oy5d5Dl2vbf+bQXL+ZVaEEPXC5SVCm+F1qwZKgcQqBnR8fEkWxzb+
F8LBqPUR0LkuvYFn+pCR1y9BaGswJhEEe5X8/BxEnID6zNkMUOsaS/yc5gU9zFl6844f0lUMRojR
WAxiUY96smXUy6nLfbSj61sjWWL2lp28xqJdGHWMZkSV3nLc6yBQv1TBX/NlUnA/9KD2Om/W0hlR
sFqfVJDRohe4MEKs/GTylWZQKUPuFdTASJUhKyfNsVg6B04q01kz6WDJBggidqybX8Xq+ozcXCR2
duLqUmUNptYKz+drZ6w/BlLDaknfRBPrYk+qQ3vXDEbA6SyiHDE3ryia/EvsB9tMjpppQLOfkoYP
mXFHYqGlbEvFy2lszECIA9aG413S2L0IgNfkQ6m1knWRj1MvzUB4PMVu1nUABZ9XmZDPaztMyQIO
bTzUZ9WQAmEzOW16Hys/9tZ+hwh3Cy6EjK6SvsXlnTU69nb+yLtdiqQ49ethXbP1Ivh23zhFt4wj
rlqXS7ii0Td3lzX9m2WAkFeR1r80I7fM/C7hlC0uoYJ0xw2a/GgcZh/YG2KvLXPr+jyxM1Ymfo5l
yiTb2nhg90frmb1nuNKP4Jpgs6EMcmHh6yi4F3c9K22uWwQEWcegdOsLMvsuqdftZVGp1n/g85ew
Cpay8RtcRZyGIiIbuzkl/LH1+rmzMRD1tSvKQcoKuORo3+ZIevyLMuj/mGi8GngAtdmmYGPYBEPE
bsIRW2yYXzofAGeO+rIovVSzpCJ7bEh9sn0NM0jZHN5zcsd5wz/WzZcIuTBFfV8LU56hwAigXTCE
4qTVYeFu14k4kPlMs1YZ5IYkW2ZyZ9vxh2xmMnra+zBUrTWLyenMxu5966SCtgIGgfYxG6xldNzy
U4cFciZk0gsLHnviNSmqTNNvAqjx8ZdrRzLY9n5W4OkO+YSsZmsvgZPlrcvZLsNNgqldwFjCbC1n
t48qeqPzkwoRQXTZIIMquWBc6yENto5ipXGeVHf5aCdxZ7oMxeHe7eNY4uuHUKhODFxQ0xqK5rGX
wBf2IVzjQ9PyROV41ThAz1GxJ+hCQu3MBVURmdlSdimTWXB1ETQfn/i343jeLvAdONabezog3i9f
8nIrmAHnH+UJ4ghmpWmUxpINvKI6I9QW13PjCQ//f5kFcIH1xVnMMhNFj/TAdCCfgGhTjUXu82oP
G4fLY7PUlJ06HTl+p1ou87WXTI+H/mrP3fxZPAxHFf5qiBH1cSQB0QZhs2F+ayySWkyaS6Va88ax
BQToI2fikyeyFa+OhLrdjiXwGf8VcxhBfFD98hkV3zcs+dnMJtfEcwlk7M6FKQQqmmYhtTkDGypR
0c76+cc9ZLvRVN3p5AACJuoYXAsfQmeJTmzz1wXoHbWcROvBwpr1daQXW7K/6Ifrs/L7UTrp4nO9
ER84xC9VmqTzrTlyMn05Or4E9SjtyibnMTyZ1J6TWZd2Ge6ZweXnd31WhAGKu9Jiy3/h1IItfW2d
zuSfzuSD5IGRtuX5FZJHWmA68nZUdszhcyJcS4wU/IllmMrW7LEwdslI8tv2r0q+BMSoJiOvPcaU
xlHfItti6USHJZgZ+VtewR8BpsqxNMAiDWiEKsL5WYYZkhH5XPG3TrTOwmKMWBjRo3YEOKuKabhS
JhLAuAcE5O6lXILtywyH1yuN0WEMv3bcgBzJ2EhH5wKcZYZX90+boxGEIA2kDpw0oQfZZ3PwGRNZ
3TyszQAF4mQxV2Hx2Q0OkWnrYoBdyL7sANUrXLymHoAkIiJdN3qif81pzNEqDGYYj+mzFYHSXoGJ
GzfSXF8SoIoUMd/fWEPTSXbq9FbiFVlnrJ5XBBrsw2zzJig0B1KzmKWZc5//0oFg229UdK/fvAme
lSYYBJa58hILqEqrKxUQSRTqpV/MIUCKYKWT0KEymyL9I1iJukbsV6JMp0osEBe3Aqigwp4Z/quV
ykN6e8uiknCHELiPQ4GMvIJMbst19OiULiGRKPAy0TW7LY1RdzhvzvJYUgwBAV+X785S8wmyWxov
OFDNGNuorKt4WReYW1AqIRHH6QremoZXrUaKRKFLnLHSd9tcywrgIplN5RS+4r3tMcouij7GE+0z
Zqm/C6Up3PHzr4oJWcu6+xm+6Z4Z/bZb/V0+DlUzphXRQ2gU6B2S9m/1IETyDjsbYIZch3ORdOKP
K5595YAjhWqA2Z+ThGYC/9W+jFRy3ANgwaTdKZ/EkxrF1eNhlY2X4zMJQTcwTFapEjDdPWtXrtlN
46eNBTuLa4cGJ9IlA2m1s+YAmZR0cWzXgCkH6MlU7Wn2HK/KRTgzXYjRhe1KhCXtN/j463chNODM
vKGHJ7uP9bTyQb8Pl9zXGFboHYuOgFrTTrytp0bI8faxny7a8a87dYw0xOU4q108q9ARWpgmPeS6
PBjTrKacnqOURka5H03AQgkA50BzGSF0EivaqEkuDkNjY0rPbk9PgUXEUVKlH8+esk9gh0UiCFx/
WMxElF9rCZ9mt+MA9dnzYyHAWzC1bjCX978JNeCmdwA9d1QaEbETP8MF4/ZzWCUo8OiJu1YBwx/V
eMExMKRDczh1MUmyHc83AqlgA7bW3Yh0ljnlmjZrxLmyhMKDANH+hmAgVq1YX3Cj/fvJB/YaxOe5
C2b8HoCDBrFz93OnXu6BEnUmHDZzoda2FxPSxuXAn6qCQg4OhYdK7AFOTx/cVyXd+N8a15L97dHA
jGu3NupYSKBkeHupllZNYpV/HG4/tHWooWEeZ3/9cxTKPlgHTrwzYNjgqd+80TVoHlmxpPLhJu4e
4M7AxvtxonHBULH+izHuJL6W6opy9jOoEGNjYbFVHNYGlmPiWDT5cF6z/9Y3Etec3MG3SuO3rPnU
UOrh9xgek2rdmhiD062Osz9nbqZf/i3BVzqzhgtnhaNnskw/rS44DoJzexdGrB4CA0G23Wvcb4Az
PJCIET6WIdyGNUob83e/xSwNKzegVPVZ3i9Lk8F1VhmjUmRxzifO/IuYb8AP2iPlYFSC923QnXXZ
YkMoTYeiVmxXREYJNqEvHV+wuuI63gNUCaj1x72seO0QkXr+RmZkbnrnDBZhjOdgB2C4V5+jSoZw
wgVYFCeoTbuxR3LQuI2wKTH+anTBkOuxigEyZr5El9OLr1v3/fKKwLu6iJMAZQIwMgs1FBqG5kNC
vvbpxEZOEoa5GzXbtcBzIkIKUhbUlmKC7r+pfSH4J+kcnqYOiq7fLwANHt2jIiEcDovF4A8DMQzU
FmwpFbdIRKe8r/rCFSPA/ttN6LIYTboLVXN0+MviBQTjiLdM46pRXycxn1FzlcLxLbbnOBzJ7c0C
38izYa5n6QF9jKATHeJey51s+idZNesrVx2W5Jdx/omrSKCsOMgw/r9uhwr0laYQFE9dkfsd1wTS
KlLouayDiH63C+oRiZAHKVRzGZ9vCl08fAfzepccOaa47xzexuMQ/4SRnG+CUY5fTaFXLtAkKiVl
0OR3QtckeKfAh2uztC1rzSgXl1gcoLh+uzv8o9KN6gDMMg8uL01jGrMtXuTotjJIjzBXHkOaMXVF
KNQ6tk0WGpe4C5Ice+2w+CDDbzRVC6Rwkf+DYN2/XehH4tSP2WPvY/04XkPaEOjwAY7cbmR/nbam
F9bmZJWNXRHvHZ1JyAfyDQxZ+eg+pPvcuEOaST74yEOTD6B2hVgw/cZz7s2duEazAOwyDRDGAmop
Y2/qb8mVDF5JQz65P8qk7Oev2JCuHRp1vtSYzOazTsskPkJ6wLu213M0y9d+Cxxcc9tzw5jET5gC
vrvqagktzwWLB3eS4bEYOlLy1J+8zRvZf//ud8sx/lQOm71iZXYBbLh8X7OyStEOcC+QygbDsN3C
1hgrn4hS/ugCgLvRGqpwwZIq+yjMRHKuKri2fFqef/UJ4uaWIe6fNtrLh5B+5WzERWafGQmIE+Zo
uTleSNEXleedNeTwLM+k3Vn7JvH3c5c8oJk3GI1zhKq5uMRdso/ex8eYV+potBaCRXk4lzLrvXp6
N32cXeNO9sA7KffA/YW2N3StVjwWMNPAAnpnVl06FtIsd7sajgzn4dSU7IEAyYf0Q8Cn06HBby2Q
xua5jT6PaFZLM9gBkbo7BQyNRlNG6EowsMSlSYyxYmRKTFLJ5RQeQPUU2nNmroEYv6Won7Wx10gm
cFflYQj4htrwISfNGRa4Bg0hjvSZORjGiq7N9SBjKx7kWM45D1I/U7EK+ZFrLRmx8ylUpIx813Tp
b+/E7fDX3funrB+8E1xucS5372Qaf1WI7oYa5tsw9rX/d5ztUOmuGL3aXc8Js/HK0McFquIbm6B4
rlsb5IZ+hIdecRaOZMWwjadYhNS+M4hWg/9cDrSkMfHPCh9kL637XJTOVi5WT1XNjefDkB0K0dsJ
omhjD6NasGaf9D6qvuDqTniogfpS5iW2Upqrp8ToWkXVdxFoI0bGDZZwRp10P3vqifmGsWjXCrsh
nnXEEAHYCc2OyIW+JVIMu3+KFJ+7v0KLgb0IN//wztixUC67v39/a2Ag8O0jiWOGRiLj7yvb9/O2
HSvAPE/vjexyfMTbhofKoHsygV0wnHXYq363w2tfai0Jv7RglUnaiqLGoVHVSlRSspyVAf6qsPi4
USZSWWHGStDudQ73mj6MHQ59vKiMysRm3VwQCHyiF4Z4nhod/V+83UoNKdlcEmDmpDP6zQavIRTK
bBoxl1E0Jq+/Jll97gO0yhaguItWAJRlQDJgiCyGAQt4SxpQLu7oaLe/PjX05Ps6Ym97ffivF/uH
SV55Opcp/538e4UtiXxkIWGU0j8vVM9Mx7WUIrv6IQ59JrQ1QblVmV0Sa7t0zD8Em/9yngXjQGwI
HZZiT86VVIl7UDIAhcTAAYRhrlFHGm6Y465hcPjYxzxe0SK2J1S1jCS3YGQ9jerJsYfFrlm3f0se
dLnZ6DIP95HROeojU/JBe4oi5dkB58+MlfBfw1JYdoy396aV7r6gEINSZPAWqRX/ixIIBN4svZnb
aDJOBUP8EPAZ6KyAKIBRV5kxBWbYHyPCsiPxJtL7sFnrEYFfC2MeCjJpOk4nPAbY0KDZadWZBXj7
cVo4HzGK/PdltXKR7QAQfz9aQ2fkuEu3uDvG2zJhU3TjtL3LdivkHMqZkhQmbAa+I0jVp/mNSWfx
nEbwj4/6kkUhrnSIsVVqwMZ+M3VA8ILT4vRVwOrLk1GnCz6Jr0yZRmiWhFNzztglzD2xo1+z7Uzg
H/qXl+umCh9QJLsaVfKO+D8L2VtyEfjD9reUSm5MLEd7hzaFvTjSZz7NOPJYKgDYPIvDfw0kmsdt
Yk9oUZGZS29ANiPSOjnymGHtXAcjXi3+8Z0BB5TBjIQTrnY+bObuy7S1sqWbRG4nTl1sTUlcSV+9
tnI9XCEzjrP/z12oJ9hq7bmoRHuczhWPLU9H0jizvmrc9D2hsuR3IGrUjRRliXXosY/PWPBo4Wpw
p/XwPAK3m8Tx0sSYCuSmKninuzMrFdOdvBCjZvHgv+/LR+rKjHNc29wiWX8UNgOQww7TGeooCo2i
RxwXx877digoodyyMNcV6rcMCqmEWnLAYNLe3GVq+yV2uqLn5A/w4RviQ4FjX9xRX9yAFNqbksGP
o10dz+oigLNAtpKggVS/vHRQYEZj22hCP+V/F250AQ048NWTRJto5YVIWWTggBHERWBXn0CjIJcV
+14c5wlPjTzPsMyxl0McU78k/TdG9Kr708pc/wR/XIpK2To6zYNJ5xEQaOytaNf613thMHHsl/jW
ONIicdQlU0FhU5ArkCDNpLmaCvNaYD1YYer8fefkTinr2wF9qSiGoSds8E4GQ3zBKi5qCIiXla9G
0qFvS3GRGXdktgymNWAvwf/UGCZQGg2busgQRxRsmKghQdqfueEx65JmygzHxG+s/lmayVUWPbUj
AuHKqw4yBWkoZ40m++ro2QJDO0EqR+tYKOwiLT0IUM/3TuSq6NFImAChCRB2ejDVSBBsWkH6hd86
h+GLuAOaV0P+IFYEpicu4gHjTEtJ7ADGgP+OG2pqRzU16FHsMcC6QrfdQ8kbXXIZQYqu/cQxXiCk
ePwtK8GxLgp/DN9bNO8gSND3k97vE3Ua8tWdHC6Rj4eg6gpd4RsbcztRp4ZZPr25lOXyAQQ1uOt9
6HHjzjMqaYmanRSV35Nr5kMyeRzXt4gdlIJpUDqdD6FUOrttPkssZTrqZ4etN4WHg93DmF//JzpY
7GKLXgzFrhkT3isnpWh75oP1RXjgg+uENUwbtXqO0s6hPho8eOsGqnBbW9t+6LJjgF7KyrlCJxWD
69c7xvE9+VZmDaLKK90Yg72mFnYtOufp+ZJHk9j2d3Vs2G/rPInExCpWOEWKqOiZVweszh+n10Ky
fq5DDaYKLHPfdUkQ0dEBMGWzhngQ5mV1PeNymI4WcCQmcWIGcxlrrK57jZFwBhJWYi5nTEAcCv/t
Uyp366K9XENe68YS38o6vbv8QsFrWWM96KCUSilJ5O575OIcb4b5NhCcUKHMvp/tdAZoyIyOf5ei
3r7DzTPnHmU7z0/THcrYbioofpnccjyAgpfIYn3vDQtmm0TT+pGj5lEPfGxiYAQrJUS801RAVqHS
XwkbmwVoUozFItmH9YhoK7QlO/xmBMFMtIy9oHYG6fgAZOIqEBND3FQ/JawWcCRsqXrj4Pl+RPid
aJFxHGVp2JxJBSMnRqY2h0cNUKZQzM1iDGciEnB5r/nqEIsEq7L21BYXaHHcmMtzZEkj3grOwfeL
jsxHNbJc6iix5MFMIo+lFx2CU6wsT8qRqsyvpa0WDttTt/Whf/yDfdzR/keWKml8JDAMwCYDXvfy
GDrjxk58QnV12xKfD2DfEUtMTdcnOG+BR+74lme6yU9i1mg1YOojCMumtAU6gYtPv5y6tK+CpTkh
3yGKe8XplxiXCoOPHs15kJUHVZiU97CHqcY1eup78iZE9h0FI39ZtpMv48ZlAcD+YTLkxJx2H6x1
/bXaHZy4kbZmpeZdH8maqXoLZaYB3OEP5nIjbouLIJySO4oe679607x8KxdJ4ImoZ0LpI0YsB7GC
2+AeazQHBFi8bVh6ShT3Uaco+sNnGQD66aPPIH8mYT1402hLjD8E9s/zTjJ1XNxhE2J61KzAf5et
iumUxPjupuQpaGy5psrojvHPm2/p7calODLQUZheOk6dkDf0c70jM8OT6saBCoWClP0GaMLhrOD+
HGgPFM04lgbAz1yAzMK01/HPZ0vDPUy95a6rK5+BgDcjlAqbbtf9vPIZQXgWypF2LzPpFj6jbtQz
24m7aNjA7kgt1iM46ZBguvq6GBOJTLrPtcmyDWQp/C+C+B++Fb/UI0dEwHH3jbvQWMXZWnoQ6B4u
oAQxvHDGZI1gpjsJ+rq4qd6p8FX7mp/Wm2/3Srj3p6BE44+OJmJDcKEwkZlV13yJVV5nHuouZpLh
EpHWIYpj34qlxc4zh1LPiMgP64yDmY9KXEca1eH7+D65XqOmzcVJpj3hXATbzmmUMofaRPrvEsWe
Durb+sVJPu3Oy+FfH2pyxqA9MJdPGvpEQFGb81I9/EJCNd9GjlPcCZO+K+3HkzpaH4/fn1g+VQLH
m9gThUzyBs6xAKn2kTxzjUt/urwvfK5mhJsKUdL+gUkD5V3yrtTSQJNPrpnrSx2hv3BSkSP6K07S
bi4w3xLLid/tX08011STnYG4kO+rzfbuFZgGZHJeARRb3aUfMWjNpS0S+9AqMIvwQETHsdRL19iP
LjydDSdCsygGfexDRlPzngjgyGbeXatClliHh7fGHqbfs3BN2Gc1XL5aMqBdTPUJ7QqcEMopYbL8
zvM2mgDBOJ4fdePStInPfXqbboE4aJkgMcLv+Vm2OCUBZwE1Iae7yHbt3j+GfJchxbcinxp8Cgrz
Xo/R6GCC+0tpY4ZljjO3nWd7Xi0obn5w9pVjJxM0BHia1+y6tqDH4BX4xSrDzsG5rGq7vGctG5Ia
IjvEIwUroUc8Zzahy5cEie9PE7AO4Hp+pXuSHodtYKvgsY8scPRbRgKQ4zNVhl52AmgfWVb+dUd3
mkQqGvHFANwJSUph81q+5nh2a+MsuZoMIB/T++iSPNTcA3XY5Wc6C2T3pzTwdFFidrJLOghvUkKq
pri/SBkf8VtMIftyYey/3L6orwbeC8wvIPCUEhvSo40UFgOyxwBJTrmVvE/Z9jJH/2gyZvs5B7Mv
6hr8pM/RFTSJp40DDTJUUkSGgEKo0Hyu+AObSJswBcsPGsT8Jxrq2rxup04oKpU4Yvu7rU4iowK5
pPXW/PtxGc1B6r/YZtIVG5OjJPY+a3AWenjKNrSyArgaL+mz4K+d0LLUb7cOq0AooWyuOQQGOvIL
ScOm2aoOtBTUAZdVbP4E8GQ7COmL61VwdXjOoR0Qoi/UsEhuAV8SBvLUIOZeYYFHRcfqYyQXZPnE
r+7DqRIqQVQ8apUuHcJC+32cUbAjQbIJ+1tUYGyCCNCtS4qR2rlKbVfA7F3Lu/HUj7VySFs7Xbhj
9aa1tmXET4aQcNggvx/AMP6NZoROEMNFo6OMBtGMCH2sGr7mJShtLiBJBFzt7tY44umiWApeynZV
P+1KJPIIJi5AUQY7tgSL+sB+sYzmunf9tOL/+VOT1GOGvxbtd68ieXhC5kd8v3AnINt4j5V5bV4x
vw1HWTYOpISO1UTUYG6GbaJ/3trBNa4mgPMQGXlqFu3Iozhh8Xgi7/r98wkHqBqAhe10MRvPYIzL
qaaKLab9biGxYDzBNtWy1uvIpmuqrkA9hffSu+PqXFaScv2Mnkz1SAihkuP1zZ16F1gARfVMToUv
4gccAojm0N7G7JBVSABvY/JH6bh8zwlEkCmf+Op77WDWvZWULEsaLbE8JIF/sT8SU/mQ0SeqiEaC
WPaNSvV5TfIGzXK2aErNsOHMOAbIsuC3gRVKbkFafe12bJbE7d+GAq9QViJwx39Q3FUeZqRQAdt4
koxyzQqmEjZS69ex1cV+s/901oh2Q7Zwb+XavYkU/xJHRWqpxr+PzdyVqEjguzaQottXXLS3D/S2
kR7KOhqcJXxfh6XuumjilXSxEUpeWVJ8TMw8jnnJPunwPceZBEUw/nAFkIC63E2Idk/4r+8GeB0F
uJtOBJh88R51IGbt1fKE+7jPpAfhYbkNBYRray8uLoXi7S8ZCfxTUbA+m6TTjY6FR0f2MCo5YAu6
oZ1KYC99nJiLed50/R7R9NqJQAp1EaGl0H8lQ0p1is4DwYwta2W1VijqgztnkjzbL8TBfqoRQUNl
M8NxGjTVo14YbEe6iQ6jSxoQrqi/pnzsfmK5JWpcj94qpopvbhxbYDY/4zkLFT8FZJxhXH/PC0Rd
oEw6egHOFVb6WWaZY564V1coaKTobippk9CCRkudRfDdDY3wpBciE2bivQFPBc39DuZOWv7j5rZ9
xVBkYLs51c1jg8S0GL0ci9I1sGlo11ZONqEa5qTQQ5mnUdSl37L/F3mkfDM4yp/0aXdHiohRCNTN
tNHMQaXD7salkmVnYDlxPPlaVkoAN9VQOxxDkdpv/cvQTtB1Ao+KUcWEVy9aWoJ14Z0IBCs9xV70
YI277PIqH82UIK27R34V1G3fFiy9XNEOZA4niYJ0587MhmlzK84b98f6I6E5IWa4ooIsAiFJipK1
iQ6zP8deXCEYcWJpgdp45u3wQVbVXbfMWVJrmnh+OGKFWLL5kCk+1zs8DWmLca89YhlJsO0M9gZ/
XaXAY03t1BYO6Tee3xNKNG/adyRTzf26UP1fHWeNWHKGa+XOYtWj/fU6FE2tAxyAkNp7oLOyh6iK
rkbts8v8z/kuyFkvD7flzhsxpDdHYtV+OusSMkoTjjxOClTs0HZN0ZQc4cLzJ82ygIO7JZUA6ylx
m4QelpBjlGThaNClHn4oWlHI62mxEG26vNjmpU4RMiqQLRaLLGW+XaFeni7DRwqvE4XCwiFq8Esf
s61reOcpL+Q17MFWW4Fv7ZSiQswZJonLlvkQKEkmgYg0zzJSX8D1Rn0RtteCibVD2MkevfiCMvS6
7AEjb03JcFKzrvcDeWP+hXFZjGYC6R7mdKghfdG3KbRCO0zAKmM3LwPsziF2dVy3NEvZbTgEiLwu
XnYMDVp0qci4MOmLyw9ZKub1vYBVLzj4/5WoD/LTRvcFQW7LtM7zCv8/lDzN4u4xdgFV9CQnmMKs
W8GxcSQwmqw8qVFqrzt/dya5QbIP8eejHqWBEpbrwZ1QauLmYPOCJfSPg4ApdjE60GokH5HCWvlN
8udz46JeH6QpKizlHENM/dNKhwzMXOdIzXd2uHVFDywJ9oHGK6Z0CRzJ9Oiz5DpnlK5p+QXjTOa/
g+U3OfE/ZjRYqTjCHj/JsTtFgufH9MUGTojJDsL2/i8wPAkLsSb3sA8JQ3jI05ykAzlFtRIzg2nq
K+z2DrHRgYaqrcYRge9om7fhher4g5mxgFXRmwcpXZwDwpz8T/VaaLPWmWi0pRVMyx2N//BZHHMr
lN7Dj9lC00W2YWH/e9r7iK1DsWSy4a0UtO91j4dQ+6nkE+axdQFNe9sYlpgf8q81Ij0ynTjNHk7r
W/6IvDSunCgTEMNLbPcpcHm8e52Sq/HeyXaChBZcp6oqkhvpcDvByT/ldtb7vrupqi9G7wd57Uc1
Hg7KEjz8KfscrZeat8qhS6kge69wO8RijmXjHHg4zaXhz/RgQO6UD8ulJ6xZxyZr6lcfFFnZIE/w
4Q07hIo949DojAOR0HIogUrRxcPK2OAByUdjaa3+IQVD+RZmJL8WuLppuJIbdYNJXeR7B9rX9t6L
8xD57qsNEhpKV8/aKoA2EdECMdHBdMWpa0m/LAVkkJjxEuWvGxrNPMgDpgD2xUH9o7ozNgeonFEE
Illl6HOWJfaVmSVTw1oHAn/3s6CTF14Ei1d8ruX9PkONNODfVON1Wxkn9m46N/FJGI2LE5+J4Vbx
BFSK3MLYb4SiV+wkbglWrxb/WIWiImGh23tosm6YmyeamzJ48MRG9yJG4t8AhGb+dExF/Y0WkiXg
v/0XJAMGXwVWqCRaweXYy90fcprNJkiPi+5795URlLt9l8mbQmyF/VIup69T1ykgBh7K7HttT77s
FmK2DxHz0ydVcbhdOfjczMv/KXVmuZrGbov6OLL0X8lGkwP6d4+C6QxfpMZdius37FD0oYjfijhF
dKMjYKX5dUXtvKBBN+WtSrqCxcnxNYQVtv0KMrCDVru8hKnh3VJBjgGIVNEyFIuiLVGlS1p68kUl
gVqRXhd5+uYTYs5U1vizsxnoF1gRjeoggXHNs+kiYKXrU4+JWyyHwONHdTNjnhNGXxDgSKXgDOG9
AA2hXlN+AaMNKKs0YK2SeZrM5ylgAE7XGXPziiUzSK+zF82zQmbaon8EHEOVGA5jr+fz649DPxrE
iPiT/2wLF1dhSOYwkdzlm2KJSugUmujbllDVrhhX6OUsXfhYV7ph01bjGnxxPrrsyzPY5+yaQ1AY
cq5P0fSNdpJlvESVsF0K0uzR8cu8WGZvRYrb7WcZEc/9FrIp59/LyQRcT21Y7Ax5tNsWa6r+2pfz
C6rUdNtXZqy+u3SEpuj5Os5CtiYDUKnVKhPYaV6rTenS3lcxis0Hwfc84G3m20BAq60SwaHHhPdQ
J6YvDQwPjXPPtU+50ruwP/W1rKjkpSeGsolDpobcX3l/N18D+dFjwQU+YDrddTLfYJuncY51ePDK
RR948HBh5IsBwpXKZ5kC9zA70xzUO2XqDA1wX9HBtm2BrjK8U+wxBnvw+43sKKnOVyDRfzrE/+ji
LBCm7TbRZua3ZDrGNtH29QwXoIS6k6O774dJ8SEiNg4wvhQ1KpJuWXaU4Dg7pdunaf8U3Yv6UmaA
cidabCSvuwPzKyR7KS8OqrXoUIcDbk7kzM2Zk5tvzl0E5H3VMBmEwH0fWYs9SA3q2BYYc+c9KE5l
URziy7cX/uHrfQuMfi1SbTH+Owwic/yyPy66az4DGJxxg8sFWGmNDrkyO8bAfyxbFkhrcZovSpAT
syLiJV3dFICpOkRHLd+D1DiAo0+aNYJrNtpbkjY60bWGQvVyqZ8gQ+/xSXTNd5oSXZlEtaNl36ty
RRXjbN+5mJ3sHGr0MSoKBNLPL6NTHEPewuDewKSryVWOF4I1JQFHOv+yciEvX9AfWh0Lx5lz9KUQ
S0nm4LzISbvEEj3axQPGMgsOQlriD4pGVbTp4rDxzQdrzKzABk3LnKlfR3emRTv6SSe0NOJsqqwB
jhdoBA+vV+Kbl18Y7oNuC7JimMBPnnxA9W9ARgQOOmoyiFHrCV1BAvfYDU/wRfUk+1zT1moJoed9
zF+RF1RRZUTB2x2ei8Om0/d+9R7Ycksg7RlkokFr7BcKi9ttsSmAhHmD+8f/SPBY/7RClFRsVRKI
xbEW23NHaDMCtwICcI2X1cZHbHIML+RbpbxkZB9SBRjRj1Gdnsa4EEOgkD8kCWFSfX+aQbrnr63a
EsWcdjefbiDyr3Ncn7vLzhW6IuAN8utGL+oabB6d1UAotx9F3Nct0JMheeQRZNGPZuLbnflR3Gm0
cxpgYpVyuYsV1hgG3FGwMrFzcdNpahck03Pn50RdyHTGwmP8CRgAVgHsfM0M7pnKgJKwBwkEPsNY
+sgv5bLR3qLIYJZD3GcBmu4AiBOJDfVRqJPWRduucWhQhqFVa46t2b/y1vW659X7adZPWY4XKRiy
hXqsVTIgJfe7aa16wmHxfPHt515kMure4OEA1KJBWpXUHOV7mCiSuo5p2QtLDa+UDwvD1sF6A9pX
9WQcfdK7hKlwzExwqfyuBuueYxJjjT1DHqISsFCBdtYJYiDH86suJ2R8nWnhv/9RhNBvL3jBXf0O
N1oY34iG0bblCtBHs2pPDqcpeuTbAqogbBI7agDR0Pa9Yva656adYTrFG2ZiXXovMHZ93OCpomzh
LLDZ3JhcFhMawRvS5JpsZkk+vrjAoKy2tO2EgdHawPKrfSq7Euxv8OB+GX71K6yCy24j2O3n8DJo
sbwFbMMQONGQuK3YbEyJBx3sb06CJl9hMcP19uCHd0KlSCWyzCZVDyotlxIvW+LUSzqmsz9M6tQr
cpRnID0omzh9Islm0CGvFKrC278xxziXn6qJL4tYIjK68ws0eGevt8dn/cUs4zxbncGS2o9Odu8y
BOIepfAqmM5iImm2bD9QVZsHRp/JBc1K6768fww5gizTNgiGKPNvrTVkdGHYMKQ1kgGE6nKpYlaI
S4n++oklA2Mwxx/g2/xOAS7WEXiIDJEC4V2PPBp2Fs/kATCMPw4H2j+wDqhO9TrpV31FJgIB25b+
R8CiuQ5cN1LqddIzovIRfWuDRRS5uHBlM2j+xA0orOzrRBFbmOAMhilegTIN86Chegq0Ffo3xfA0
mT/aCtC5guoqcR0kT9MosZ8Jl4Rz7lRvGJ7VQWsLZnJa3RwSGzR5RmZKvgyskEE1dpb9Al6PYMCR
SEaShSvbzuv8x12VLWiO/HsNVCEzhez0RJkID4mt2sKW/NHKHogTd3rV4DXnVzewPn8uvfPlZDMJ
G0jCNAJj2iJsp93ClH/inKtG+oEghp54chdoOEQenBqQQu8kH8Xw5vD6tcez2NlKmIpn2pRMF/gt
58Gr5eDCAOKp1x1KLUNhFNpjRdDYjCL7owC7yYmn5SQ2Lc+Pjglw85jQN/qXgJNeAjeiCOmHH/Ci
2nPM6FuJM5jGhc/MPxwEcysTs45IyTou3uqqzmCJAfrBUh8dlKNjy5QVwKAGnpi2A+Mf7Pm2NqH/
k5j0yHsdcn0tmENebawNxyFGxULhGLulHxkFqD+BCp+N12Kh/+huge2eZAfSsXbh+Sdjsib731rm
zIzG0JwyGDfumPalkaZFQLWaviUwqdO7+/GJzSmOzPxsqDaEeXlR1doH3QlSMO9wv0AKILj2Mqye
sQnSWl6mg+gf22gEwAtsEQpoKEpVeykMmYWLu/eBx1k9je7M76mBHPcQMC6jRJuDED0jBK+8Niul
B6fkOp+nTfBNI9zqkyCzfxgJXJ3XvbVQCGjbosSKvk2Wy9ObqUYmM1eshUYirQVuzvvRfJbkCxTj
w9kER1yGIg4Hl0VlTckSu1kb29dq/L5kMm0c+ExyEV6m0fxXaarCTnNiV+SIDOgHPXnLCYkPCTgj
Q1FtSF06q7us2axFoAJveLwoSV09g2IVEbIUs3hOIkgySQCBEsiT9VJsky5osr06PBhOjsZG769Y
12+U7dSj074R62C48a8JlRHkb6Mj0Z+9o099bgrSTD9BpdIttNp2jjOoOwMyGH+rWqeJJcxMeP+I
J0GdYsDmp4mawG3GYL/bfFK6VYj21US6w0ggAMnYM0PeLPhJCIz6cIZpUcUdrjmVAbijamdx3vU6
siUOS0ey2yL3Ft9p2fmPX1PPnwc2HBfmztVe13cM8DnyUOL8SPmmoonNT14lhne9iYEV7ECoe0W9
RzaDU+bfxqwHNHfQGO7FUK3TDqb/OAS1kVtDzimcNPyIYvltBXdBk+INaia79fT52E7LwWJEEg4X
y8i3BZBS+1S44+ltFhonQyNaGJ/pS1mBXOYpxVw4ARlyGq+pK70KRB6k3MsnAnmAsHqbY1ZKthos
SFgDVAPlJNk1o6bBF7ny3ta9BNvE/TGTXlXuxqQeNbqYeBZmzuqe2p6IRlm/0qBs3mFRokd4IcZ6
9cm3Mr74sL7VCgebwfT/YzRJbjM3rCJeE6jnDmxSU7oJcOsvbrV3o9CQ8VQU05CFpPoQN6zQpftr
rOfs2uUBRf0+6KGpmwLZ8gCH2sJfLj7FUuEMex7TYK1V036pyqIY3G8VWseGZoZWh5jeZZ5Uxhg3
TqfoHtdUHHViSgw8Xof8gt04nOceMDnOTPkSVGrk1TZ3hoTzndJM/FUp3SecfW8w3tqSC0lA2bPx
8a+s7VnzB8awtBHYNTlByYK3l+dVacJckpl0cCczQQUnvuE54mcZkawQVltS94Rmb/S+TNBd2Lew
WTKc288S5RUuuoCd1tr79gQIpExH6ZIZnW8fr5xv/Rmkd4/VDoGW8aVagNDnoRF/JcxPCZF7Nyxq
Bo0TFgVTNh7Uua7qvlQrSDgd+fZR2Vp3KQl5vl9nyl28pTbK5k7Kjk7hYZZsij2QW14YRiSx3LdZ
2rBok74XBBZj9yoOZ1d7VGePqt3E/KKxJAIYJ/fc+x9+ot0qc2Svy/HMNoPtNuOUMeApIK7zquoG
7i+41lk4Wd29rSbF+7FGqXNqEEdkUN/hnEljfJhxaBCXA4P7BJjinbOgkpiBlUSQ2Or9MMITkjSV
D2Fl1jCdXHhxwsJ4qBebwHUDRi45p3Sv31Jav4JChgOPk3mpLpAp6zpIXPJJnpDDTITElWD19cNj
qsbyYwHJ4edRLKyAtbdA9i8d4mqb5ZfzLxjDHKHX+nrJdIZJdUrRT9OplWr6ZzWzoBo31ydyXuSn
5o7opxPxGaIc4RqGLpjsHK9Q/Iw4qBa/2NvflVpGfoF5+MuS3wzcezLslVlRse7+pdF8xZutph79
1zjxsXxGTq7HD/KsvCD2hYN3nGsiZvbu4gmZyuYWyyXn7eUJ6vqadyt4N7j6pVge0VrNFDOf9aRb
oBgZoB7OcOA1cx5FW5cvZC3hpg+mzRWsAlYfkcdCdgQQO4TxYKP/92SIjUTNis8bMUsz7jSGkOww
VUspxYB3LXri3PvgPG6gBxZb7rYMJk+F5WHsaVQCms0LH7cRjgRfAIi/F6SDuYAsj7EigacygGxL
Ijy7RD7J7hYd9ki16MTvrTOORDUUL5JVfRtCAzpIKUeoUwWNfVtgobGVuqOOdClOQHQbB6HTd9m6
2g2xn5zICGlLALsvO4kLbFvO9xi2mEo3+IEsrtADs/ciVvAh/qBu8NJ1lf8wHxHb0hra/78Zs/63
d1XLXhbsi7goLdcuR0cxMyG/sIdmAb8wbL/IRbBiyfc0ezMe1RvYox1921To+Ps4NMHvAJZJQ4Up
aUtWqVayEq8Em3HDNhZhd1X+pqY0BRn0QNoIeYknu4zfQnSHVrSmuGUuNG9Do/p56xwsW2nCzLzy
lczSLs4MRqnk+RFJ6thFymkYmDsiDxbo8nQeJj/9kQQE/0TPvQGdVn75CLEGE9ODpYf1YpZggST6
Ne686e6Zv3IJh+zXBz2cH6Fip6gmYs64E+9hpnBSh1Z5GHIciI5vKctTzCIrdK/4sM2qzcuNGnX4
L1UzL/hERkguv7gDfJpG24VfAMBNtHGhdGT8fuPRrjriPIXIcek0d8TXth2KI8KsYftUZHripJbZ
cgEAjGDcO8sXtjVKjn1UQ6JXCqljkFRMRSri+fs7dWoUxCeE8/amZlM0D+K5Yg4aU+daHT/zBEpG
fAWfLmqzHSBkx746tGmw6rxqYNyftSbPVDB4NyFL8rddH32EsJEYUc8bO1y/7Jp7I4vDoQBdSxLJ
O61Ny1NncsFh4Bef3QpDUvXBjSIyxzoLnkVgmI8CcMKRVZYQxdquNops4ewfTfrYCGhFu/1gowbK
mVjRoTdsggMonAbQKWhSc5hATG7no3usbqqcucmv5/prLlCVAgWhTMlaMnrIg/hpLSz2b98p6ElS
mvNgP8w41yeqN8Y+NUwQHoQ01PTzV2ARvEphO2mmUfpIUBrCct9be3WLtJCYxUnWr1wNux+v7mlh
jr2y49ySFg5zdn+G9Lc+f4aG8dUiq5SHSQqbOfyfBvPiKt0l0MSgPlkaTMRJfXRmQSz6iS4AXRwl
156HyAuu+Sgyd+UaESgoK2pKf39Ncophxs3yZP9OARWUM37MLyu3EcPgvAmTnW5fSkje3T+uenTj
vUO9BtcH2fTDDTNm8BnP+J1QIRYxQ1U9DSYbPBQ9dgGTW5yeCCOqUz9Jh/QoCo0ZtKNsugGK6MQf
tqLFxOaqwAJt4KhnZIE1hnNPlmsENQr1GGLOGvBlwjSeYnw4SF3vSjW+zsJUeFPRxczFlVvVCHyr
dSlJ8SSJvNrFGXdkcHpn2HZ3DWAW1QvUjtoB/0LFTZC/qHFfs3DVUKJizCYNdKQAz3vHtAJJFoNf
Nbkro+tgu961pPe71FwKcI3fGPKK1nYr4nrGkUUnCz3+DVM0uoPfqx1svUhFcUa/U9HR9/pWD9Jp
eHotEQHN7VfDj+SpTYD/fmoQAIC1eBF51CPrYm+rCLB/nXBGpSQ1/es5nwT0raDgCyy6WjDwBOmL
/yWYGKRwq+KyaPiXbLsk/GOfN7SwnNp4ZZgTlGqtKCcAMHHu2/C5zkJxOo2gN8io50dBd3QpEVD0
9Sz42babWmyKVKpUjKTu9pd0t8dn1cGE80st3KYAUkgyhuV4J4joJenTDwVA1I8/WvdW/ws3m3Wr
8CgbssgOWYsZxlXv07ztYC9b+/BwX9p4NL/zXpebTPRlwd+UBGqZ3ug6xm7Ij2Uh+UJFw1D8WMKX
ZNSlqXg4pl22ENseVprfgLutc7YnOBy0CHsrKwHECnVMVDGOVqElDAu3R2XtbyoAjUgk3UQoO3kO
rpasS1jQVMHw4EVI0Eu54gNkReLT9qFu1Mvq0o23DvngIHex/MMG+kGzNqEiAK606K6Cf6JH+XPf
hSGG/+O0DIqj4RyUernzXfqZVPbz/k6p/jl5/VlvUFmdB+pvjuFGrzMstDGSSrbo8yLppNIteWUM
T2zR3I0vfIocbrzQtRZJRUmePswu7dWuyZUaEXi2Pt2ehLI3TdfREcVDghVzD0WHkm4D6wRQv/H7
gNlFECv8zvyZe7ijyDYU1JFIsZ6+i67DXTde99lVS4yO5pzNeH8rtUdRyP7mgiMbgm/JSp7h8uc7
hiGmFcVvx5/Yrm9j0qb33G5sd7fZRWLWjHc0txjXM4YEM9h7PX5jBFrq5z8q4T8yuSh6rnqlsKBJ
5BzuIzJLGDdj6S18CmI7DDPH0cDrsFmBPDajuwC5s2v2ZNPWdpSBHxWWmsGy/0+OeF3mkc2zByoo
ycDTxU4Y508ZtrNdYQVPPfd2iufKl2bODioGWeW4j64D9Oepidi0VcIZ7TRuR/rRGl81sfKKqMwX
zChCrckWraIwNnh/UsG4c/agcvn8zi70Ypr1ddGehwyslxS56gacwOrysnpWwfw8YzssWXlRgoce
3aP9BORYrDFGbN6ONIN7pVSLfDf5TGTSjkppMmuBibJdvWk+Iei1vViJg6K7WZzdOdPj6vlAvpho
mwahQwIiwS+BPsmO13mTDeLf7E4PLTBpoqTpVIQwiiymSj3aYDVZmbreE4w4mywemvB/m1M/L1e3
imEPgqu6mHoQ9aYTmtfQu5WG4l0iah6UhwBLzqaFBrP2Lay4s9gZJG8Q9kQD3PbZ+tkIx+0cDrH1
e7MmC1BmmWhratErYuP7aDUiP3btiNU0HZeup44J8Y9FyXQngSj1i5AZVLim4O6JrVjyS/xsKqnv
5lRcW9imTyxRVdEI+80kd6nutqO2wQLmNAg+5ccbwtkj6rT8CVN6T0XhbmNSnDc1YrEu64O5PwCm
uwNnfFZB8UpUnQc7RVm2JzBl2SRjTs7nmllcQ7c+m0GTRxyntKrW499JlsMm9V40W+DPFOGqRwUZ
/NlcmMtZ10H+iT/NiXgenh5e25sSYOO0LRrn0wUrQLv5nTEjbCuG7NnKt+IzaRr/PLkUsMiyf31W
IA2xd3Gj6wvKvfV5cnd+8l0RD/I7Rxpry2PE2sg31CEIeVDZOVKbno5pWH9b010nUhRbUOZJA5IF
uYOCpJ4F5DYRJ6nV+nhIDZe4dmTyAtejKX69l48YcobZ4o7d6jz1J60h6/RDgLLPRCC0yNtlNOiH
vM4DsSTtELI/EjeQaE9u6m8VZchr3lc1trgkdTRpsdexRnuSKE3W8VxCBDMPbt/PVk/gT+s15Cif
3wp35lue/79Py/XC4ejOF3lqcOpD6htfG73rTLyDBzbkOzWpAFtAPwLryZC+TxCXdfyVlk2oMqcN
7MxO61gm/In+MNhtH08Gr8vwJSDuaOM4X585kHzWW/+bPaNORHQmpi3H4Ah1vSDgHPsRjx5p8Hgs
LgvWCqE2Kut94SvaZGpBK6hQ4rCggqu7mOGyl+7kr+KlgQwOfsL1Rb6Fj1Va9c54FVmZiSrIe63V
ObniXNuqU74xmSmWlpg+RFtPDOgT80o1CcdNQOKCr/OpOrIO/T+UhZOxWhMua22KhL+Lahyfzd4A
u6uqWsnlG1hfTno5w7jvT/oZ67pj0r2P1q0hXa7OsriHKpzV7QKazXAqNniIPXEEBFq5mkzGwA3f
8qiLsg0Iy1nZ1xvfprlMy1uMKLYFWQTpthvPVZfE2IsAeV6bEtx1hqY+MJaeOG3hYnZX8uz7tmcl
nGLlKz1pyorheJgDI0EESdpk2FF3y2Gff4ESeCWbR7S7AmYHb4rrRPXRxBS3XQ8WwkRCIUx7Xaap
T/CkA/QujoQW2eyrMas28Q7JFQmZMYaQI6PMMlcAqw0qJ4h6AfnBPGR2Mmds255vmeUn0MNcaYxC
XsaX+eJPJZj/1h7s2FPoud0j9thGHM03llvl7fP4vhvrYZttX7A0Iibt31mMOnFGzbFWjRmChZg+
zi7UAx6DCJGYFn8GsP7axUkenbutYmAEJKNZlA511OnuvKYiLnHE4SzsquO976wMbq5mkL807UUB
e/4p2fa2ZyY3NHMsWMDL1jupYpc1gL3cv+usGpZNYpyO/a1qSTCoPu5uU8MJFmqCFktriL2MN8Ct
L9pWlYdeE3xz+K8HRE58gpe7L/rSJ7W4y70WQ+/ut8PX+Gtn5JCMPVIwk+ieirN6lailk5YcZTuU
0Lp1LlTX5MOO5m0+Jj1W6EiX9OK64Zpw89TAjGhfOQ4JuZ5/QOCzUKbIE8bpGNWOhOyd+5OXA/Ah
N0ShvccGCYRGcBux3LN9Gr0wB/Ts1L7csokQqXh0Sr9+rh/6L0zgNuiev/I6qK1lzy1XVqjCHRHd
UaLHEKqiCSQOsr29FRE50TzQxmbXzDG28mgG6GLhFFZzyswlDBbrJ9hQgMSI7MleqKobClhjOkWz
Wt1C+bQOTJu92+w9mMN1sIdLj78n3Zi2xNCUTVhEmiZsizt/Z2LHzI3jHvybnKymUf6803BKFw2m
RbXjIXBrUGBtf3UCEnQ5cgI2QUTrhHo6UaKsLieIhdkYWF8wGoBTbGa9l1xrWbjcD742DAzbysmI
ksKCQi+/rpOu6aKHYiHbNGmOeOmvZZcPUZlBWpc/wZs+kuZnYsU8ps8ETzgNM23mSpx9y2MjV4PE
/uZXMqp6G4kTR/GTNqRoPqrhe3cggLpGV2w7/dr3dy1/t1JpoO8Pjci1NBDyIBI5Dg5r+YyATHo4
4tXA1aXZTej+9bXyum+ax9JoUfHlRsqCT2E2oNBveuXEc5ge4wg6y44makDiscWs6VXFjHrTj9U+
4v4etaZGV+aSeog4DHWHNTNx4m+N6mYGVd6ILrtbVKQ49WbcsyFTSyhMlpuMbH90cx+218Q3d0GC
aCpDp8Iw5ARSVebN9yLl8mEwiMWtNjiWjE1/enrjFZsAdEZzgYdDjrIVlltyTNq5N4isNpHbYL3L
ponwYJUKy9awBMMG4Evj1/eR42ID5E57SGh1c/8xeTRAwv0iwFoq24GLCThsojLz3rP4y7orEen7
mWQmEuCM9U32WzVpuxYq1i1h+bL07uACLqP4H9I0oveUFFl4fOpcu8b0/+BeWlvxU5H0cPQ9NiHL
ye2jLSPyEWWwBPB0C1AyfoJl+K+j2XfdDRGxzOOfsFxAkpd3i9lc+OR6/MnW5V4FLG6cJauEqMbx
jD3h5fIk/Gi0Uf3DwqKrYgntCoJ0TonR7x0kTHrzs5+JnBUZ5HRouFKDk5vVFrewroq299O8GXER
lpOa45WRxTOnzqRBm/2/cakLIeRmYgbf+VbFioLJ0rFC2x3/UNdcPBIp8KuHfGoYcnLEEbnqil9f
Brm3nqTu/Jejnh6oqxSbW93JXz5QyPC3YOKpRX5Co4E8MyV1/n/AmGpFvvwprRTI6+ATDrEm6sJ6
o7nT5i/D99UyDBUs0rlZoDDaBIObyOJBD+O7jzVQ5ZdPkkPHgzj3T1pkAW6GWy50jZMaZvvSF3iN
1wp7+i08dQ+hE7qi9jDkctULqelJ7vcmxtUbL5wt/kk3MJni9zDuG5eyU5BJW9V5qlGCKQtWAFIX
fiD46XeS1qhdHrW1DgfI6k613LJc1kgpwVl6y2wiwXiZhIx6qa93baStiXyT5SDWkPFMS4DrEWHU
ZR05iEdP+p/0mZQw5WEProFEi+2mMZz5NAngTI+mT+INoROmW0PhuwjTsgIg/MdjI+PxVd7sx4cD
KhtBfyruFmFiO+CWmUnWVaEWP4EOKWPXUAnCnO1+cdBij77vVB3keQ27195AIWpyjE8iURpcVDzO
G0hm3iFD+pvcM2VGYi1QbUt75PpXECbRlnxJJ6GhhN3hpIY6JjwKL9d3S+N5caiTgXhXCTlVSJ/u
mAqsb5ckDR1P1Bu+CWk8Inf4MF2HImomLEuzfM4XCLdSVmTezShDIL4kEz9sk9yonBZbuLYZgM+a
oPIiTigqDMVB9bafmomGQr8T0bf/FgpN3t690ibvsjTZN+M3hOyBftDNa5S7aix+2Rb2bPyXkOS7
Zx5Za1gbZHznUDO3DNdGmL66wOJGatUlEZuTpi+HJaktGCgDoxtnTQWBa07oRUstOL7WHEBKmLvc
BfcJGs1zmtFyBzSGlXfYvUEkb4ifLDC0NiUAutcrfiLKaFJN4OiazOtWnizB9/5jgt524KShtSKU
VmuEoUYnDkAK4XsxQKQiP2uQAZ9QmFvvWCb0Jk0iD2Lks6HCccIgLH689RP7YgpcQj37BbUguxUp
iMAjaj06uxGbyeQmH0jpQR6kB3PfpzzKe4JvppE+19DWtXupJ0ZW5nHTYHemBWU4mlOjakn15sey
Dpsdc2a5wjHoMEzRb0uOx3MjUHrp5VlVAs6td/INbHYMG5nu3EL3gkB5ko11q2ql1CgS4nXNok25
i+vCgJcApoVLusaEYkZ2YQM7LPvDD+mhJESkqkwlDuzFjnjiLsYMFYNt45E77ggequfWhbu4isv0
IdTlMsLEwY0FjIuRSAiao1FMnB8aQe6WQzWZPx6Br2l1Drr7YgL+mXunuBlkkN9D1/mFPQ5gjlSL
cv450a1L+wzVXohIsZC7m3p5IR1MWGdy+uUzLbjUQ2lbgYH3+hrqRYbJ4oKb1/bFQEWx4aYzjeg0
n/kuJLJzH7ZuuYM20ppqUZggTKr8/dhQ6TIynrr7wXKFlRXHLzSfyu86b5H+lEz7rbmC5l8sSQfC
j+0QV8OA/2kEEzz8rNwfaDjQj08VGUJLyJYab9b/NlMNX9uQoRgOgmTZ3JG3mUjN4T69xObfHGb3
ZzBYe6wuQzwNEb2xBtDpjAJFkFETvB9QibUkIOlCytDkH1kmfjsOkN7lJi5vEJn9Q9LC1MiqncYh
2gAIj90BUVNVxwb/to6oyWsPQzrkdAUllse61G2v6XMPiomiaYYXgBU0EJiVPrfHCA0vlV0gK0YE
DtVxRwWc7Cg/MQifDLsPd9fmhz7zHxs0DsKvZ4XGSUbCEWtV6CBDmteWzZx+tixjzgk++eE5lZhX
ke6kiJ2y0bmJJhyBKG1AbVNLOYR7+oRKtrVG3Ra8WRijESUV1gH+TUIK2RoSayTRj9R1ktRtx1uV
c3/94lXt0MuAZHoZjuGJOiq7gqqCi348UgM5BrJRVaRdX3un/af8tnlH0gw98Z6EBhyBbsBJiEiE
DxKUzPcg8ee5XtQTIiugbX06T9yH6Z0AFZKWuM0kbWEKsPQ9CyIwaPb3YOz64b01D+G33W3k/U8T
SHhRTSvOfSdfT31E/qqRlikbBhcGjlJ/XX4vJNy2ADSj+tzd/+rj1c6+kpR69wgF3vquGSslHno0
aJTpup40t6L+CVGUULhFduSZcCaykFTV7uPiHrpJh/gEg3f8IC6qaK6iGKM0qGcx7NUZ+2/uUfU7
8iXT48iFzKQ5VTnf1etmR6TH3BF99syM0mAoTmU6vXoQry3nYFS+wKFhAAdCQM/H/9gSbZDA/Em2
FDVM0kTWC8x2s2n8Bmyv0xnpt+koWgzZFpA9GdDZEZ7d6dKhxZ+U0XvzgPHIl4WnOfcPWGYLkQaZ
bStyX4c0ZM+OBXNp+oTplylj0BWEkapVS5MdRLb/vjhwYrm2585Tn4xioIZLPr6CmmXnLs67W0iv
B7HTR000xlZ+V3KsrhzoLf8wvtJKk7E/vrTfsv9Y20XjanIabbXz7j80H3wVwbrl6yHwKntDTftc
5T4UWw3ZnxWqtNY3JXEzegOXafZEZlZ836i0IQ/D4d0XLqx3ebGu/s+AlhZYmAw2iviptItii848
r+6HEkDB1GOu5OHnKhVLkeAILpNfy9pfTMQDpAUdvoo4YX9bE2GUmGYfIuo4fRLAmpsySCNAanQf
8kJkW0RwiecBlnVD71rGJNXQZ2JB3k6CnPsSbl2giHdB5JA6QM70qwku4ClVHDV3UPDDBvhvX/wS
Omd3dsrrOKPduA79VHsEJa7jc18oceeECos37bqEGUBGoliSdJ6l3R2Q0qgG7tKbU99NZM9bBrY9
P8+Rn37TmFyNMv4IMpEyNKHoT3SmqwJjVxVArEVHeovyq/6H3KIKPV/i8/1gx9fZhAlGYjyFSfFo
g3z4Oo07qOJ8LWtc+UOVS7rt/JJKn8U0j5edIRd50ZfB3CS9+7YlNjCeBuZNjvZ6dKj0H10meXlA
/ihoCdpWE2BFbOt2KXaqe2/Eh+PX2+MjfxMqJiGeiFLTeHTdz4gzCAr9Jvbu8CwVZBS6vkQKXpeR
AcfTphTfKkqlA2mr8y00SsguQsXGsVUNlKAXL/V2d1ddkaPsyJl10AWNIwWyd4BT2LfodtOxuBRx
9Oa7n19ck9xYF1TiRtDnbMrxFLoJ9JpBtbRAPHdM43ahkKO8HDzzqU4TeahOX90ttWcRXqU2FdaR
8xG52DLH0Rd1K37TYLyKdYDnjXz3REdpQyX4tpjCo7v2sxnzR8Ngb2X260cXrLqXBZZT0g2U8Xt6
4UdjWVSqmHjlh+wtutslsGUv75TTUSAJADCJdcXthU8aWCy5nvkegOmTXOrjgfAPGadnhSRNdJ8t
05FQX2AA0eim2R16CC9GfzpwIEXRcv8I98qNIkfe1E18eisKmj60Fx3Ml+METRiMmWsN34Ki7rKM
JgNyMWjNU6H7uUJa9eKMq3YUQTL+4em6vJqjtaLmjFJb1Gw8hjZry3o0G+fZCYd09a0gZrokoxjk
/ygtWsWOYMogNSd8dcXTSDnSPV31ailCaeWQnnFy8mlvCahaEL/voFM6uaDZJbKahVVhnnwes27t
jn2AySIEK47VOskWispDUhwGp0NS8oZj1BPJxZV7fm8KktYVLtUFT+IHscR8jSfYgcpexUBh6nbE
glnwt3F7Dw1ohGvNMbhzes1ROuJQKcNiILt9DY9KoawRZt38LeyBG4IGOiPBgeK5p7c7Nqm1+Pfu
nxJs86A1fhydQrwmaNmiUT2r1n3ukUHu73siTbUYOqUkq0i4btTV40HRVOkfqmpHfX8vNZGhQo85
gdnL3d+Yz5y08OiB9h96akgDRcbsw/RSsF0qHY0o7eWJ7u/xyI1+uxlKmhZJKqx0Q/YioDohtCgq
jfZwYFlbGcQMGlMimhSVLRM8d6WFm3bU5Q1e7gW56xxp0Nvw3nfVrnUnzS7/NAkzwKFiuwmOVV4u
by8rjoa5k/0ffOCdOPK4qYHIpj/YL8hmhPqVckenw12dNwEBR7GvNbDtc6mbcPqeTF48swX2z2Wm
O4n49/TvJwEPwA+Xz7340s9VbYVzankAuA0TUEL0Spw9S9QwTapiyRu2sdsT7d3/gY+ep2eewH+2
9NLy+SXHvzYhE8kNxBumDU/PGvJj05LDTCvjQ6AwAR35n1KkZ94zdoh8wX0Uo53bTXqfsrWXvRfj
joFWnHIQuFg/f3v+tc52+yMU1bBeVdBY1S2VdFxgbwPCybl3+Zba6zsChEdjLC0+VcEhUMuzPZyi
34oxqPt2rZMXyjrvzcP+B+/SO7HAiOJNN8BMAhn5yIRTKCAH9tS8vspQ5RihIMtrbjF4uskLy+BI
P/ODF0qQQaWZKwcbTU70ZtDXSt+35jAJHSqdfwq194efaavTWIjlIsddYie6Cc5VvGXqcHPNdTgf
MPAQvWpHfzuqXuXyqo5zkXuLB6ySsdVv6RXxw0X3ZqRLjcGuRiV5DBVADq8M1Lwx9sib3eGr3sH3
wrsiCTYNWT7wpAXhr2dovwX9dMq4KjmUb0HTO8HCsRGylnXlbPVutzrVd3czFnyWTZB52sPQzKhZ
ZUMpMfGZ3TEFMN5h/rHdvRN7GrY/QBKIg/7mKM2l8pIg8Qw56Vpw12WL2xmpvE/lKstt3ADyzMTj
pX70PTo43Q9RUszmcXVPcGl3zPbuoKtCMKkq09Xb+6ShGe874PHylnUEG13GMFbcTTgVb09CAvq1
bxwGOm/6otjdA30h4lkeYE3P1Qaq8Aa+5lUcsLTagZG3wxYboEkf7sMoMmJWfDVV9mdIdfQv/VYR
95dTvAz+3WTEL+env0AW5ed16CSV54P0dDnTM8X+DGirx3C9ftFS05MkhmRVKFqMswXPbkUxOF/P
nEjvzzQj3yXzSLpTvxZRO1GBGfEq8Qp+Oh0+gNAuyxvCqJPWojMZuRE4vDqwdkVUe1eid6OS/hj1
/KmW48wyJFL2ZDXmbycyNRg8OuOMTnuUAZZid6PIHBV/46qewGwHTcSAE/hVBShsBLMRQnITpPHH
9WyLUuSOzPamM623T8UMJ31776ejj8YjIiqwzV/bD+ZFhSh4b/EHQYHhyf/pVyhKIQj3vAEatgOf
LGler0QuOcwMrkCtqSTlQAYVdIKC2iAduYC+nqwRKe3BmXcSErXon2ilZuRgdcelXilSBwpd+ivJ
9FAy1l9cp4IXIumS/FiBZ8vfr+2CMQlda4i4lTJ/X/6ygwcZLGSWPsu88MsQriPVZ3+8zZ769jsc
J9vjescqvWRSkFcPYWy0UJ1CexZzT3rrOV1QijqZuVFVMfTdyQi6GHAt/uHVHebAPov3o3x1EJtf
pIfE7VkS92JmwTtHZQz/UDENYJUfysGEPOJMAZQD0AOVPQRnJxfNDVR8aU0ZcY5KeZFQSvWTmCgf
Simt6+IjX4Mx4VH36e9sT36DsMPuURXCUt9RRDSupCbRK8x3JvIasAIri7WHtwlPN48VmLRRKlUD
YLNJWf92UAxbnHp0LgE7jdAoX0bCjvgwJZbNT70ysj92CrWFqJPHIXhkIzUWQnCvPv6sUQQ2yT6g
TNbMLUhQ1IBU2R101MLz2gD62/z2b3iLczqaoO964PNjwUPWzi45/SrU1YZPyLc0zRY1+o+XCC3g
qRl67yGs8ekd6a6O7XJtwM9JRH3XfEiTwkVeyh0Jcag5Wz0iroXdWEptNvVq8wTxCw1FgwjES/Qy
xrxxtcAYCzF/87hGQn2uEsAFUETgEMmXMzeE1Y3ME+vx85/3PI/bBqCrUl+QjY2bB73X3aLLVuvo
DpHa+KuisH/2RS2KsY4mfT9SLLVOVj4xqUrHB0VcZi1gIsCwicemC3J5hh0cpgrOOuVTM9CW5wQq
fd+zwJp6RDD5vFXoY/Vw+xi4gU8nCn7+r+gEDHuUFGKt0lqPXEicBN++0OntaCSVAeWWjMryhoGP
ggOsHvfCjofPE+Zm0i0Wj6aHBsdwiF43oSSrvivwmKuNLXge2Z4gLC/g6m+kGHpY1Qy23+b94VP4
tMrMB3s4IIELV+pZdTcwtRPDeDkdadas8qg8PI/gnmwbJrLkeZojtDayUYPY56dFs0J1Mf3R9eG9
sfZ0blG+vXdjGIm6jfGoIiGogPYICJNtpJmWYoIJOv94ayMJHfXXfxRCek4Rss/PUpMOJv7m6BxW
B0/i8dmrIC/pkzj48X+hHvGATWtTyeDEnD8UDp6klpqB1F/+8w2Fk2/UbhY02qzVUh0N+wjrARvl
Rh7MOdbFGRSdiXU9hq2orFT5Xyad+oyDYcBuoPcXLZF8yNED0mBUQOMHNSTSXq4eUjqoO8Fi+wJs
C34C+XJNnJH8BzLnJnVYG5K8R7HgIM6LqrvjOHtbn9VY4x1x6RyegRZy+VN8syM+cQVjPJozQiEw
4uCV7u2TF18UTCSk780RViXPFXpc5Bs8oUpmbJBg+b8d/Dt+WWILDKDSO3vDvb4DBNiagQlHhXy6
gxBErYVb8HG5iMFE+OSx33UUmxHhdumsF8rCMzGDYMbRn1Jj6f1goid5OOtbmQwEplhWIt7NJGue
S1DZpEgWBOu9sVjmkDgFsp8/GsMjcB7k2Qya6la5K1O/mUtaMxuiKZCxmhK7PO6Uf7RWT9WVbYvS
8gelNhi415KzC0VJnM2b5Fj3LsnQNrT4qw9ivEW5hlH3/88H2jw8bphhLa6jyXKARGIZyO7a/nhw
KXfJ084EgQqj18QMJ/OQ/EBRSQ+Fy68roZcZy5eZ1sbD58qGKj2DvlnC78coFHtKEsMKGhWA+pXQ
8tyAfnpnPSPQkk7kjmt8M/LHQNjPD6ZqoxFdBBiKf8OL1ONJleazBeuhhasDSbonH6iNTAUKY/L7
2aaWfjsaz/TAF02sbbf3S3akXT/bpZRnQgxqXkmFmnYffgvzQTXlK3+Af7b/rNOhMdD0uFF7VF/k
vUFY/yo5qfKW68dPsgAenj0H+qcnrK5jcoazZnNrSeVSx/uI85xWPGphpioCMfSDQXG5PUGFeuaI
Jgla/r+shAaS1acirKBuGRHo9mfb6Fm2LJUqq208oCO7xCQWBZFD1lQYeJw1Io5OV+V/vlOp8tnw
hKcdfOsWhAHykyh+555/Bf8B1prNDqOu88WnilDbTVZ0vYsAlNY9DwKqj4Q4AKv7Ce2l/yDuj+uX
gT7wAWt405bV9R0w3bUxMMwF8GxUYrzo+v/4oMayN7njLFwzbRwN0+TFCgImzQv8UWKa5bYN//i9
M/ZAizKh52oz24IK6RPyhftrqtEUU/KJNusHpQX6irpNR4gxCHs8d8f4YbUXgAr7Oaw/gC/H1ysq
y1Glrlt+CXAODaEVoY8emL1vCXqyKc1hdwwMIAjOaPdfYvM5de3z6TqOWpCipjDwmxmDBaJo58r/
9JfJQS0fBEqJBhlom+urxl6Knu53avg5JXNNcV7j5iQnlR5IwmRg4IsruyCOK1RmQkws7C+ATLER
ZqyZasDxvijC0cM7w/KTOb9Y2awUTuP3qKYJUiWiubcz3knO2Zgim0E4rbqacJ+9ihAgvws4+3yb
WQZ/rStlCvzB9aOZuRICbY8wopAD96+6Z2KPIxKAN1SSt+9+E5PBC7Aza1qA4+NSeo5+nPubwUM/
ueBs3Zsubk/eRNCX9+X7wg5JA50D0Ds02FC7AYLcauZmLCrOsNIg2uWgsG2jvjmhlXkHbYhqoEmp
ylt+d3KG0e1Ypo9kJssrQJoZ5RENXaJq44lFqeslWmZuv3MmH1XGcwYFL/UhoCLJUY1wa/uNENNI
S7j76qCHgRgVTrz27uQVFdqQgaGGRjyWQV6PW9d7T36KolqPKtMAp3iG3NNjhiWgX+bL8kn+y/ax
5ZuBjVPbANt9mozbBYxZJMjeSKVa+gB1GUUSREpsxk3DP/dAzQlZXKJKbCZQeEm0fjFsTAymMilr
suvHVnkOTJSbc9bhtgbwTQB5J0oZNvmGQgCKT+lF7cryZ56ICeQuSc/OMAlJDnmLRSJP4hsH+ujL
143bnCG+bRP3JTr6Ch6iMXMGRwSMOvXBQEa8cY0H6MuARyp0nCyGTqErGPjVLOpDVz7kWWwOPZ/0
cGEwYgJ4ZU0XNVnjkbJSoGfkRynZOwdC5aAabQP8TIOewJqUQ8U3d8R3kXhSMsjQw6Hyu+eUPk0n
+mYBj72RwU/8mzRXj7jnfAYR6mE7usFXBZaQnLTeGLyZ+qKZbrUN5+0v225KgoIodFvXwDaJamEI
06MFQ2RGKbH7MXIHYm9CbwoiKstDEQFX0MhswwZtMZ8OfvrUS9ck3Bz/jAjdf04Pnx5UshFufzNe
R78nUGvrW4JZ40tSgk/e4VNDnQf2Ln3CkUQ3dNBqx5RoJUucBUwgH20mJXAIB0IWiBbBKn3HVZHB
NTTGmZR/6bbpowqxDUlGRTKVFOMBDTQzA6LoYmU0kAnC9tCNpCxVEuEMpkBvDCZN0IyZqt5gVRSz
WflplctqRF0pVnyD9EgETZS/L23zc29So5VrAu0bShjMtTpbMHkK1Oppz0sKo49aPdN+v7v1ClIi
EYwvPGKWRB+aobevKy1Xm/zL5qqSVC/WYhkBU2qobF9jE2lV+tcQlvI9BfjEYGrdLfl3kOXOD4du
hO0YafnXIGDhHEVdOnXgwZIccVjlj546pIjWA4nXitf2Y0hgSi1q85MpEevJIo87uMYh3lCG4Ugj
LkgqIgtdiBsLZeSg7eXU38hesnAW6Gy1MNeiEEWa1uwtBTjirjJOlfE05oFG1/O+QH2/kFNEMoy5
10uKh53lLWjQHkv4ly1o6u0XPuOMUYBQQZnrXqTvIEakoDt98hV7zzF5kSDUKw3W4yoh9/aAMVjr
25P2HCszKaVTSyfR3f7OloYPMXeo5sV9pmp8GmDTJnWLDOcSQ/SlK6ckRKWQ45GS/r0C9+Reh3MU
dk7NTII8TE/SA1+YiztfCs13axm5Nbw4gNd0N/lh54GDX6FQNz/uPKb5ZltapzugYIHAwvZzUm/2
6Z++hdLKYA5nVlqUHD0EedSNFn5+B8tZbLjGHX4O1h/jBYIHW02Q1e20E8slXu9vNicZENItwjy8
L/NZboBNYbpUHmsf98Qp2y0rlcDtWNpdP2R/ad3p8Gnph1M2fLHa3pLpj3pa91YyJbqDg0VB9n0V
uzhxVQxayZvufO3ev4/s1RAprvaF/PCd30Q0DOzwfS//KfYC/Ufw441VVVEArxRk7gDegFd5RinG
2rEeGv7Pr5eVp/F+4P72PwA0nuczY3pdkeGycK/6++poV707q7YAD5AEwMV+LxEADqD5Js9XN0G3
JgARQ+d4W2Tx5cQmQQkuY9r6RF052lxbk9zlqdsF0Ml5Vwf04K7wmWBTQ2B8L9Hf1U7xt6hkKY1/
TS4ifJ8HXTgAWf042w0V1/aFiqHt2DlYfw6hp9Nsku6qfECx1UwGlp7eFXnmIS9Ndz000AL6E3gs
CL/AS4bqKSt0AWclii2DK2nuf3D5WD8sG7yV4aNnMUXvj/esISox1IvPAJOVlZy8RiYygfSMeRhU
4G0ex7apHx3HZMbXKt/nhTmhyX7qs2eKXTX0rtnn/XIcKKXO5iyFH6ljGKo1jgfY/VAMDsxk+cRQ
Fk/wjjfPdkzeHWYy7/Brjfucay5I9IvgmpbN87HOXBnW/+gTiT96E1539embcqgPnik017tuZU8f
pnSzfSKFWiz+HKwTHsGpnVsaxzlusoxJL69s8Zci9OREKy883FaT5sg++iNUsgqFGbHSn33sJZ8u
R9379gXtj5tUhRqMd+owxgdw607N0GF+wKfAlI6axTcZHrKandxCeLrfV9qT49G3GhiIXmSmngED
ITSxS4w1LUYuUxoDWNaUhK2F3dZAW/wZitgU4NgUoavgwC7lF/4RT+nHBbgGYowTEq22PEDh9iAo
bTzvQ/hTMXnt5bnjrbV93cA6uWBbI7kxahgJvFpy1wfOQOHnmFNzOLnv0K4Qf02xvab632ExlFgu
UhJizkI8VlwkppxBty3GSk8ZVgZKGONAKzfgNnrzbTjCQHSiIWTvKKpHdwOvZccZ/offmnN0aa8x
msgOYXnSTz1g7cNSbc6ZvsFW7RF8KwytypdcVX3jf+IC1No8SOZ+d4syy88ai5Dl563yQC6XT0/n
M0x3NWY1+Tjp7PkYrMqXEZQ58wmDKLltZYwGh6gl7d17shD4lbWR5+R9pzkvXHTEhzJ/uvQ10Q5z
AzAgEqKhfSrurMyrvI2igRI1a7gnIKPwsUbRNj3t7dacjt+vMCUG9XxUqpMFGXDc4bIfo8haYw3R
HH5AkqxhzZeTv4m5/nFvb7hAlkgR1Id3kwWOojtQ9IaNv2WE3RnaM5aOyPlyRCfAz5HXfC01nPRe
5dEkYhRwYs9nnId33dPEVTaIxdLNFV2z4xsXql7pioO0PwCvMDtVxzJ4Zk22AzvyWPaL4FodOONe
WNgfilofXSafya88qOE3FcoN3G/7s7gnb9Tl5lsafYl1wtMBG0V2/5Rlw+vv1I4UXo9c6JiJEvr0
PzD2PfEClx7LrlCh3UrGFRE1WZhgf6BiSxanY1xjHznkg4sA8D7cax3jPMpCnLVpqxXb8yBPYJDU
WV/FDWiSzVIgnjhJpta9pT366rYEQdDiitq/H2XVZIQa4QFDYN6VA6gCmCRE1xP7uqgviLico5uQ
7bW3WOhkskA64/IMmnFFuWE4NFDlImvT3I3tGtrohmNr2pi14E8KTd6y5zrXEnlUcaCj/4wwbSAW
PXVeHkz1/zWdIvrEYWbG7Ym8iElVHlT6E2MC9k8y2I0xhOaE5o+XWgYpaL1SDJgV5B3DUXDbuXaZ
9fsvzogw9fXOeNNaea9BSur1pLaLhb6mLuWLuPlFSqqw1/G3DOu9yBUNKraAO9X7DSGsUN/glXn+
gYFkUJ/oGjxzoW6ILZyVXdKzc4dRK4a8PXhemCoZqeSy9YRuwF5+jVsDtOXYdK3bICBV5rYSKyYT
LukJKkq5AGEivcJh6nEW7JMr2UuWHEn88M6VMQOHzHpaeRHqkBA9l3OEb1FA53s70B0BfFp1nucu
vOMlxRVbql+MrlhpcoXfpaigPKmqhDOp1h8SyUtggfyAlhVFoBR991hzvD6eAUZEvBKcRIrbMzHc
OTAbMJjGwLUlSB6Tw/J/+DfOoMawCugmY44b56RUA6n/1MphE+Rckf9I2yEnSZ8XC0pqzV5RaSSz
+bmFgt4RgIgPi2MW3zvNMdQcPzHm4GcB8ljOxszFkZU58AHgOW1XDeBU3K7OrHG3oF3YGCRw7q1I
l8VHwZPI2AkQPUX9N+5MyfIxUGU2sK/FmniCDGjA6eYVSjh33WzpA7FbHbp2PjYoJ8CAf/Jv14Qg
2wMN98ckE98qWQvXsKJHFuMcIdQCv0yqFnTeRdm8S7r8v4+ZwiQkK1+oEnF9CNqIC/xePJRvRmAS
Anmmk7JzeSw2ODCsSGuQZZRrE3YivlZjZa2EuEYUkSAhEuVuzalxw26lkSmYvWxZe8lDGhnlFz8s
o8bo4pFYp9QT39A1c60QOzI3s/VY66N3NyEAbHZMBEK5cYLf38EvCLg2u/1PNX5WLNOpvGW72+iM
p+3BhMyzt17Ps1KJWHj7+evYlcAIfXbgJElO5fV79k4BsYg+s1h+Qc1nh+JwLs1FKAW0IpIUkm/j
Hl9BFJd4g1CWyxhliwkonGI4rhrw+aWpsjQqwUA7d+B4+S3YxmXIecktaNOfbMoOL6rgOf8naMdX
01p1m4Ptmw1nAE9TXpe3iECM0hfC+3XI3OivL1GPs3qNp7/YJWCgbbMJusq1XCSqngxpx2nxbzZe
qFpvglOGu0VjMHhcNx9qVJZG93tkoly+mFDst1f4yM6Hhcmay1M+v5aWzQQAAzIOKa1zwwD4ePEA
hsN6NaEyZ02CSQNx8o/K+n9Isg3B2gDr306bWFWK+LMwd/BB8F4qpvluuX1cqMUi2BmThKhbETYP
gZU82KB1hPZyWgA/P1AAfNkhiYu6Sr6GDyocXq9Wi9EVfY19zQ3zTClntZo14iVAhb/eIpsMbuOJ
3GJ7ABSEnCO++I2K/nYDbMMzyonLkTUfL+5OpuqBLE6SkBTnWHu2gdImX46u/MTYABxeBrVMGQdh
PWYd7sRbsI/SjK2iTIs3J65AIdyJ8u96RAY/DnrIvVSuV41xSsXitM96sHOzNciiZauzx0aa67YV
WaGWqlkI7tu/4cOI0QLoOUWF1uH4+mcmH8IDp94mkoOz+3OKtIAULzNG7SRVo64TSsgz+SRn3xA+
4zoLr89t43lu8QoOHtyduXoxBxlB1BKzLoRjOSrvXAjUA/RWVvH6N/fHCnhKcnw9KuG2zc6XVHFT
jpp3yjbvu5zaLG4q4osR5CpozktZ2yoekj1NRqu4aFYiCrUFxtB8O4mmyd+nV+Ux2b/UDJLgqsAj
I9dDV+2s/daQuonsHpHh9liDv06C+nY+LvIj672R4Ree1EEuA+aWA0nTbPMMKGVgRMIGPpLp0LD7
s5XfogUk8BDqxIQWh8/5mjXfF3GsAZqbNoLaBchez0mKt2gd2bOfAgtufHZXXLLoBuUhDao4YYCy
7zXr49aBdPSx8T6J1jaM4hcWtydqnUMC3ZVHL8sYHrDZ6JGw+l9kGci90e7wkeoPVRbTH1YfYEYG
O4KUUUFTot2WOCOLpg+2teNohOSNtgGp01IxWuW+Hj2nhEf1svszkFsGbCc/Z357D42EvEG3oGaE
2DWOhHQ7yaZLq8J/JMMAKWTOVcOZWzEvnI5hA0xof9hLS7OYFs3Hbx33y9yaZJo8EcbHedDbzcMK
1fwGsuTuUhzzYkCENMSAKIl9QqwAIvMAb3yKzBBOJ+4sV219ZM2V54iBzAEUtXAVdKU0PeLQFRKc
aYpGlFZy4if/zdF/UETYlljr6cTwF3NdIgfdgfiHHMkz9bDHSgxRQgpICasZwwFXLHoe/AAHgchp
63M6x9RX98ZE6NS+mAeJ2oY7drCvU02dokTgdkin2sGq7vdTH3fApeIhIUH4ky2gofPkM7cupXvX
EVdmKoFA2rTTboxcjbIPHsNUxABNmEa+ynf1nXXSuX1FqMis2IFtELjQj7MFx4rHHU55SKCs5UW7
I/2SoRuwKrgCaj2jaHEn+BxUtZNKwM3QVc+TBsbJgeRSmW3U9L9tkoDyW2TfQtCytFA/qPvZwrL8
Xy0ELb4NnYrYlhb8NqkcUkv8KzVxLtqQpVgbqBjpDkKxrGWkPvnNqhQ97BrPVAnFUURS8MI8YX7B
xlEVS45snQaKRzevXNJZ4kayErfDcHUNE1OYEDVlyAhpeSjic28w9FymTUh8XGDsdCDsAUsL1d2v
2ufm/yFebtGKJM78AgjBogJ6ZzBYqWO3urAZ7/rITeN/tUegXO3qjgpOYVvwdB62MPh+0JcWFLN3
jSa28pSEbQszsamg2slcCAduJqFbGE5O/1BIjrh9CnznrOM9jD9JzxUc43U20JKeUgAlDecfDhan
lv5vLMz9QjaHotLqmgGqdOqrBmLKSHuCUvOIWFZKN6bTUbgNdZ2tpehYNaTQEFjryU6Kl/hktQCV
zbYGrZd1Az3H1ZgdKOFoLzmFczcir1ygTyGll7Rf++DkScf5dXLeLhwMGICJrVOixXaZDiozWiRk
3x9b7AficAwM52fKBOzNiguLR0BdCQ8wUbJEBnrXoZ4A7uO6YyrglXYaBs68KwaQQ0XRf/Ny0+z3
MmkgCQgRfPIGSk27tzf5R28b2IX7rSpv59qrTeweZV1tDCYR6EhLBB5lzFxFLD0v0GbAFx2+jVQA
jBM8PQY44rfbpswqGHtsvv2h3WuHl+VrjQNaA/KTxzLylW9ReI9qKrdBdAhQitHz4mzGyqljs01r
wpQLz7DnpvbjaXqvix/THK3JGv0gYN6NagXvmPPlDDuicxwBG0U/MEzZavG4thI1x42+yv0fWUIO
vutpQfDNKpenfiEJFaW3V5q10CXBzNG0ZrlaHbZk0YSIU3JmI33HSO9WFn4zVoDNEH4vxrjN229T
URC2J6i6TtTHkFdayWqGg02eKkpAKF2ZB/RjwfmBGPo/qc2Y3F4xYnOEFyU6BYyA0qbDWyjPTt3g
ECQYY1iHinNeGlXmuV3mt9aaO+TC2Xv6DgJVNfwymDfN3YZltpvq1LkVMeR1tlWhwmaA62BFWoLP
LkiR8sT+TP8e0uIR36TCdHSW32PFUGCYz/cwcw7tFvumSCIMNM+kldH6uyFdt7vFGy7w9SM4gWQf
y+9wuSyEwzvvToctLm8QlCzWx12UrhtuIVGkc43MH55FcEs4ro4EkfEkbBYMVwRfGPA1S5Nqc/w3
Vz6Q5F30qFPPZOLZDyHvhatQaN2bVXqEoY17uR1MTqSfwdUbFY9+hXKCENdLCxq9nh1nrTdmxIO7
Kbo2K0zB+yyzqAScKMY4kFIFKkugUBcD8sl6hvIn4w6yp0VmWukm5KCcG0RZ7pHrcWrhNWdShuy/
5gZ083XyliM0DDNmRtNlzSN9DDktwJ3GlucxMsupB7T3PLNTLoweCpRcUatjGFQOgY4pW2ySSIUf
2Zm4wOwsDgqHtQbKdgVKazJhZ/aQ+6EpNvxRQYi/2kPlrSJcjHBDMBbbnOjMaWG6VRCMZTNWLYRq
EO+qMmJg0t6hxh0iWyCfyrTbttaR3eZcIyZ31HKYQv+WUNB89/O4utr2yY+PKlz/959AkWUc/QOW
r4VdDYMtE4bJiu2rdebZmZ95zEwdgrea1+CpZEsltGXKe+fSplhNXwETVXxHBJ32W6Tz7GvigsIN
TV6RaWh3TamluH3AuyXsN2WYin83e+d4Q//VaCpVNgTMB7dyjtAEghpdWRz+wssvQBhCXXMyHEJu
3hsIiQVJRGvGQzg8EUyD+FdVoJdQTSfBR0SkdY9HS3WhTUksL5kuiNRZa3aiI2E4Z2x6Ru90CqjK
Hna2hYTLiXNAoccUnQxY1P/WZOKuSXwXQQSJU99XKi+Liw4C+4A5ARsWxT8FvNAt4qWn8brmaHy5
DVLwIBi8Rb7wFiYZyV3I686OdKpKxN845+ENAQzJpGUnt+tDeVuK8yk6Kzn0hPHRsYgTI/0ApWOX
hHcXVU2tsQfOY9dRvTbLx+6TiEbD6xpl5/2SOjkmoYWSVKlwvTkrtWQrbit+ZeOjTF+cGCbAhXMi
6kr8oIKD0woQKplrIiUa2AWCQT6Jf79yQ0+iO70nmA/iyq5dgc/rg7ahROgWncqXQ8VHyxxUctay
UjU1ho91mmj2soDqY7mIo8Kzmp57ScpLP4Z7J8uyRUR5qFXYYhIB/9AEMX36C8bkMz8DDYduP1ql
iNWaIf48Y7TtqF36eUeC0zC+8U6FWVK4xahJnExh0HRu/OA3h5EDUV+7xmbqV/270aZS+/A2ZcaM
ML1Z0e7gVCS2aSsvFV5tWhqogDjpuuCA9ml9D4s7RvHXd/NPr5NtIPBU+HHCWThKUle9zsbxIHNi
MzIWSfJp7NC2ov71WAou97I9gk09G0MgxlFVh6V2HlJ/kTFS+Fr4o7I1BYOUGhALJDxjC9V9Ijel
glkUlrbtG6YkYZd+EC3bRoFHKJzx0D+vYG9SzipaVqd1al35VAoFwKsph/PC9L8oPvXVOrC2ziWO
4FkTiapsnJLVGJ1AhyM0VR8AmzFB8qtaTU3QnDDUqc4TlhbgpdGJ9Z1Z1TI9zI4FN0DKsmq5QZcJ
iHw48tPk+WDr9UYOWG6D5ouU00wIpYSmA2Iw9PSCHhnlz2AE8vSYxF3w/6DyFYNNxjhBZJvPJBNp
NQf5f/HyHi7aD7WfS12Iqi//YWpg1oR7vTD8RtXy+eYuqMVW4Ujp+ljkixie/q5WjMeWjyVCWGJ8
MtuVFZF8bFBwJla//DZIxxFVtHloslidHaMMT+t6qU77k/UMVRP9vlKMNCYcVwZfaaGopO9DWHyU
YCgFBYwm/B6MooSitSLv2JBDSMzpdJ8Cv8lOFN2P/qI1d/Xlfjo02MIYT/R2Eis/Qu/aVEMMjR+i
PRDRxAPcXVzzUP4tRwsjxonwh+AG3OHT0/5tBgVXjKn2Q1HS/hKDZrm+HaaHuq9oCafAU0wssraG
RSbfJr4wh7QJ+1oanM5rZO/0n/l14n1v8zC5oFDCFd/gFTqRaV+LKb+pRIWa5gD56p2R02/qe/tW
Y1f265dYOF0upH/y7WWCkyx4WV8Vqtwn7u2or483Uem/W9nBmDYuVMukBeD5lXD3MFXMulycEVVZ
PdgIVfuWyLjcD+7ALy6PdmVL6RCiwFRIBm77UZeuCZuBZ1JinjNl8SzVy4t0KG27SsS6jyo6sm5r
CtWoLtzyT3wJv/L0H9A2w2rEtd5Zo3IqkbHDLjfpmfUMsg7PAxbHG2OT5xxyrh5v0Nfy3HSlMFKJ
RZKtG+3phRtfN5aAxbkUJ+Fe9EDxy+WQEZGE/WqH57hWOLMLZiAmX/9PzLM3uzB8O56IxkQCuPPt
eHWAxI/R55lhKEXgd15hNvWC+xHbSYm9ik+iG80oU7Fx+slkMtifDz4UBgueS6i/23Lz61G4R5MC
2GcL5BkorLFNXz6G/XUj7I9QVylol/xz6SgfO0fSAqVE6ozpNk2aMFjlBF+Is3FgBE3F9U2qRbjA
vlneEue4boWDvXTS7Bb/jWufWVs8tIkDTK6jgG/KpP8rHX8HOTREMa984QDoR9f0M21y85LTXPvo
LZlyjgDf8k5ncpgFIm1AsofyLTnqKF9WYp8MAej2xN5x5ZLwAWgkYeoogRhbg5GydPBI/oL5Vw2W
LPem/dqg9iLsrCgPeKaYktooFF9tNIVoe0LbTb9pwx0JYjBstuzQFuNWSzVg9ucKwn5ry3qKqq/d
BRU2yEI5SjbZXXaF1OzPY+SgjeZNHP1WmpZ19q3EQHoPOgfrhwqcLmznY+vadtbWX/ZALMErrt07
eARmva41MQuXs66tbU2+z3HyWywjqN8ZY4wxmIYpmffAZMGcQ4DAL5QZDoGT6BMH5JHiMiYHHBMg
x7QT2JLL7t3X4cS9dSRs5BCZ7dl+eTJgUa45Z3a/3v92fkmXDTmD6d9XOZt+TqK82lawBkQPVlwb
PmyPFzd0QKP559ekfNzgGzPbOz1JW7VORSN+clkMRo4o3EYltUdVMgzLXqnumVeor4YAqm3tHRIO
oKHzPwIC6dVngWRmSRe4+pccioeRBn6GpW1+0sAU5r4aBUznw04E8j5+32MXcpQJhLv8ykyC+j9/
6RwAedSrf6VLdBWUCaIxg1wIKBC9fuQ2duUCQ67KmU22UwSWr0dant8C16f5LAtqeY3XZz3YIhsE
tDZyX9J/+WPV5Pg+DJ77D5rDoDmVR9fdRbhUeYe8Zi/lw3xYZRwFmItBTON9AueWNLRUwDIacX0h
bM9Qt/TnvwzoEhw6rq2ixEQYE7yLYMDD+22mYMjfrylxp2DeWRcO1rYCxri0+iZ1fp5/JoaFkdCs
X+8B+69JP7G+0ApayxARR07nrzCof2a+kueloZF6ica83eJI9nQWRWbPHx+O8ff5CuCqhMS5CpdT
ho3e8o17UwBy18ydkSMRkE+LhSnPFCoyneA6lxUKeY/1Yqc9bZLD1O5qqY3kkh+a1VDSmguK/ssV
lP87jTHyvWefERpxCiKyfGAAlSlg+3v7AREBKtCYNTMHASA2284TdvflEkd7/maeF9jbVKq+7hiH
px4i7YIXZrMKRXPdHYJcmyu0YcTv0BPE1G7GA9i6HmUcQ+fYVFCBngvZ2Op8HSH0TBCOy5wrMNDO
hCeBc7qoBpgH6FiYBItgNeORI78ySWvaepivcNBRAuxONIXn5zfIWLDf8dVrGVxljT4yKQiT0GTh
NnKcpoN+S0kIGITCtYNltAGdiGMESwXHkMHeWz4ReGjVL/bPLJRfZb9UrpBVI/sNd/VIkFXUav3x
knn0tbrmHVlemoblCPQgAlWG+IRJjARdZBNwdl3CUfPJxc2EJGuhu/Le5rtlYkHUJy0Lh8L2224V
BOE3QjQNqpPpfmIcscuda90m92B53beQGkb+gVPBKWTP3+kJDhwUuCWql4oL8T81hyCxj1FdzAC7
FU/KjYKICR9pih8/pVcSP41aKG6NCkVzFK61jXpDKXrsZuZuKTuucHlDBRLMM7zyeX5JxX9J9YoC
EeU/SW7i7M5fL8VTmgNw4evfv4gY7G/vxjzuj6pwSndCmxH+3wEmq36vYv5/AWvkXoOpbX0KwwJF
DKgm2EzpvmVrUnhq7eVmJ4VqknsFLI9MFoRJ7AC1SMSprJNwd/QuYbWZ4xcomB/NawUEP3NBR9L/
1aBstzV27vTgc01eiQKkALQ0NKeKTZbagVZINQK7u7wS+ZR3lCKuOfGx7kA0VybQGuIENGBmJC+A
PHLQfzMa1Hk+0IqWNUwgRu2Mj5/J9eVssXZGZMVqqVvNdNDoihk0cXWmyUNq7Qpe++qXYEJ6mExN
WXh0/MWnHjo8Nz5QZ7zFG0sRCpiOvGXx11EMl10v0wubZBTRk4ULXmkl4XUyQuT3WuEMR0QkVmPg
zoygdDXyxG+aqH6uxsahpr+NLWh2hwt1ess6tC2x0BHFi6IVvvik/BwP2LNjMsPTifQdK9SNSpUO
0tJd9HA76lyl15cVVu7CRy/9RPby1OK6BZrKLZOpr+FRNfw5bqLbfR2l3eyDs83HWgEht6aNCTuN
VqU9QikiLDhypOsLqUrqjU8pewdTRGPGWtQGJ97c7bZaTJ75Wi11rmY+I3Cj/2huPu8zu8j7oV87
BJY3un1ljhWYLN2JWaABu1jT/0S6+gi6vSwcX1LEbkRtl+Y6EQAmleXxxtXo7IRibqeNOKkic6RD
78NhXCxh2WhB1SSvCguiPxwLU3R9cSrhH7HRFlAa2ydXd2Q19vYyrnA45iX/ELR/IcA4F0FVaXU0
1WtraOWWV20WSG/9rcO7D/rEodlkwneRTqn/ZtIRhf9pX+G3+55Wpi2AsSnaxDlJOOChEnT03wCw
BUHLybBxKpXAbPgmF9roBRRIuboivRIq3mUVcQRUBmcg4kiYjAiKCDnf6ZuJ/CwezW8QpSvDlIag
0hzSvM/C1B4dBGhQvEZXWPt9Zmy0QUXvffa/0VeiSxpPDFJKNn12WYMSB8bfyjM7v45AjzXNbOeJ
R3xPDaqxNhZ5Xdyte5VK95BB4VQdBSv+ZEYtADaZHB4heLK9qqFouNVZNkBP7itAh4NNQTPKJz2r
1Wr6icSghU/VkCs/I4T6CR/F4ZjYRtqJlNExp7jwQU5PvsSCmMzqo3Ca+cxFDtHwq7U4YYgIBeke
T22PGm2w+ls614ABFUradvNlEaStcPtcO9PcfU/SygETwycLTEdDLJg+JrHMjQi0kYXJs5ABC+3W
AeggbR7hR+LACaHSlB1TavHimhl9sP3N8rztK2sUnZ4jY3+MYEmIcRmRJISO+8oqHWk93ilt6hcE
EQRRpsi7C96uxxjHG7psXvPj9cCIIx88cm9r/9id1QmafGW7DXyjCuv96r3bkBwfZkAHxEbIMb+P
u4L+UbA5LZa2ycxtFzt0qQEhnrqUl+jN3hIaxAaGFRKsndE6deAs3XftmF2aI7ard73IUBtwp9VY
QaKGNFgk8NR6puZ6YCyOHmBWC2davgW9fDvV6z3P4vJCzprnP+fAkG3bFr1hFM3fU1fv4VZ/yUJA
b/fPfaQdAsobNTGeZXl0dEcaNaq4TT+gFInz3zJfvfu7FLj+wbMAed1X8D1lLMIneKGOZhPSaQL5
CXc5Wv35FIvCgggEDgQcTcF4nwNdI+6giatGQdAsOEGB3GzMi49YjQ5a4X6N5HU5JRCdyLab545k
/iNq1UrhlxOkkBEguamRX3JxPEvHj3zdQByAfqoASVKLOKkueE3zoHJkMvb9u0sVSova3IsPxSFw
Uv/JwuTTchlTWS4aTWaYOXnogMDBrO6L/a3yfZbf4y2xCX/C9UdQDNB5BuiQZiu0u1Tb5J2jc2Vw
iyHjn9UpnMmlcyxZt3X7rqHOqQSpv4evLKUbt7VjDRosFgMTHBfsDlVPNApGqe8SxsjgsFbH9OAR
9jUYMDVIUcTt3DYrsDXWfGtuiNtM/GV0tvevxsUOOcdTL8ajw8knxvjiwqIjsCL4r9e2RfXwLJ6U
LJ5toGZO531pptGAP0YSozGf4L1r3GY7e9LvhatUI6UJ7TsDZLX2LpByQESzPsYeRLx98KjNKhAg
dONv026xfIa9dSe9gTUKgIQYUJ9w08odQFOk4zbiS8S02cbiRB7i6OVnoTWNdmjqU37fBF9NwVyK
9w0jOLlMtUxG9oAj8SF0bsCqV1ImE7eUAh5b20Wpn0hmg6Qbv+maU95JyKoD0d15lm9kkOEIlIDE
tclz21N6Sj5jeWCryTwbc8DcHV9YG909fENe6wq1lOuTSMRyuRTPz9m0JIl5Ul4NYMA2si2UF85a
437baZF+UXPflvRrjYDIyn17vv/uWWh7PSsCfxPjWTvhGOPvia4Q9iQU2fsoOqPNJpK3kMufaA/5
RWXxocYssLEoji0vfdneJFaUWiBC51cEEmOkGu7C8490/Sp57PnGfg1L+lPIKzPohxGazn19OdfA
f0JYow8KDCiqucTPXrWHxoe8THm23FzLy7ee9dUWEzyfKO6rfGWHUJA0i3JOIjXLhy8wDBh52Aug
lDZbX6ZCRVGTsV29cdERRyv+VrP2cM27uXFqJ/pEevUJ8/TF59fTzvf+qfkAsuHpo+NT4fqUkpiN
v5CN0WTLmdcdxng1wrbUirTZOC5GHr/BYsF2cJJPWkwdgTg4jR9z04jvrGI/++EbmIxLu4aBgYPz
jUpop++YOCCQMRWPYCa6f4LOIaF/m9gb2wXqeoJERHZHyEV6z8nUaJmSuUZ1EFjb774MAmvheEeK
rv1BC9byYn/6EE6QLOGf2OceCnN3oEXpCJ0jeoMJwvJeem2H/zdfngjyWpCBIi7WrVSGuL7Z7IKl
LZ3Y0GbAs7LRfPGHP6VJLiaS7s0Nr77E8ZK796FiKin/H5/QKz1CmxTDYei68UNUJjbBp1EDwdr6
a2cOmaw7v076mQk1wkBOB7gekmrV5sx0/iwmi+kS786bMJBYR3I/DzZNXbfQwLOU3T9k/YrufIgu
HSgMpAtiwg1TyGvS1t270mttVLegwlX0K6zvNgdxc+V+ulMuvLlD63Q3o193hyJFg35jnqGrj8Bq
wa5HLmjDOLmpottZw3RwFF/Kx08lEA170DjypND27ZfJKpRSTKLbNVUTCXExL1QN/+0XnKhCFDPe
+hTDDW4FPMVGMSMx5wrsT7oHm+K/io4F1WRBLEssSpqMRntoLPo7bulnjiYVvIwYuC4/dD8VUd+4
3L1s02ehX3sHYM8vWuu8NqL9CfbqO9RPk7x++U2oFeB+FclQjKrrUFXl45kT7odoeiP37HU8Jo4q
+qJYLNRyAuAEepgfls1IIuCRayQ/Xv0ZI5NziW8eRJ92B2wWRHNAPVNSUsMZW/AhrIclEMGaae5q
/f/pfGZqDvr+dku1gz7azj7p0PW+J+czxQcSAAZwW89DaHn9geEAMh8MiXC8ajF82L0Cbqf9JYMQ
xnGeAmf29elUzS4RG/3lWSps0qnzTZkKnJnYR+eFZZsghGcg7/aZgsWwGbckjh8gHHMBWqdFtHtS
AV2b9dPx1Yph339wozwwNTebziERHAwKwxDpxJvnCr7ZtsoS1NC+BrmbB89N8VZOmbzXBQQZtMIn
5pSddFEKJwXPif7oyZWAcLNfSa6yupl61wtpHEjehn7S5cf6Rf/IQlyxJuYat7IXdusHoOUeNzOZ
NV03oVjuUhdEJpG3DtifIv9+YVx3bcT73uOCrpV5E+PCg4c8dB6sKuXZxyxNg5etmeVUC23KkyPT
oftVWePDOEJTklGicniOE/p/L4ZJZmrSVM1ylBqZcQ38g3FepXiP4GvvKfoIx4Htj7oLjFEiAluE
nePuyYt8/Uc9qud6yckeupVRVh/d2dBqWIDyRhPXgqzMeDr20+pkU/RaMfi2DVDF3LJAeVJ9KPne
wjZdVzjdNbaQzKFVV0x97ah+ula5IlV2Sy4PwFVQsloxGeTfQviIqQ9r2rKLkw5jiDdGaQrqDJ/T
C/heHaVOVMrtTwNJ38Zjr9J/hFKS/y/UoQ2As9tP8biL7qGWS5C9V8uaecms02NcwwSJwuiqf9da
ZvSm+IYkGaxQIo/lZ9qKgDQ85N4CrW8ZHchBk8xAFWkLyAG3dU0c0sDPgCbWZ122dbeeB+INN9kY
yqcKmCchvwfTY46bZZglnqJ52vp4322sgM7+4H4CwSIDpj0NItjxgv4OMmk7B7Fj3DN8A9g6rfyp
7S49Nv4zx7sz5rvJKVP3Zelz88eHaWTdt4hEkaqTpMq0Th9l2BiTbbptGeS4XhJ6vjfu+T0jHuNO
V4sHVAgdlZDZeh7M+ZWFaz07/uXudtmVS/nJlIjai265ukcc397FdoM9C15GnkiYd54yj3cKVcFD
QtMQGl5pToP8pgBz3t4rOrUiryccONycWdIdrFxSLcYw+BpLmpa4bkr36SaGD1Zt8reNnqjDz4cK
c04P3W38f+pQ7laKg3aQlpG2waFMWEcYHFTulAAtXnvVTuifMPTeRR8zqMG7h4FLSgkcJ7lmXTaS
pKRcvGstUjuOKqFb2g0eMQAnjNOTU4ZFHpR+tyaqFmMHu153BLd1oHLRMXfgwts8nSaY2cnrjsf7
yVCkmX11hs2llS67PE/NUmAFQEiWgrkgOaeowg8iVi5fSb51OMnxelJGUU+crBnZBAuM3LN4FCTc
ba6gNaCoI+Xutzc6z60bYz0Fc4Yfk9NdToXRveQKwhlsdlk8ezfTd6RameMHqLxJJ3ZVWo9vlDtF
LF1ylctKx1LaEiIzpSNUQOY9+8VyU2xyS/HP0xK45bbf/V2SBCY1BVSUSWv7kvK/tzMJD2QUg8dJ
NMOUp2kV8qKnYIcGwHK2/oQH0VD8V2yQoIaDDfIKArcAHSvBrKFrMDNgt9UL+Cd+1lCyGqPqBFiZ
rhyzOqQEWEzwCH+OpmnPxWUlKycFDLwJCKCBOMEoNoWS3LAXEOagdBWjKKMmTW5YdVjboO8vxT81
LZ11pluQt8WsmCQf+GlRXS5sCMs9yuRen8CQchnogVyh4bhj/1fKqsL69eGtXbW61WP2sMkcsHlm
4sM4emqCIVUjIxLP9MDA2Tb6O1uNYXzxujHvovfXuNAkrxXhSNTchduaNxweyZSTq03Wpp/QVki5
8Z8Ee8KZdytI6vdhSFlxW/pNu/QkvTN5BxzSpj+As+hix3MGHoJhANZQsLq9iEKpAAzP7RWiXRrk
ChqkZv3wNVI6F14XjpZt0ebj+BhcqiBcciuzgeja4Ng9vbUjhSB5S+gndUWyQHZhcOdQlhdojye2
IW50Y/NGxdWZAfps/LiJ2Iv/rbiu1jery2AnnhcYtO870b241dF991tQhEv8m2RMAm4e/jMb5Rhv
EBxi56+rL6qQ1N5NwfCppVIfUZEZYIbkzCAtmMKsqRpJZKVa38hrMDhngLS4pVacspPetWj2EwDh
ecFYqEB2zs58sTc/SgnG1I7Rk5aeigHpTfKApgTUqS3WvNWsgmIExjqA4/YVUBIebi8GiDr5X4ci
7cr+bRyW0bVhv3QB2ozvAO4X+DYp+/gNDZgDTrELsq30rJlBClLhT5hfn9O7rcIpHeF1jMolUP4X
1oJJwm19sYizWmy735pP5lEOmqnIe75MRxm56Wg1/kxjk9WUZTP7Oo3M5CEzUvoDos0iKhChp+1b
oxBia1/X19zSgrJ52lcOqk4nRWtWTgz6iAYGNoYPyhBt3RZIcYgE8svg1Z7rXm1/zFf2wjk8+jEi
eNFrr9ZeOs1Mm+awNEHbKHZmLd+AA0Ua+EoS9CZgGB7hH5Fp28hfu/gsHE5/5b8Jq5W12Y1e5i6o
AlXFwXD0BEUKLjPdk/ujnEyGGUnWy0La65CyGZKF7EnGEvGPGqBcbdwEQWsrxKAkvi3MH+Yw1q1r
Xod9Ftlmeu+qZZqnAQi4fiHdH/GX8zA/TlVpcFp/Qee2peL6eviKfmwlXwgRl3x8sELOVXl64DNQ
KVX2YHwa/xL3QuHtOsOLN2yXYvYXRavoW8WPt1xZ3th7xPORuVyDlxWm7wFHrLvYOylMZQN4YnS5
twbwZZQewhMVKERJZU1pd3nLeb1CykFHopGbn/cvtjoRKASj83E/IuyW8e4su4XulpGgCUlfiqUg
Dxf/b7EJrrkyMT6Njwghxhx3V90gJ+5+ar0OqBwO+wJriwvzM/poooUSlq5RQ8iTGjtiXvOKkFRK
cuZujpxHRxPyK29KAHBs1J+hEsK4TJkELx7OHjEWcMpu0SgawupgaoQzrcv7KX/drA67+mhZSGvc
Cyo1F+uBwq9JVl4itcRQSX5S0qlznV4GVk9j72TNPRZ7PVmvAsGMD181LdqveSB27pog1+bYn5KC
6YeDMmEY/LtxfgzNclvOx7Z4KCWaWfyQ+ygjYHatS4XW0tJOAo7gr2kBUqNdQ6LaQBLcjYsO62HR
licUoRpYyszL1/QCm/eY8/sNI9KyHn3wWh+I83sx5RqDGRqsZxYnVJ/hPb7sp2adJgNalWD95+dH
4aaz8DOSAO3hebQd1lZDaikkOgRuKUKijq2KMHA0ot6cl1qRkBNjOGmH4lSOgerqQ2chk8/nV1Ow
qea7V5ipfs2NLuAYPfb1jGBxCIF0C9NT4DXhGRLKRk1BYCDi0dgse8WUE4Aah556nY0CH2DNwGwB
buN/6TGOgrJsky3csLRLKPsVPrg9ETW/MdGVTKCmKAWOV3TR4ix3YKpUQzULAGRnD94rRG6o6mLC
O/hJQy0c6V3Dg/V7eynyuusvLG9/a0PIVZghcn/lbFhOkI/bSp0x2oVRrHyaMEeaixFMZTrBlFT/
U8MwIS7uqhQZOen8H6AB/BjlmfqD+L7rlkm5LpXdwkm5rloE/bEGG9ZRSBunSBjbJoe9T/OnKRsT
S4Km7XHN+q6EfQJwKNdgiHVXEhFfkPLeQ6jdwVBbOICgrCT378OpkY7xVmDljgGa+44KCSBr4Nvc
YzYH34EtC0OOSBoW4dcSNcfMbaCERsTqF0rZgua8/JfPeP2yR46+xzk7XtvtsH5e9fGzhUtAse6B
qbWHOdcKFtivYTF3MO0JC3upcleUO1o/5CpcGubqjphzXE00MUZt462AY4VHZq9lX/TFijhxxXD0
JMouHtHuxMSwZQwAZK1R8QIOEmy1kuvMi8c6+oHVmZDFYa2r+oR9uCHv4luWxa2HYDvxw/O6pUS0
9oYTf/TLHPF5ViMPzbrGjbARFTkRpXCUKiuOf6jXXS1FsFOCruOHBbyS+d97ZYveTAnY8F7TWD5b
oiwkRFJEvqYgYLxlnW8jStg1PFEjpggUkcqo+g4OnyYYq9t4A6ZZVIavYrODdyWGKHs4XKvsz0by
bw/pilh4jJhyYvtE80SR3rqZezgkXmJZuHvb6R2vxCw8uLKfPUuJ6molEfFgMtvqZmd9VkUtk7iI
51QsB7s2Qk1Cmd4JjCNA9yIU48byXE/E0kF6H33SgrAj8o0m7gHxGTWNkIQ6zPm+ngYIQlZQUOue
ut/6SL0q4v172JwaGQtmIzfuuFTMoSLwziNTQDqvTo+lgGLVj7kQHiRwjXBG7BzP6xd/HEStrSO4
39CrYQnKPw3fUAg+M8RFt/z/6aOgT39wtc6qByvNJzGyhGZtNn08vYPrxA5aiqW39SOhlx5CXia3
RN1YFCicJO6+3H4x7Re0NPoG3HA56zm4NukfNsSvFSePyVzQHYTTZfbto/DTAbxfmsbpK/d2UUvn
5A7y0Flsl0S7MMpSzW/K9/ciiSeMwSB+dVmjeCanH7F0U0rMdQDR1bd0ZoKFOqqWGUGD0NyEbaew
zRNgYPs/4X1w+g1ljMi5JGajAQc8ZHD0AnbEotLm+sYOXbfFW7ESqU/WxqaJpp31Ngr/x6ijzkvg
Wawrv1fQ+JaJotHDViQj6X7OOUyfw66hos5zHV3OZomBSqsHwgX3OFIhj4svBtKU4lnBq7+czkUr
PAnVy/P4vbbEo3dbvDBMr0t9vUU9LjW8oK++l+18sEByp0W6Bnetr4xDtUC1ffvW0RNDYuXhaoxp
Mf+MDKwqa7v6bbvsN5dZON8Kk4lgmm9ZCbOFaviCPaFKOEEMM7ponPCshA1maD6J1snsb6r/wOY2
Rbzh+tmy2uijuu3OWxwlgMoGBA2wb8YVY8rgX1gu81GYBQy9hWrLnY5CbtNiBkbY8kFX19kBdAB5
EbV/66QFTWrnn5mMHDV+lD+MLtwumW5G0a2dRY0ZswhEN0YWRxPKCsAeJT31Q+K/Qiis4gl/FtdB
wKeEEpigzTqoCj+Vt7JkCYgL/u3YZLLIaJkewloMtiquNGtSQJGWhiPrErgX+pnwPGlXsaRrXObD
xthCpNp4FGe6i76MxyNyCaYk1Uf6hHkzGeXVO0+eZnxyqnCX42izd8h37N1RLw+2NHMSBGTQboRn
7YmfOemF8zjFBl0Q7PFZKEo/ZPvoQbICFr3Nbvtu2JKbLWM6B4JYIQSAer/rQ5S+av7sUBVhlfO5
Ntfm05gRG+BsFdTsM3qN800PxhIcY9crRwLNELpO9/K8XRWssjBzftTPxtvFWjzpB9wsAdXoNwEO
iE7XTrgsxT8qM6nFrXk/Y56lRSSE589HEyOndWDiX0NNDddbwg1LrUszOOnk1+PZIDCB0ivdyWsg
QghVg5HLnupY0H1rX4IYciZvlZOwfCX9WZbeMxeP0V0u0VCgatsEbaq7x1IyudnWd6h+ZkNyr+2W
Koz3TgyMgqhCKqSZPAeagM2o6LvRwtts/DqcMy/rzr2ZJGm57jJsVobHjYnhxM/eqQMtsmwrZvbT
QRptB+UpdZhkgFlAqlB33ykBqaWRa8arHOb3JAhhIQjkNdAVZGjNaDxN2rVxLVU7EZbRwa8ed30v
AROVgcAfOqb9fLH+bozaRhDmt5EHSCtbM5kUF7SlMw3Fn2VLh333GZlKCgAILCnP7YQwuAJmVPQs
9DbIRrKRlbQVavJechERFZNZsqwc+zyg98IjLp02yrnaQ0ApOkBfRRCurrM102i3sxuQYxXd9OPS
HicpPpD68oabyGKzynqi287ENr3zneKZhKctJ89QhyQIbt9CsNToXJTUpRof8ByAiU6cTlw2l8j7
FWxnUUt026TUHzqR1URmpxTe4uBB3e0rsM6x/YDxQlyqbRdxrVoShO7yv2eFPzHzWJDLtVPlxkqe
17gYQWq4+dFfyPmCAOgALAN4bqjXrAx9XG+eVc8CBkivqORN7bMUXC3JQChnghW4x9crVj8iyApd
VnlbGU4RX7bkBQxaJJDznF4xPEjx3kexhc1FU0iHh9QP0w3DnW1SZHEJfnJB68CFmYNDqOpdrXR6
4iJt4sxHLRQDOmm6j527Cs1DGJaL7SWgdT+tZWG95XCIkcSHA2/D7biMz+5ZBaXwbIvUyvTHfFsY
6u25vS2M5Fg51n5ckKO0hrbn/ZkcpBHZ7In4Ylq6nJZa6lhC6u88TqNDcYpb+CG54QyDHnWf+x4t
5KMaXaFIB4ejgfIiCzR4vrb18B4k5HWCD7mxaqV26Fyi09Iyho9Exjt1yTdkSNOBhjU4imUgu1Sm
KT4tR33ktGQQwi0L+a7GS3LwDNXZRZUh0cUHWlIHyAHCeSkkWc59ili/6muzI69CZLu5wJ1Z71Dn
GV/nEAirvaN3dROe+jOyOVSiFTcv6HRgt29flAOViEhRhTFM1acDlaQsWNq3qiRU5SOScKEX9Nl4
0iXbQEnUQF/qEW4Q47emo7uOOCUBdG+EH5BPUFW5nMR0Ob5j0hk6ZYD/+exOSAx2j1CXbQNg+J8Q
mpzaivAwv+4Bwikk+FJzlzkKEYVR2+2O9ufeQrIWltg6DVK0+nnzORfgbPW6OTiKGeD9SDgu3aDC
L82StHOb5nBrlRcZs9yZ3wfIwuXM86NOQfEeQYig3EnRjjQvcZ+dxfkAcKQDHvYJwpkjDdqD2VkW
keJmZwbe1pl3lNzQOhHxLJLAl8DfzYDsHxIaQruDm6ljQ+qWY0l8h9LybuztR0XVBE13bexGCPsZ
jahRWC2/RjJ9shstpJq/NtO5p+wwfnFrirlHEMvkW40Gg8XcmDaj8t98k7RgerOd74vZKgPzoF/I
qEgTFrhIzhk3RcbX93VTtkNcx7/4mRelV2U+/JFVJp+VeQQKcwzJMQ0XlfyLd2cpwR4Bew1a9wB1
Z+Y5gPJwsuNbnNq2oH9Wpy3sxguRKTjDd5oI3vXVIUF+4Ch/IYlxZRg0teaVTiA0vo0CV+DIs48K
Ixe+WMw2v1rn1anGbjW4SwvpAoIFFS5f4+cOeyqCHtNFzhjfDa/Zu3+jt4V3nVoe+UeI5UcO4+1E
Cc4thDWxZvpmw5SOUqTzANMdiWwmr9QUNyX39r1rL4CtBrQhS4Rd/kikIiQItDJvEquMycwDi1Gn
DVKEWSy0A274AFOwNnV7cPpn0k0V1YhLu0Ob7ZlxcWGYyp5MsNzYwe8mVa2pfAZ2HK2pbEcxZD9J
ugNBINxSe6eUMLolE4f1VE2Q/TvG4vfCZ5smE0hEePfT1KvBrLUwD9GkBGyGQOrvAnBMfXs0+vCo
/5oUHnzMw8ogr71R7Iz/NZyWASCpG8dhFB0osrO3li1n27viGKqRd0MfuwOdrcE1QpzOLBXfjwHc
OA22AoKBOFM5SZnceb0T+dUbAx8qdKMLRbMDqzcBd91UhUrQAAOYBrIuIFvdLcvluBsQnm9Y4rDU
D17PJPcFBQUnqpjiIRmvWAGMgxiuZHohDiY1Vhy3QI5m9VMhGxgaVVvpCxMpbjyoUNoMYnXbT/Vp
W839iQvBIwI6GyAIUyXyJ2iJXykYI8qIaZkP0Sshjd/JeMbPwcbQG08dl6lKlRXjtUxA6ef4LseV
7ghB805+5Pi1Of7+I0+40g+mDAr/hPGSznrGXBDkf/AlV0nOO/GgxWBdqFQN3qa/7aT9wZKmf+oU
ZsNC3ySaNRGcxKliApmEAu7FT+i1drPo/L3kLhtDTx7PFhAigPE3eJ8xXfJCsV7WX+FVM1Zf0Dzn
5Ffka4WzljTMn9BuPKqzh5OYhyR+qQDVBHbzyByVcIIXmup1dq27Q++uobYpdZq9BWK8fyfS+wTF
cWnFOjirMw3z4CJmCM+1B2/0xv7iI6fo4rbfu+1/fv4H6FO5+KNsq1mSpLR9oe+bEAEGJPW6WDRz
Q1OSd8h7eOYLEcLhZCn9tacBF3/rb2QQLzkb6h8S/JwQsMVrOfUsqQFx9lhJCgPIzi3ybVK36J5s
gBxSLrafHF0vq85z71pohvad+9gmcjrDrU2k+Liesydq2RvVXKLF6KuPFf4/Okgh/XV9uqK5gViD
yUiFClvpj+Plp5VXv2E9n/2R2h55WXctha7V0fzI7n117plO8ADfpbxKEacVD4NNnyHiUBKnYTWe
oAbmvkXBEt4wuNXYnFnZzyjfJ7oek2wjIBTcwfxdygQTtG+jqVLVLv/dPtPKAwOw0LuD+p/3dFNc
cohdHIs+N3xV9whDJzEjBLeQR7eq4+hObnytIslela6MdmmDfmiv/UPdqKPKrIF5ZFmdpOQPnUgL
Fkfms3yyiXWEYdb8zJZ6mauoHFMFaQefqRO6pRQqxUrtXh+ntub6OT5wF2x40kvQERBEsEEdoSu7
FWTyQdnqVzyA9HZGjTOeGHzyIFq2TcxVVTb37be1eecaTnyN19j0B9sqtSGcNPyqT4mvv9NdLPAN
horrJ6fLQ3x2EkAtQEzVI6qOh9hXfSHVxDFoGL4YlgbfiMdKROtzfnh/Duq3To6oHs+8HVZWKG9h
1p96zxcLj5xTPYCBMvOjkKabJBFe/j6a4Il9Re2o322XRgfIA5Nx8c+OIuGnxVnlC1/EsO6xyfgd
aqwOHDPf6FQU/3kbW07O4qhtAcEuA9O3GC8rSvNo2dEpJrrQS9gz5zjWuhEO1QGxzapdYbAb9jnB
BX44j/qC7/zcafEc9czFv6u3MdfXH8GUz3xJjYxMhKdtRvYM+E+nH17hTSunCExTR0NXym94G9rF
CYguFBsJgMnNpeyssj4vG79qjoxDMbeA34tQyW8Br9doLAwPRUtQqZPrE80WuoYlAQkKAkQMROrI
c3f56xGi0DleXmWQfRFYL2yPBAdGIJflWrSYYMMHfgZECZ/fXA1BvNV27hyKUpdmBOdA+SlBWy/Z
GoZV3bw5gWjTgvw4WfQ8RF8Vnx4+PWY0mDjS0BIEdgim0YkPPh82mmnQPiwDO+sM8ND+LMNPQsqW
AtKclFhi5LVAId7Smv1MJ9jv3lOBYJ2LJokH9LNRU6N+J5csLozlwhCihu6HxfmT8hZgh7/NQe8E
HPOTuBUYz3AtsfXXkEdtObLplyXI2mQeH+JlKx11u2y3ybgXhNBXo/X5vj5J0uM43O2OG6CP6+iW
gd9J6Sywo9F2iPf4Wrh1Jx87OC7whLPRI6aQKup0jJ/juC6NWMME3o4xwU4ZmOYnSb31oeE70Rfd
be9OxYUxDmrDKSSCkQ5s18QYfSZ8CGbtA3EWRjjJUm+toKU1nqeaO8hKPh1pArAyHranMh+u+mdk
0E7HbNyEjtXYtgGZsT8SEW7VlrTN3OO19hoYU25Dpp9JIwfZsecc/c7scJQec3x25Dl2CfejGmtY
N80odvP4Cs6XqFo7sQVUiTrebcjL864nhlo2p2VXG3ZTQ3Wm4VQt6E0ekQAa5QTDeCcpaUi72KCq
1x7DT7c7ugwYHOJ6Pw6beTtO95+MNDNKip4suJBV9SM9LM5aHG9UZ09idGdzgdGxRXcXwFuj72sb
6953A9OzHnTV3K5nQl9yb0ilVBh531OvC/+kvaWjTjBPtxxU4JQ2zwIIxRtxus4CUdWYvfT4+69l
OXKRng4T4FCFHMHlw3Vn0qpxKH3MRqxw0mQl4Wz6f6OHD2oKn3kU+hHNe6QDoExLmysOyIdsS3BK
gAvjrLl1bA27eAfPrJoTuqD6ozVt+aqQvR4fTfVSHMP2HwMr11OjPvuA7Ej1f9S0O9ExtbmV263m
3xTopn2llfIEczsgY6PGxwJw9Jp91Ph8PKWG8V+CwOdRHtJ6xet8U+ZNXOrSSfTkOBOLS3uMkCj+
FC+92i1aVoKz90aDmU3km3BiBhcPxjxDfSvTfEfbFYXAyta+a5jWg46NsWZGnxRk0oOEEFxMc4au
fRNBEKUBxG26CmJz2EtpviGVQ+ddgxI5o8NjZeKtnO9TPqzA5tSNp0Vno0Xmz65Q/LKZIixngsfA
XtF1IBC3qgr1fRSTo88HVt08jlKB8vg+jFfG7SZ6WfKI466R361ztQu6fZZ7yaP3nCym465prC6E
HF88Guvo8ceKnDdYvjryHwptT9u0SZqj01I7dy5npE6mvuSosTu//JTD7icL3k+tgSQCA0h9inI7
ux5YEW0vdXHFgdAe54OfZL+73J2SBVyPTtFaQINtK0KnhAnO3fMqhoYTSUVBS3OPqqWaiMnBaLuK
hOpR/bqb8Gj77IcFjlacPp0Pr52K0/jeNAzuQlGnC5GpQRuoeRWIGTdYzntljwJ9IOFGkzLy3G2V
jtwpPIkqkGp/vUsVqVs8Ibm5uKGk+MB5CwYFRquIV7Kzr1gW+1LP6Q97OU5UUGXGJuYfGxZ5ZhDg
4JT4/8ZF/UA+BZQOPid5rXhObRiw6nB8IHOA1oTI2WKfYH8QbpbGs38ivXt9xhHp1thamyRKfE8s
p2ODhhrfCtXeEuNtl3ZteQZANoBZ6Rk3olTvR1lD23PJHZRhXkn0tRAqy3tqIYomMTg1cCpH/dGT
nsED6Hm9eH4JvqCHxKV8F9GA9MX3nj8H9SrdQxEWj8eGDBH/4O5F1MBe+iXRuwkUJ7fPSREaMHji
Am/X8sU/0j3V1o6xac0AGq1NBUVn5uHHh+8Yzlq/QihZT15Sb22uKMUMGI5M5Q8KyJuPI2PMfvaQ
zUTxxPd2bFb2ZVlbzzQMPqCj0gWUOM2Bi8YiChJ1be64mG95qWBW1TKXWWo6xUDsB0eiR23NKaqs
9jyX1JRE2OrwTFMbNcnACPDfyVQWX6JOwNibQFlrpvEH1Eye0cNH64Tgc5C+O+eUVRpWt/iiWr/f
wp/dqiP2PN0BhH74U4lGr9B3o4Evs9fOGN1afO1SspDDIvSS1ykGqiV4cLFc1uKZEaC5yl/6dBBY
kYvebc2jL7OQUh9i982+azXPxkwCgibuSMj3C5yfVXX/9zErC5+mww2LCffsWuIMZFqfYGWcZTvH
Jqz4pXCM7KGVWr+/r+QLLpwPAu8q3/QLsCn+AyDAM0si5X4/3Hsy7Mk/3ggJKBRG8uP0VY2BxwK9
76s9wdrG5JLhEf3ETiyVM2AFeinpJBsp8mtbjJTFN4p1fTJCKmhiyQ+3lPQrlSngaxiBy7x+psYx
xFTbcNl52tjVMCOskWQbAakgSPUy5bab7dmgjlqNi2umx2AEJgXaiGijfj2kikQahOqenrhhtdVd
5mfjWP2KdOMJrf9HMFjtte21GTNrP3SCz2u49zs0jzcXgKE66FiEHESuvllFwFo+GwNaESNnBxVi
prlUsK5OlBlX5dpKUCgcUxVL/DR+Css6Bb3DKMDWJLU9BzUndRwKXWX06NxG/mNtLjwcLkQZhym6
U0SNTFSL7QoHYDL63erm/vKI06pExf/1bqhw/crZkn9/5CI7FUihhjZ9c5a0ziubBumN1GmIRUI6
iVXK8lPVxtVI3/0xNOlBAeQ8ddov5EMCRiu8U6OUsM4J1yinxmeP5zLXfFY2hSkBD0srfTA8K4To
GvmMIQfFwDtV3AQOCNP38Lx2+CciuC361OxWxdmbCi3lmqcUfzXMhVDVeI97nTEHhh+IenT2fm5q
1VL8x/bVoJHjsgKDEKeXKmLTgNrRV+poNuzl3MLcb1fgZLi/YBXyaft/PR3jFOk+Uwttdw0EuYVB
GLW19NQHtYPl0iSOvPN5yFzyTEAxbUYLteEGZwZlKjuu3A1thfaIYmLgAF59WjL2omHox3enqlSQ
yshxhk8Rdgo7fqm/co07qKC/kPlkT1eS2AnS2IpOo24TKZgJxuWqb/6upkrIHGtFhzr9vLWSXx9C
QzE0Lu+f6TEdSbAjFj68I41n8l7+5FhiyY1nvueS8KEuzodaOUgUHoXQNkUjxIoJWsHgJlkoWFGB
V7k2MLIwuQf4mtLqn+OIEBTtaV+80sErf2za39iWNIBBNK0ko2Z+tKgS2OYmwndRLUiLar4gH7el
Y+ULFl6WE2ljneFVSzWIFHAfvRj8vHP77F4EUGwDkpyoRVdK16lSctzs3/Ex9V8dFA/aMQIz94N5
MTfnJmUKAtzrn9SppZufxSI7FDlUOaT95blujH7kEyQg1O0HbTvIaR2DewHNai08gGAbd0339JRB
EwdqGK4FOyBPi43pa91hHX4fFYs4kvjvjZLC9kU91ZkvjcuX5KgDSTkyBND+30sub+WXlUwAgzs1
x6Y9fwkPqt3DZmgYSicCvS2yNxxsIOGXJrg0DZHcYLnowMDcFbChRZRM94cYlZdWZfOZB69AC5sv
WUF2fHw6o/788rz2hGagWlsNwTWqU0ntAHVzEP2pdmxx5f/bjKa/bZzPwRNqWNEvbW9WhUphmbR/
ihhEFljIarKHY8m/p1I5PTgvZVUiyZJSeEsU8GazPfSAHBzEc906owDD1xdOxKjiZY5lyC0Lpd2u
gxopk3mXEjozPhi5coHe//cNizcvd48smnRzSBm3WbU82HsfmPBap6Y+7I1JRkXEO9s/YeXdPPuP
K3r62q5UwXtCXbaDefRNHZQLsO406Ju8Muacn/hCvUx+ok/KLnQPLlTIR8zwPfhHjrJeZo2P/71d
8ZA2Pise1vQ1lfr7cufO4HO/eVmtNRb0iqphIeWifout3A4ONw1pbDqdYjWfYPQTz+nZgO8yAP7Z
IqsNei5ZxLdKY7IQtxe9dPqQ+hzWIvNvFU+BL10ChBKYzpNq1tuJ8CptxHN7N9i0zkOPFPkZ8k9A
iPPxgr0LbPIGEsuXKLDI6nM0Lk4j6g42D5velRUmL+yPoTcf7VudA7Vkz8TDLVSmZmMnlozMDUQS
gyuixARBt4gTU4wQluexAx/lPZRib1b//4mgaQ0IDg92Fg5rwPhZBSWvNCLRS5ndTsn4pOaoYFE+
FyXOA+F7ElF8avQSLfKD2wQAx0HYFHs+d7Q69gTOAEYYuuT5DdzteSXWSX0rUPe37O8zzdRBvdJb
UrgvKb9/vfrX4e/V/QZkRxryNCkaUijqIaLjLbAdvD6WbVN3iSJ7/pm6pDvt3xRmwpSzjzBb7a2T
ukRkz1pcEG0Qfhb6N6ea1HlOHTaVP4+vZXaqmET6NQS5EVnQRwnvGnRpsSJAfnW/HLB/KQ6ZFymW
qJcc3Sqp0agIVWopFVw/icqT9XziMoASELqtPJviURk/Ws28PyjCWwDe188kxaA6dK1lEXSJmVd5
0k3tf/3zhL7f3NgUkbC259Z7xTlzKA9QzmVkdV/a/lbva486k+Yn2XciOMDBGXXZ/BNIsHE4JKsn
pR3a6lIUB7mamngcCen3yE2Q4dYBBeZQ0I/7BNNwFAoHtKjNeO7vM9w5szzMqnuw3r2SzLn/ibRF
YeY+Ovl1+Hq50S0wJbd6b3Kal9wDuTJvqZvvUaR1h1KObDgULrsMlJg4eVarDESVV+vuvQtHXbE+
qimq3twx7pS3Mgr6k/alx3JH0A/aXbiauTeUExhlcS+aiD5XXr8A1F5+eHXbDpBpfceZITNOyZIj
SLng6QsmjmAWFZ/ayhaQMAEHzT5Ku2u8ZU8BXPeo53AzzcAcIc0nZYlK+ie0sx31OfipV8OyRVE7
xLaQhf0FtzJ5VcMm85Vlfza0y9tLYlFDSbeLOaTFRV5hN9bEBZ9pFZqBI+2g7zX0qvi1nNmjAETC
k/iIyNKiF9T5keWw+rZIZjZ2tKOAOuISOidj0dwzm68SAAEs2hM65qx2002vRCHLnFgFytXpvHcx
qY54yudv7pGqIDh5UwjPKr9zlpDJRaxvvQzls9TkgF+XCOtkzLaS00EqHZA/3qXiMkTwoeZsnXtL
N/fZTM8sGZUJfjarQ23yklvGeB2M1zarfnZzxPFPh536XGdDvUICy/lCwq4xfRCWeqU+Qup4XGyk
6Makl8ZcTNaWFMEwtEkY9R0Z7pYGvDGDvbltgD5L+T8nJA3Ff90lXXZFKrqOxjgG0K9ZaxqDmZ8b
5EY2AFutOeDmqarkkm6Ntmfp5vG99hyGnXlQpzO6lG6UZSbwo5XTiQEfgtKWlCZCZkFPZqR+qIym
1icoWD4Tyeeq25JcVkGhW2lzvvDVgKzNBTPeqvn0UFAiWoCTnFQS1Y7LE9l4nAGTO+2ZhY3UBDJx
U1WjSKmMangBhUJNKtIAmBbzRo6FjHx3HGtdpN+uqfKtOBAVVoM7RpYZO944VK/ZXBkiAcryl0bL
LfU7mnomYlYaZvfmIynClvLSbgjqBDqvoZb8n3DrFb0aw8hJPmGebEcwXimDH7j2ljnU1fxu/muz
UvIW/UShCBRl9w7q2Ju7Bhr0NHBr8/KNWYS3xEqmGjHJMQL/RFE5a71qoAJuNgbKMoY5GZcRhhMV
KUaq5OXB2b6jMbhNIypOv95LUftupS4CpYzfX3Prbou6ALDFjA5/hg6ayO4uc5WHHXbfCePhT0ga
91CqhUQssM2QA+68ADBeUI8oSUIvBL6yYG9s7x8btVTZZsWPvep4Yli8cUmI2664VfdGzN2wtAWE
oCPV2++W34tXmzwm/KQeEpxqUHmT+Cek3/CjDBca1dfmJ6IHkAfs2JoO0WO7eADdu3DKt9jbGEpm
MQNUh93pBLXKEiGef3hUY2dXNIedtBOyzBBrTAUo82g0UBGUz+LBl8eiiGS9h+o1iIhRzH9UCBK7
tvnTJh9q5shIiJgAFR3cD3DNcX8G9nTZOSXw2W+UwG90BPBWUShqW4h37/yw38nNPEAw9BYh8dN/
yqGFJHVr/07UGieE7YNGpS+ueHWY3mJ9z/YR2FU4Rg/cKFw8zz/FSt5mihwOD5oVZdE9rfqqDu6G
VN9Qgnr26e8CzK1fkZWJipoVdhW0+jH6cSNF6eifKZp4TJwvJ22VUKBVw/AKmmGYzWweAI7YvDkv
ljuuuQDuEqs/iiRPqFJKClvYmS8qxheqAFH0pc0STuBy/Cizb78xKPt/hCIx4NUBwTUBUUF+1kqJ
68qGJr6S5J/Egn4Awn4MgmATXptb4T5ck3jIdeR3hJhtuOGMyDVWnywB6UqBI8PB8li8kHqq8uu7
80IpRx00wm0gSDbOwQO9t9WC8zVolg+qfS4c5Gw77hjmyz2rIkQlj1oQTd1KhlrhE6GnneBaDpVL
aqPEV2LGK9MYlBcMcEvkOvytIj31s9fqkVfz+tAM6aZdDoxxKmvPoTVt9drbVbPSJF8G7qImfpdQ
m7hqRSJBC7AriVVY0Uo/RAj15kM09XzXXfnvnV8qoEPrRXrAG6cU4v2Wzl29YQPl6X71HT7MXtD3
7KCESu/wp3OxjASTau+XrfNfdVzcYtrN+GnO2e1MordlLjBjDwOyiNcCVtwkUN+4drR06p4wC52b
l/DdoNE+0WGG0n8Wh2U/7Oov4IKZ8hapWcyeGkMvb4n/PCcbSHYF73xN74HsEbptsUT3J1pL7Im5
51hukMAbFbj3i8g+bpUYPBdHt9d1iP9Lih1BcNPfm/UQgcFF2Sb0y4xJhP4ZLs7eh3iRsx+TjSVE
V7G5Y/h2n01wmPyS6TeienvG5HMqQeMdxQTTqF17BQml8dif5wqXP65iDZ+FMuDS4glUQLPU0dzX
ZGl5L7ySXlVEotqLEbDdbyinxHeU4XaWsnw8ANEGLTOu2KJzJX3o9jWXEBKu7sp354TohfsnCqrh
fUMj4RmouhQk6Sp2VXXNCbU/jHM31dDV/trHzylMf8cvxzWUAB9RNcdRCuNTseJLJwaREKq6/ufl
eQ+xx9T/ZT8sYk1ITmqfStCyowv4vUmIpQgyn/B1hwpDb2xWdJKVMvMsSqw1/KlkkO01ywo9HB59
atywqO1SLoNol9xa6CcgDvIUUUrEDv+IhxbsoG5McsHfmxX22snmG7ReRCfhdVsP+/6TF1zbsbpr
o0vbmQhDhuMKfXph/SLNG+Xyi1jDyrE2L86TBtiNglQ6ZNZIS3uEWqfH+8Rb1pTsDbhFeCVyCplw
2H4MI8N2ROiQduPcjqMwib/V1Z2pa213NnU+b7PXjts9hfcPrvfFw0/LaaUkeo9IhitYh+yATKPp
cog7mdpiqMZdPO1bsQ6J+FaKaDsyBqI4lqAyODNqh3ORPHduAOHT3tveSUpCrSt3CuQMM4w/aiSf
86ZlPSCwH4CaJ7Sq05ymnzUX7Su/uPwP2LrklVecv3E9ICrzf9hAjJbRSsg6JgxWGoohDrGvQ7oi
OhYXkjFJMswyY0SQXhHNLEc38atWFxetkFfZ36Fdd/cQw6y3OuWPqAH+Hr6mVDpcTQvOtqzfKgCg
ZG9Y65/VFU51bjhwC5jBwQ/mFi2zAuyHBaR7wzURBwyXBIw8OndnPGwbyEa9VUGVlStmdhbnyuNM
ZaHLSPGsBU/OkbqQ3GetkfKQBHog+b997smQjdnn347WwJVn/gT4O+hE5FfCUL9GWfU3fMa27Gau
S97ZhzvyING2vwUDHcDPp5iQemcXEUONOJC6dgt/0NPDHBduX6v354roVnplonAgOTjtzOJCBZ8D
2z4C79ioU8l0mMI4QKDQSOFSMUZO5GePtO0FiEfbiUmpYEuGYzUwFgUtJshTB2ezITQA5eqWNcfP
EYTNr3RIwuPXMdXRk5d3S+WVhCWO7gBd4hmn65tXLJxRhoTog3Pvw1jbHxU4voH7CfKQOcCklbmp
HnAtwMB76FCfEHiiZng9sR3tzpunsD5ryVCojrphPD5BYulXD/mq7ACgw4GjP/SNKMvZIMperXcZ
edkblMSLt1vaNc2OtAMCnzXzKtj05AkbMz6LadQj8oRIO13sStdFaL757Rn2T5b4DIxbWAKeW7By
mid/L7zCfjQPE/3KlhnCxxOmp7mplV4FPBzU77z60pqgN/RXYP9j3As79nWF6iYWkzhpD4M3/6zV
HMitzx9fM6t3xb2/SxP1LcPfYoyabVkF4VvmBrun26dlTjT53xLe3ZbQAQoC49AxqRnf2nDqtuuo
u9GB6zHRd/SBwiAr3qmxpq4aDBeFBzikPv//MbgxqlBxCcfhbmLBznVrsvzvR65pXW3lgT+A2HZe
389DFNd2IcLt+1JCHhdO80LQz4pZhaLK9A1I9nz20yo+nTqs6cJwkgTfSsX+ddKGtCZfOIdqmCK3
12dhu8f2kPW2vJd7lL6yNPQC6BtYtLpbSV+DmTn41yxDpTaSzgqxW2P2OCZAK3Km9JLniKC9u7qg
/BHX/eQ6Be/zL7+ALsUYMn3mPbDP0yDnsLrcCDhe9lQ/ki2XWDmWe5zt+LZ4QJpLAJ18h++7BrXE
ezNnudpigVOOclBrUUJmm24nE2D1pGEIkvV7+rHFtvtKzQv9MnoyQtzbuiyJERp+ZH+IZWigVDaE
ZsXGPDN5gKa6/yie0RpDLDnKFDt/ePBjSs0wypMNXttBr7iB9p7ZYyKoUy6de9rfn1n4Nd2YOtl7
muX4sxaQrNI1loRmVoQCtR2vk9iO/O0Tr4ybf+6OIhYR9z5rLuYP6uSM0R/tH/MtIQY0Ufc3Lw5k
wKhjs+cJaiYUXe8xElAXwk9mWn1WL4BNZN9qnr/lr/kHIZS4RFLGZrYwAezMjhYJpOLS5HfMQNN4
7rLC6q/333pk8HenmaG4h9pVPBUM3OgaR66Y5y7lAoNhHipeZo95hlvpsL2zXqnyOAycAtjUheIM
BTg84l5wySvzL2npe1mzceuuJ/k+OkyA8RQl6VFNg/0Yg2yBG+86EYaWwhcOykS7cdPPaoNdj9bH
R7301nE0fjMtASHE/mfdalQXSMqbWPNTy80qMdqZsTBOPYzGrZFqe+Fs/jNAy3zCSC7FfZ8M2lR6
bHaz8S2x6feVgGf9WOay0qmZPyrJfxf3h1lcdPIytXSy5k5JIz3aadY/hqclXDjpLhSta2dMJOAQ
C+cobYqKA2xGH9237gJTBPYBoHJN1BBdafUL1K90lna3dj1/HyuWyq1AtOqPa8HKUjE1hjhdjm1c
NlnrG8XkWbk/Fp9M4hsvSKs73WaVF+0HTxqtUossCsniFr1Xuj6XBv7uNTYmSf1pU1ULU8A9EHXy
xb/gm7ivPgaB4ChNYfIoMyUTJdK06X/Avs8Dh1Cu1r76OYQJG5u+Dgz2HUW6ZOGPrYXJtDCTnaRy
tMoA0oKXB52H5d2w3YUZEtza1WUdRfnx3sRzOVN2WhWaHZyVYmJw7Cy2A0OUrWcSBO/BfHk9TsdA
2zOaSsrTtuV3ilyyhi5JeAc4qiouta3nh0CNrY0r8o8bTs/j3PuLoTTimE9BAgpteGyIj0nCRiJ4
C0zcDxVx4BvdRWJG3RBN/SDcsaJGqyIY1BXiruxNxLfYE92+TTpYlrUAfJCaZZ2sLRPFj8UCyL1w
/x0qSY1OZEl2RdT2fapCiVpi380dw0Jqw0am9AF8hKcp9vB3YJw6UHqRXTyr0wSdAU3ePXyIN8gy
iYb6Zrieft84KmcRpvnWnD6kf1IEO0gNmtS93QamwL5p3LzY9dy5y8bgZmwNdKqoVXddKWguu0Jo
gX3HSZMtvPM4HZ/AN5kTvmHeKICXPbk8QIdM6gYocJgLwJGuIyggq7I3g4pyFAvbCJJ3ul1w5Tg5
5TtrAztm+8xM8fI5YQkpMUWH6GgWSGE7Y1S0WRj17QPSkCRWfUH9RWU6N7/02wahNa7wUqabfXmD
SErVP2yqp8lwjHaLcYoKn6Fu5knt15XJcDrZGEy3QoP+2iRsGCpwIb6/QqOu4/E/3MOrnZMlRWRL
urka/mvI88k6x+mKj5fqJwgqx/unaAd/ZnunTdOLPQxjvwfYJIvAK08iaEKj8vcDusTwq+3h6L5D
KBVusTOIaNQaQiIvh70mIhQnjh8DWpVvisBnstgVv8Wbv1/yJn5U2OTh33HIstDC9gIJYTcUVVTs
qxT7MlqaA6gnBl1V98NvnoOjZBxTEZokOLuqz8WCwktgSk24c70NVEvQ0jDVsszWqvUjDwYkr8ZU
nd/eanH5jdMgta/n0gKbVM/iyZv547grjp7NthwOuGncFUnDeAKrgIER53e+OeMD9tSfuibe8RYy
H4Z+Bm/XwMH5GvTbiI6rCNTYeKn+RdK37b9mtF0yQUKhREFOpVun5dcCjdHBpi/WG4wK3iHLPYOe
Eij08orCTYa8Pv4si0Jx28vgzmPShcP6FLQ/ad9H+ek6TIxT+7tu21ttFo8iqMNIdof6nT6Arg0K
FG7gJUlUusSSm/unUFz8lcAB/76Q7PCPKu0pY+YHZoQfZzTu73AUqQXJyEFIsX3gXgADMrG2xApr
qlnErXfzTdGaKHelW7t8FXrLgm48jT6Uga2YNZLSrs4TenNexLuMlmtd4KHHtSX466cnqtCm+KXU
dIkh0yEaBMKTRIijXEo9+ND4mWEJjE4XjlD9LKyIKUCztVqNgz1YDwAMwK8kypOxdHOvqCV9JVfK
Tu4LJA/OH3gEjk30sEkKLRpesqxOGah6E6nzl5EEVSyO02KLycW2b5Tr+4xk7sqjggQDDLBVZWWS
KPqPPOWGw1p8hXPDlmMma8RxU51XRGJG6g9Rk9odY3TUIuonqcbCSZ/ADlnIjhuJZ6kLnga/pvgE
zdtGRvmejpnqLfVZSgHgHuhRZJjQGzBcW5S8zPwIyWoxROViND3tjumRCNgwwq6ob1jq9yaeYJm/
ZrXnN6DGYkEgFwNQQNtpsP9JIRYb6OHISSr0skNjQ05P5J/2nJrV9vR64599wUkv2ZCU+Pb0we4u
4amZ3M2nTMIYm55AACvGczZhND/q+Z4vJ/DTpDGxC9MjAKLkylH8rVHcxwTDOK7D+Q41MKebBePA
PO1tRssaSxEWn+vxqoujdsf42u4Ew6kbMjN/323v+PE7VwheymA9nEt3TiL4jjYnrMRVhOYHVoZR
+U/76CLyDJ6nUkoxE8EyrmecbVI64bz3cDL8uVU9bam7+uQGgiI+Q/X1YGBruy2baBv27rK5jDly
v996FjSoC7tPrRipy19OXaSZXGILVKNcce/WzIJis7AlwICNGG5sN8A+ysOjwF7eMVU9885wIfjM
y3QVd6Q0j6rpVik0x+/K0+P8CW3CpeXTBOEJmWk6XvSUGa+lk+j4RpMVHvUQuOhzg1NpAGSs+a9Y
GjP3HSXquULfpGiU71GgPOkXa3hfuu58eFPXjrwnZaDsV21fxmn1rllQJGjCaAvHJDeP7Uw2HJ9f
bg5myE11nYjfxCyutSVuxfChpU2ENAsAVqiKOqCZqMlZvRWleg7e/RMuQLorzPzR4vYrPiZ7XGPU
LWf4f8sGA5Bdr06/ISjHFan9ffUTv25lJdFMO1z2Y3xhs84efxqZ/oEPyU/GAOumITjuOLcj80zq
qwLS+W5Nc3b4LsKTvX8k4ANLPL8dMnq86LfjtVhEseRXhxiVPAh+TCt5Pq47Vy5fzpgqXJxWkP1r
+qzScx4PrG1Edui3oThyUwvv2K1wV2N0W4vjrXfed+XUGGOdWKZYkTIsI1ViTpaZSE8ZlZrNzjJe
D2u2zKEYYwSt5yp6poRS5JgIM4phfiW94BFFxCIynxlveTaU3NZ5RR/yHscLvuyfocUFg6C5c5kz
GNWYRB1ycVHjwORgUK5+OqwCYA8h374762kEn74sSmmTIK08Dp4L91Tq8xPMMnKRxbwCFbWNcyvV
6NvwW+tWSP1K9mRYXwXIlR0zdNgPjz+XnXI1AwZkcAFHZzX4CV6fXnpePjILAIHxGG4rW9TtdHVQ
6yCYgSMbbWo2so6gvYEIdB/34xSy7WeBNNFcC6Vye45xkaPS1QgDz0M3W5HvOVyzNJ+Hus4HmxVb
/DxvvNR6LveNwUSKMadE55HMEk1GI21D4ARf+E2aKZyOkwoFPBbIcLOhABVYv1rVQaV6WmgBaVYd
rNbYB6vfE5dkr8DxFCrD+LxiM+rXubbLipNimMT7KmIy21QGkJyHFxbXgRGvFG4XOyOr/gayrqPF
p0XWsUhCwP4GkSgbTccUSYiDqZfU4g8PddFDAXvnTTgD/x/WAX3TVBKWimCKmYDg/+1y9zjL4cC1
TWuQ1GWaoV1S1GmNa9C0t7v2IVBbJQwI6FnbVZ2QSW2exHdG132nMPDOFOe/k4NH9WuVk3n7vu0S
8WYeosglBfYCBGmBWSvYbgNMoITDTB4jvFRu6QHoptRBKZ+zBfu8fk5tc/YpD7/dv8dUKe5giLcI
StUubNKiBiC2GoOnzBgKnXijW6bfN3QfKgCFu2DjRw8TL5rOaS8IXFQ34g/Y3bgFMo0TOp0On0s2
A+Ovf2IiM86FKSl83ZbfaEEA8mTwaEih7bt+OvnAaLtgfIwTiISWwgJGVaG5GeCSdV1IoG5IjyYr
Qedi9n4prsW+wx5iWc+ArByP5QHFwBFRBIr2gWg60KFD+CziVBVIz4FdWu6xQSUxk+sWZ4u4XcOW
cd8Pp4HKN0nyMdTOaw702VET+Zx4+OZljER0Rz3oB7DeqSuu5atOl6DriWdjxn/HZx3+V6KShcsY
igKA2DGPmwFiHuN0HyJUzBUkUcQV7J4K2hDN/khHNyN1SdlGiyOflxT9K4NgPrRyp7yF84ZeKOrB
tTHqZGfu4Tcepgv5M85clqewFYnxw4LEddNMTv8CjUfmv4pnfHktdzK2zBxEVVSW7a8LvomhOrGP
zQlzdHP+vrpOYyiC0m5PWhTNV7oWt5WodlsIfyWG6mZKq9wZYOT2OkSGUZZJQtRoynBek0xw6id/
bYeH86e+lLNd79G0TkeuXXiNjuou/LT9zoW2Oyf086uRAvTUauMRBmTnQkO5311AXRD9HZeVCcaM
w6pifl5LtvJ2ERN5A/yr6FqNG/3SiabEQv2pBpcJsI144sJkUhVY565XxluWuGBG27DXYp0Db1aF
MezvHWX8O5VYr1jirz4aW0WS/cOdbk1pCpmIaCqNHAFvDigIGZHubpdDH67DdfVHAhflinLj3Y4r
uwOthEsu6uiBQXH/+RL8w+wMEp4cmW0+Fpft7lsGL+6eqs+/iKUpbR76oAXt+iJYJ7Wj/StFX3tc
NPWixpGw5cNS4A0fb5jwNqd82COwJDJ068leGdi3pijvR5CN9XWBkngIWlcbmsZK315zV+NSGYyZ
Bkab31QkaDYkMxtn437NjGPXQic/n1jvMXBpCibiTg0lRp/n/vekRWAzUohDbk9/XLNgWaQzZR2F
ouSodkECBx0QinUuoRlzAvuAoInHLAhnS2AZkxwHYg3EIEKRiYaEgPidVZr8m/nhyqUZ0axYBQG3
6/O+de+Qb8oYoIWycfBVOKLTr8QUAhHr4pHeSpitkNBbWnINZEpACYaKBCsWjmSrHTIU+FTyvo53
9ZSuT1Ju7l/zbmaqbquEs8CLUiLg04C3zrmqtOtO9KwxavFLO8nBnKmibVwVszDTFwHow1eBXbiO
mxRgnZ43S96L75FLpOTKf2FGdTsxxdDd5XkdIQ3euN3AUoufq728JbDgfu2sbl6C+Z6nOknEN8in
RlUlS9vUK6zKhWa+S03tI7DguzsD5QzVL5up1do8tLStdz7z0cmPz8bi/Wt+fcnC3KsMAUPWnAu8
gzNJFw16vLFikgOtyy82bF+vlGNJyf6C4WYXJrBveMsDIYjvm0FemgTfYuzp2OKpR65qYtBq+BWh
n/M0EPyIFEIV0L/RF6JKCAUDl2Tf1Q5BG1XzuXDDF7epsS9PaaQWaqkbb7dIeog0+nw5ASaf/Kz9
Gh6L8f1NusQYIFtYxgYrT8x4NTv1wE/EP/PMbu8UTj9+PRq8Mi/q5ztuD1LAmzg5MuYrDttrbIsK
swPvsLxKyJt+VW6+SrUYKPSzhs7/z3sY7Sj49pLW5FpilmbYXh6iHqyAhwEvJv9WCQ0nXOUomnh5
FG1jkYbT3ZziH/VSl8RHatjiOsEqPtczXJbn0rzB4gEKcJLENVcVKx5raM7f+6i2h1H+sdqfDPTA
vDvTj2J981Wgc2GhbHbkg9NfjmpH8H6sciSDG7jDHKhsQhP0zmRx8A8WPMEeTzsfxyKv/LoiM63d
hhmUnv/TUrwbf2V0XeHphBg4oeLBDV5RbbvoyhCvMK8BbQ2Uga62gZ21u7X1elJzxsZqJFjUIZDP
ErYdaSiGrpYeoNsIqCqKbD6gUe4PzMcCuvOlmfEn8P+BD6FD+hcGCtHXbPcS9N21JiyWQ5DyHg5e
H3MMaMpoBgdRppp4Y2xfrWKGequxupUpYAjkhLw5SDR5L034GktwU63kkI0SoY/EpTVfh76XsiZi
BYImcMJRO5s3MijiTAB9gh+0zQA9gcSgT448hv/PVgA6dsHjwYi61SG+9GKr1PPDYYsQfA1ZejiB
0QI8t6HLsmLwoMvKcRhk7s03aIJzLhSPfinCzlSbAttmj8HLKy22upejtWddoS0WJDNo+7cooj6E
v5u9W3UG0HKA7oaNRMLJUmW0Wfgi6OQLQQ2PjnpDidhb7xw3aEa7Dhvx3Eo89wRtS2acT8dTJICQ
JrezW/EFszHfCLDwhmUSsRsL8uyT1fxWbNfbXh6F7dRJ3MogCYNp/nodbNZnyjie6qAZzAFmOBns
KPO76pdMmA0MjJOd4X4pPHNtnoVFotw+aMg9vNXm6+FyLAMdx1clWj4D6Lev2OASbmXeLlBFKt/F
Rfh6AogeqVGp8YAKqZ5Ub6IPBP0BvgBfRImmFaSGRdfJcWd7J/PsLl7HpYfRfWKm8ZtxgAVrIcsE
Q9aOEfFxUF3p2uNftptj0D3HNCemz+bEcsRgfTwIfQfc0aJoi0V1yrq1Rh67zinNkuOpB/FD4EiA
d/n2Hl5K79rMJUEtdD4g++QSX4SAZ2unB8EbOGKtcv7gOeNidbvfGxlSvpGczn5RBXtiBup9mPds
md2gkhOPEjTMfD740wtrqmJmDLrdBpwzF2rc0YNRlHiq40EFPZ/o+/FpIFgWIIouwr6FdtlQhvFy
DCQ9mtRNbRJpQIV37c+iwqqQePsCCY32fOKdKDDrQyPs5aKW3a48loKJy0aG0GYewfeGGbelfhDa
vuXjZzdTEBqkdnqDeY0E2jetvopoCMgPbAO0N7yperoDPk79lSINAsvJ+H4eW8V8etA8cX/dKkmG
LCvm7qVUL4D2XKIBpZmPyaAYlqUb0rqpc+GSYJQmA4VmuRCg/TcChjxSq+bm/KTg1W7z2rvwaZYv
QaI/qhjFYd4Ww9+7O6Jibykb1gKkL+vonszy83uPBWDSkA9SZJYqo73p5E9+JW2ijxdmrlgcoDOo
U54JcanYz9fp3nD3TTkMLkSbIpwv4jNSQorBx3F7E8lnohk1ZsIvPLGjBTTB813MbWPDICZroNzA
cEucx+hApOEDe7z+/UzDnXLuVZUQkoOCycSd+YWtVU/NtX05fu6JuI4rj6FAdld3nmAm9rgYALGn
OKGetXLAq1n3c3N7PbHq2pEzogZGS04r1F55ulsTF8dx6OISOf5cO1oYSbAleZMkiOgSlMg9Mqje
1mSDdXRKkeAieLDBjsXBPqozCQ9WUMqmAJumt2AxrNPXdSzS2ghPDq2Sb9kF7tDqaT0JqBP6pKxm
PswVMkPbBN+0Y+D1uTdr+bi88eLZLCdWWrSkuSSIkHsSC3dRA9SqQaRqoLMeaBSb1PKqRGXdVl29
t4I/TACvl5GuoLI/AsHa/fsL9iIrTAUrbVQ2E/ehN87Q78vGcT4z9uOIujrCq/Px0Tit3VzQMBwt
L6fZWz8JCYx4Cz7fLV3tRLmFZf5yz1PIoJIA8GalUgW2OXBq8HwMY73TATPqVKRb22w0q+5dgcjy
j3dHB8629NKhlQvZl8F06MyWFKkQQTDtiFbFsS7ioDGMqXgQQfisX9CDeVq7aetmfnRi6H0KhobF
I1J6DHyCI04p+xbXCs3an2HX3XYFJwHhTniTwSaCgEHF6EA3KHD0GYR3RIvcamnIU7pmEcRwxDz9
ZWhuNRAUpUdlwIH2z/TPwxF7ri/CE82uEDgHchFPqCHVzqs8/Fq7gAM+MjT72AOKcHlE76poXfL/
idK8WT4Vha2tsev+9jS5hV5hRpTQRF9EoTsC9IPZOK7IM4gjyKnmsUaXScFasMfPBfJrz1UuxZaO
spZtAFcY1AShtfpDqJr/xHFTCu834irdwr7Uystf/BdHHbNIAxXItis2kQYXsGMpMUgx+9BPo3mM
8E7ZOT/hovHO3lkmasC/8E0AYEcUPc5K4HE769yrubO9qcNBz447szcMjrNpCyZqzsx3M4rnBXXd
PFAqOLrZBYw7QOzjr4bAWmyEenbcRFcVLpg7/Wxa4/IfMyEXSuZhoihZQt0HcKgbltU2KAGIwoRx
kLP9yGFRHpflrEvZ0LZxgQaFi/G1H1JETiUK1mmGubJlcVpaNWPPnY86pWcpeChzjaLAtQIk0ffq
AC3ggkgeVS/9m/xl0r0q36vw16lpm8D9IdmhG7KsFXy20mOyGJIHkfiRP059QEL/YSb1CJBatbU2
UXAlTWsloxLlKCDpRS7nkGaxH420kL9CefyNidG4IS5VUuN0vGWD1iByOITgQRx/Bv6qw4d+b8qz
9Wct0dUPVv+wuwKROpjKcjl3LeLrN6Ud2KRBX1ZjSxX3cuGsHwzGUnXgF3JUgOFcrtQKjUEFqD8H
Q3Vc3hQY7vVm/JTZ62UGzTbxlfs84GkTGUaITqd2SgkcXQHxtEXGOrQ2sMKsC2ealZ1nw6L+8wdf
chmilRf1djJfDR7JnFyNkWR/uANHwKr7Shu0mTZclxeoLPlEdwloFnZtWDVqkpvro9an6Gf/XNj5
kVzTZYJabFKr/268UZZhejX8TSqnR648MBzfOdk853Nmz0ZHgA6hpf5GPAdOPwExngmsStINAhrc
cUB1x9bdzs4OV+Ev/HvXDPWHLBITxYjBpL47u31hK+99G11Ms9p6k7nUaxAQ0YXWCsQ6GrQRY8zt
IC1Lz2eqwttrTksPoQtw3RsCcxTIBHAF++3F+/82MwpNHnul27vO+0ZRt/7zzzbsQTH6+gvkXIX7
G9l+ySJlTrdn8X8UM2lEExze869vQen6jg33vNwCD8fNw/YNoeNWZ9WAM7J+OER4QFRLUvcyd0cB
Qel/AmXupg1dYf6aW+yiK2fopp/ybtQ03tgfvlL5nCFniXDKjFsM2IqSxK4arWzByMf4fdiqeZop
Ep7V+/mok31/Mr4QXnnLit4drfBFW1sHI9jMnW7WtVWN45rfYfClom2gEdwQ/Zw+XK5w9X3qA5q9
2aIHQOvZDjl2rURfeZ2Y1zeIv/or4VaMf/VnKDBMg2GqSB0x707s8X5TAxLfn9eHkN/DhxT5JlKe
3f3GrhtlY/B7cGbvvU0IyhaGmS8q+syBETjcbZyjEqoR/B3a7c1ZDJIMPN+Y+5oTeECeSPYMmRpc
hbEzb9z3QiPUCgvDboCBPez4Pil9CjjkBePAkPjHqrtGncjaHyf/CQ+mJioNd5yrHjaRXFGOJNk6
pLDcmhPRIf+KwBaWl8X/wTiSw/+Z6Jhd5fGrGYcNrQmXRGx4GqX8Si7TqMkKfLkpRyJZIBT2FeGm
wi8sylIDnr8Ucli7LnshPqDdkFkEcg5sM75P0k2ZunvIt1BVPkGe3YkeIcDqgFCEG9PC/itFuj5W
XBaV9giXfpuX7jbJJV4DW8uGIgTo3Mfg2sH9lK7FYM/z+7xXqsrqNEAXWoer6xJY7NNP1TNr0HpO
OCXZ3G6qC+AyzOLgc7eaFs57xupvaqs3pADUKzHa4CTTAHqI3cPVbKNNtxvxQdv5uGdjXVOKkBzW
hjO2r7Y5kvaQRMu9s4pXRrPGKw/2BLnTOwP+zbuibSv47s59a+m1zAb9oE79NaTayeA0uBVvQD55
Ei8PRPLlHhwUSdxcaiKnNbYpDqOlXRI8ekk41Zf0Uc7CFHGbk98ZlYu3SMp8mmoh9QjeOo5GfADH
+p6sYhEyVLYkZod9yKhMR7q8UkF737fcsByTHem05zN/m2Ajq6VpiRggi/Km4xuWq0IT8deRZDRU
0d0sKDBvNxnTNf+E44ZnJnfubTwChrzo+4RlQs15oCxXI/w4PFYHBnOwdioixxRxc0uVhar2z88N
H7H2HBa0sw74njsrTNs0OOyzZIBAxeycPxvGXAlbPZtaRuWGi1CUT45WKYIdVpTa2h/JlKAYIex4
QsDmSHEZKiDgm/6iYAH8BMjNq3dbcof5PgsyhBIhSbH5mVpvM89WAj3h0++Km1iHULY2XlcksPVG
PlcFLNBrMDn8H2KdVIbnn2SZJCxW+jjE1UBEZjZAPMwpfTeQvlUz8p+NKHpayWLJO5r1DonC70zT
O121QKc1abN76RBcUasV0oZOw6+0RPqHP44ZLvzQig/rhGhRb3rG3KcMz4VQxIQR15TX1CrY0txh
HGWW1AobVPlE++RPfIKmS/U/5M0AUsfM2sGwKKMEAayciZBgCujEEjhsVrgV+9gyzVqel523fg9k
sNSIeH/5zkV1kjrtiKWnKEnH1YtGTX8mVxUzyVpEHP7jQg05ebxmXXoC51mXIAQhpulDT0HNxRnU
mx5Mlk/dIq0WPYE4yjh8lXbfVhzH4L0sYl4Q3AcJO1yPfoxzMtfQsxdbRmThR3Ar6JeHh/Xogq1j
rue3C6Xx1+1v+mmjTGGR499eBCvgDURt+xQ2/6FlGHTh+/pchon8GK9c2cGjT6A/WtHrrJde3KH0
hCdnLTGR6FSEBWtNN0zeRgw2eYKzdSNJDu04V8Ybxv4udRnmS3zIU2/loaWzl6h7hteuu3i6v9Yi
9ge8CoGgPB1kdYYYJ+xw2eweN5nUmdWh2fjgLbOV6AOXIoeSBkMXhb0QNG+WniSgQBM/tC8+cwrF
n1GT+Sn3w0PoSYzgvrfvlSJTcXAB83PKoYVhgS2cin3y0MUhoVYZalvCVnBoB7PtHZ5VIYcu979D
Or03IGrMg3mddPGTiDEI0D9lmoJVWVAqkzpfHx5BE6asiiK77pR/fXJqQNAB1AA1/Ovzsjwnw19J
/0qIDXZNS042YQ7hBn/GAieaad1sOsE7uMX4pxndRIifkF8NIg57MEGNiRrBv4v4LB5r72zZlwA/
6m4X4hkc8+J2Qk/Uz+ikLlDC653YJEInRfGd62AdNFfwCB81QBWprEVX89Sh0EG+HgZKsdicrNxL
AMGXpdxVnjjNbP9FULSJtYVswNuQfTfD4sY62i3Zlgyaz62+M+8pTqIL7A9gbkjh9NzRZUAjWp8N
OxyZxhoOWOt45QOIDCh22bBTySy/ffvEgNw34p+mINCZLio9XtWB3wJ2RnFro6xr3oc5kQOb7Tif
XWfItChRR2UzqRD0MxqT6a8nGZoIZ2gSSMZR11eHrJRxQOQ10ePtaMcZNecGjHF1XoWQE4ob3C+E
VFISkdX1zujW5oxcb73ekEiQyPaon6u27DSb5yCmhr0XH3H+dEXMqw9GzUAOtKOeAWk/5Q4IiCs0
Qce1i1BOD83qJzDOrvTeLmhhSOgHOm4ZFa6+pPVvkGDaCWOm573zx5i2nyA7HiAsC6UXagLDxZG/
Igz2xkuVDw5+Cfz5GKIw065FkGQCZJZNnh1h0QkJ+gs4yPkA1KNZEFuDeJiI2lIe8jOaAGBe0YnP
mOhWew9lPTB3/nHkpAq4ZHQ8SxOxS3zZ+WUhP99K1dsu+JcPLxH5ddDu8/MJtPovqj5HtS5FIB2W
SZ2MR8Uhlr/bo3evgKb/HnT4meHXw0mvwF8KWCdSbUPhV6qSDCpDVCVbe6oghQCR6xcddjZ5+Xg+
CADo+v3eUTJ5A6RzK/7eKclL2ceLK6u612TufulaMpWzSPnxXfG/ke8v137sVo0q7qITzojz6ZR9
3stk39KPvfkb2e2jKb37DpKVH9D9w1WOHO8OIkItXclACoLOFoOoRY3AGztgAkR/r0AIJGb4ZTUU
p9L0iP/z8jeSUd7dbPA/8FzKEju6fPDT1Fw7SwC7Wi0uEHNWLzYIHUL5ammAu6gBrZmUWoIPqHkx
LznPYl5gdwGfJxc/dlxSVLYPO+ujDEq/C8C9F3sHXVAyB+nVGk3smTa0dpq489kBjutoRLm71CA3
tdjqGdl2btUKzz0sl53kk6jlasPmFohCjJDphflHHDwKNkXsbsM91iEEJu5MqxD2/x2zUiA4OqYx
z6GTT2yth1/u8MeAb/7P4g5qcfDeoX5btsQqEM2bzArncPwppjfg+fvwLy9vkNaNdqOr7p9JvPc8
B0eSi8/vyNc6yMMtJ24VqmB5zvb7xm14i8hXHf1jhu80/Qz/4ZYPwkujGy/EiGpGC8fv2mYJG/Iz
h9WxVcGRD33OarlrImtxnVX3xpwmPDh3kAM9yJ+YIBKtXDWelZCBbE2qBclJrNmIHUsXdalvBfMh
zoNma7EEJds/09ojyT3K/T1l0QhTFFYxO9ggLhGVWUw7osFYZei5savgHwFXAfSDzPxd+AbWKpaE
lS3xZSc6MMEcTaLJEapgXTKMwl9otqrNyCKV/Kg4MccUaffspe0CS31k+697utC/slhvYBZfXnax
xB/CEqA5/+NHyEVWTwFOR0vXPhXq+dLawx25LQ0pWwLk8BNevr3LoKdCLDybTm0P6bvLDyY7DttW
Yj18IiAL50lJeSaWdEBO/hs4DXAuXB0aQIR1j1kNKi5zwR+n40XljuhZdcDV6oUNJDLXlA2hmqiT
oHdR1Oqw2/iw1HBT04iJp/OGAfMRAHeOrmeVCtA7O6xF2A4CqYlk2Ux4yD/4Pst0QlRg311aLr0L
vrB4VTVQIqK5UZzpTM0WRzwc5GTD6ifhKD6KwFR6lgigqKixnUwE2o5esEogcvR55UiwGSbO+l+Y
5C/ouT8EJvUwXNQyY5lOLVmaiIH905NXbco6cvgPt3D02kDiQ/GP77KdZ8QjF80nL56zlxTk6BGH
nFXnbND4vDUVqw3GeCRsJ4wrJYY0yMK0eNO4BqAuBAocBuKUiI7tQ1aof6E3rtERa29T06bXu0B9
UVxxPpmFtcjc2cUC0xpHcO/zfyMKxmDIF5H0mg5jYzlXRH1ioBys2yvVHQJtMRY8fHRcofY41wr5
jcN5GsnguGiKURBfdq1gnQv98iOhHeA0R/YaiBqKLDXS9jHNWCVo0Vz9FpRlXY0EuomXmZk5/vWI
9ik9IdYzJo31kKXmdLonXjk9K5cQkskeejTU+tmzroldz4dJSm5rhdGJlt8M5I/e5yUQyvIjPapd
iwOV2II4gBQmUnQ91NjwqefYsM+Hc9mV+eVrSAvEzK5vsVQriRJ0YRb7q9S46fT7eHoQcB1a2XsH
2q5j3Iio7PeZ8W3qK3lmZ1IKrtV6mfRZaY7uKV3fmsfpo6i/D4Rah8tnlys7Ny50YLZmyIusN7+e
LFNxwlTDCioVVxwpm1ui8pM56cw1KTMrXolZncAFmf7r9lPIbDtWLEY8N5iFogx8TI6NU/+ZFMY9
AJ/IjSdZCDyF2iYQM30MJVo2xY6OMH+WYfmAJ3Jwj+gTZwiomqGp4W/4alTL8l1UOT+lp7kPj2xH
HBfaVSfNlunOOhlZ0Os4/aSIQzOZPa36cNg0Gra1p6jLXrba0pQB5GZO0zaf2ApyNfBLejoDsA7W
mwGLWCvCNfOApItQCCiOGLQq2CpzHzQcpws1zvZ77G/LpzMCSh9euXmZgpdgPY3juU8b+dN79sCp
tR5CqfzRb4Q7kbGwjqJ4jxz84+ug2PKpeNemx7EoDgyhFR2itXk2l2dhHi2hMq8BmtWCsqbyOX6E
BivGpCo/Q1XrmGJV5Ia1mNxGEAaTk0niVnI3cNKdjb3mtlKwvAj9pfcI/kROfazqTQEOyJHsY76m
5DsX9V411Kgkim7TczAquonvT1p67wEeEcOxxgCEQm286iWHFBStArMqNOrisR6g6KMVWK13EzkC
73AyLjhIifsEhBThxDXZcKcx0kTFQ1tIC7GgTJzO5AQcBqRrMFtKkrN6L7iiduVEXr3c7yr9lmeF
B9n4ktN7EYvSx4qG5R68HAyYoD+4G66nU9qmCS3yyqh/VnM4c7gza5VSh4Tss12gcvO2UKmFePYE
NAHC1IbaEEaUmk43KjVLJSbcjt15TE8kMemsKv2wxtx1rAB/vPjXHtcwKBDsV+WPqB4JvsZtvSeV
PeHpvR7h96TtjnVphFjzPnN+5+y/5kCnQjGMWLBTijVnnqiJDQ4fsqnGQFCdVswjW61wCz5nImfT
b/y6a1bX3Yoe740Y9k2XOydct34eV+T+e3zMWCpYcLFXklyipx9EGl+TlAh/TLTr97hpVlJCjubN
U4s36tFSBVSLzGELn8dPvlu6o2qvSiydZ3LH6apOh2AeahRc7gfRQK1MaiwKsdW5tidK2QVi+07e
LjlKVSKU5Cw9ydLm0qxyYckzYAy8JxD7odqIZq0a3bK/SiOyOzAozL4rV6wQ//oMDkiWcnbPPVii
ZWe3PgH2oMWwjFtbOYVNQv5FhaRhEyZyj624n/UVXSCC0RqJp58lzBE2OPQZO41beuvxLsOewoEs
sN5A6L1zte1qBrg5NfuX0+nUGcplJjmmKNfyH4j2bAAlBhazP1wcKnj9AgPvtYzPSAVKAgw4mqfQ
r99Hu83d2rwCijxntNFIxVTYcvk+2oiv/dmosfBZk6mdJBPmKSXZgHzG4ZNIG7Nq+9UPS6htTXfM
otc30GcQjyLSR/fkONg1Px4cJBMlp074O7YQTCerkszCUwbFxMrCbRJYw3+IrnCRr8twkIMjke0L
Zzg8brgf9MZU3K4zcoBBldlJstbXIhs+BSN+Wy/wURB02vn9b1psCkldxujQdOjVQ/24VIWSxJRd
Kw7jCrP+Y9wkm9gT/zJWSiviOYqka0ebmzjGvhlM1njVGsJNuuDWFE9398zOikF+2ct+XQIro4h3
Xg7R2nkDjfQ0XX+irAbwvTV0Mn2y81vIXo7DggAP52yxemn7ARJWxv12vqD0ptmhLbKGk9bKbAXF
K9J1ZA+PSCK70OFDxwFUFfvy+kpLhJXfVdSkQ46utFEKCGglkjz3hsvzZTQt4xS2r6nnYQgEiP+U
KfrnjsZvEMvJ4VSzdueirg/zTUfjHa/kN1s/JOMudjFMInGODcVSGqLLbppqrRMF9jfO/9DNCv4O
yICjI5kBkDjnczEGnaCMd04inGTuYEvxaqIWyGtNXr76YpHGhhOHcRZHTOAipWLg7/Z5mo/3HcSg
jjg8ed5UoK/RV3PB+Uawgy9DHckXPkkqSddcewxZIkpDUUy4fMopBd2Mm5GKV5I5lTd/8XxMEqKs
cD8/Bl6JDFJcdQsPma3bzkS+Ni2Ij296bgzLJHZyvAfCx8asrCFo6fAsFOjUPDWEgDd6CQUoFyVD
rwh2L8njykL2XrDZMZE1M255k55LbxlYSfQiqfuMsP6pcLR6CJDxQwsT10pa600MaBIUxiIycna8
4UseTvsj1fnqxrp/RHddxSI3SE+dFlDh/r9w9WAlk470dDWNXaO+emgkOocgRS0GTMplHUA1dN6Q
nAnPtHTdTEa3zmpayd68+FvzZr3VwfDMUBbQOhy4rQKIqhzL0Bd9vAqsgUk/IGC1rHarZZ3oxSBZ
3iUKypuFQj/0z62A8f6QhM557P/TZi24iVF2nwm0PucS17ncYlN6zoYMHWJT9duRWPv/mhThcTpw
It9WhFlkItdkta8wgPw2x6XsoOv4edZm5mopFE1utX0uq5YKOXxUlXCBoRrUe9/I6h4j/6eMJZAQ
Y9+8ko09n0s8Z4/MRjAt3T8R7/n6lFbg3zsj48WKGMKnii3BNjwEXFAswz2fsX/Wh0jgs8zIJRcQ
ywaIw6g4XkuX8kFJcoxgaUIIrTa5/iItwvZ5bZqOXe9p60j7/SgDMSW04x3nS4P2p8aLzIqfJ6Z1
SeiebkvRx0fCyrxxOrVYMQv794F8QT7DuJ4wYVp3pFvqmDI1mwUxGh4y/OmoiMuP6Fcdqr+cRG1r
tQBSO7UJHv3TGzMf4xZCONLh2xmq0LcF2ydT8gTxPZ2fhm9/v5v1ZqYfbJ5dzwXYvs3ND25Mwtnq
s5ylYTBM4dHHjZpuK9DqK4FvaNYacHU8+8JQ8+iM2Ja521jIPEUnf59qf0ZkcPTjXqelzU9bXG3k
rUIQEHMvNbrSCXYn4aCekszB8y0dRsLKmluhKuTBiU4G2IlIAjjqvYTJk/loQ/PBNn8sqn7tBVpW
N0FqQ/dx2fLpOv/UeSM++wzDuUmhghX5jm8CrFr1KuZoNQPWhw8er/6TQXU584NlqY2kN6JDSFod
jgYq86G8RWzJxXw6e/mHyMpw/u16csmhZIC91PpBVS5Qy8LoknyuHgjEDZsFo/E5bztxUuT2EcoW
lqkNUCgkHJYbhjD+y+y3/rRqgFF2bmdSQ2LNj7CD3vVF4cmo3L69RwrPVzxRtdAPLypim7viBHv7
6qa7O4SEdOHmy5uxj1zs4dldZt/AK7fOUjT9otGPAKM8h0DSF5FXh/dw2AuWkjZ2xN0PfwCZwwo5
NBHi6jQ0kabRY2SGy28po9e7EF8BvZOhhIns/7KTeSE6pwIAKPsXeARrzoHZbVogIW5VRMIkLNrO
NtCnq40hIbKOgt1ErS38giwHJ39Qxt4+FHUTukLASX0+jVN9N0HFppJowc5UY+JflBjUd1FmudBe
jA7pxgp73J5EyOMICO3ok0DbV4HnPsNFWOS1W9yarlKXrY0kwk0GHjGK5nFbFu7doP7aP5DcIAeg
sxEhlw7DGlHdCReRGOg81xJDDG1zZ7znu4tBLdL3A/PhWprPYHJwGySVHhdlYtCXL4NJEcCwaQ4E
M8wTmdQvx7OuaHDxpq8+p8lJdUkkN5g488bMxCVxUCHcdr2aU5WH3Ro7VTWLsT5LCSkbrZi1RwTD
lInZP2b1e/m/kz5ilAtZCJOfCudwUa1aeLar9gERCRRZ5n6v+r+5A3vvZ00fI3z3aRhGFPNF0GZp
/6utUKYR00tf8vkCnWG/kJqPMg3ewQM9pVtaL5G2HdnIQWOIOdaaRYv0JgbJDeuWx3GAi6U/e9GW
LTu6n0yyPR7agq5Im4yf6q2fpL64axr0pKLSo6gycZIx5FU0dvAAKnLW+wlH14erADuaOhHIcaOP
BX+CLxKr2Ypdz/GyBdaSTNyeJ2C0u9vJPVnDvm0xUBMFSf7RtSC6ypBGx6V+RM+nGDTXjB/zDhIT
atBxWDEz09YzJe1CxkQOXp1oK2F52DJ+pPEciFYlV4qgrCMd184/oaFK8lGUnJXIALsGXwdFG+tY
DiFGMQ0Do86qc7AjzDz7OrSg0lMo7vIR8C17bdmy4iCtFjzmY7rDpgA9bmGyRF7g+KJk51W4/YoH
k9g42gznj/F9uRsp6hO/ET8sU4ibs/Mb2vx+q5DAhrwV81Q5HkU3fjpL2qamX2HmCLCW7LPKTYfH
FVhxoPPax+DlcpGmwPKEWnz3rSqPd6HAsNaMThhqjQK9wAJFRBPQ1bYXQSn/aGZUk9+GusKihe6q
CpCFzXtqHJ+J//W5S5PJRi0IOvTHcAIjP5mdsdWpx/popasV1TfVfEZqo/Omm8NBOhl5z8WS1Gib
f4fr07StpRr6qZhyG03DugTcaw5fQ5kDj+FyeZKK+OjxrWhfz9/F1XwwlXo7NnnNsWHsyyasnZaS
HNk6AhPsRCNHchcllsYEhMStwXpTJHNeW4k+vjDvKbeNUOubcrxh9c2hLEUBQLVnBrGJHI70wa+G
f3n+KDs+vU8LwKSOz/gewAIOClKZLMe4Zkn12/JNfjE3NCQCjzPE/fqMYmxQToxDsTmT5U1l2mY3
hccVECzsqibTHw12E6qhhA/lRdGaFb3qcNbEmTLfERdf0SxYzeaY9l0hybq+wtOvAEShnEabbtlt
9tRRizuApKdx9omjQgwZ6CM6afgFKRbS7V3WUws3hZ8wVRdnj0NJCCcU2JMjT+srzq8UEH3WV3ww
C4kqVWMDjD+zuFXlhv47u17PRuTLGhHsOdYB+FEYpmEP6MjH13GRiFysh4a7xYGJbSRpB0wsDsZS
IgqIbXH8GukgO7RMsIfKVxxlN33BT+ZOEpsGwNuX+oMSL+gNp0v6wl776WigG+SKdN+FcZSs3XzM
27ltS37DH85VMb23xTrkbo1SDCCywF74vCyYsr3SIwHgRP+vpTQN5JGC7XC+CaDSrKpl6uWqHUd4
G2o9WrPsTB3ilgeUG+7B+w9URfdkt8p5pmuknvyQXT5DgYAF97tPO8xVkBhTWROpll7hdKaMuBRF
sF6XFCXR5SexMweyZ8dFRL7Do7lx9OXTOl7Bz5VnZDzCx2oPOos3i9W7AgTZwA6R4d+QMhMs2gWd
xdglmM+FHRonPwmXgqRhkU95/gOerxkG6JC6jB4y0E71gfw7nTeuLrm9TbKrHqbjHSdUe4yekg5s
MDGlv7Z1xVt6+LrGHKMQblKlgFGFm8G9VETN9SNYaNuP+l8qnLyphqnz1RpEt6FpKWqm18YU0zF0
S5mAFMxLc5M7k2+sMQTUNkdosDw+fRgkUPiVSRoncF1j75KKk49AmG0SduMRWOGXINSDznbnfemX
wvbcUxAcF2BN1qybBObuDlMWaaWUjOwvhNSLFDGPz7M6jTqJoW1gI7W8OVDqiu/ouTQKRbrDc8by
b75ObyLBO8w+YOZVJpYw986QPn4ypDnOc199C+HuAifTef87nu5qAfFceeXYlIpppOWPYDYfcIPm
iCTH+pvmKx9x44BYAHDInQQ7bsfCQoGA+4xvEq/kJJKgCtagCUjdr2IVNOcaomGf6NCrr/q5FISG
MwP/JAyjIRB1GFCMQRSvHtHJsdR1FED2NCt3L4CxheDT3KD7yFK9PjxJUdOMaURm6j3F3kAwmbf8
lso49H7mQRpj4APOoVF5+F5Lk2ay+4/jgDpm4az05JL8kuzvxMZLwcJ6y6SpV1cp24C9Da5D6pPX
/9xaM4MqlWobUPGweGl6dKo3cbESc8ifNzlYkTnQMVIhIEEJT8QOX6v0+COMj2Je26Zbjnt/PuDT
I6MnaTZVjludow73ZUQzT2gLIcJvSSL7igVw1oe8hqjQbJgS67EkbcBgjHHpUXk6XTGu788ChUhv
apVaYoSbigD62WwQdqmbI7lSOSggqYHv9uP41Jh9p5UKVMpXQ8LwNWr+LEZ/1WKqGyUTQhFCXeJq
lI+/ok0jY9TfUHaUQyK6mREAdIfwzxiqmnd2qbleNKd9v63G8+2sxXL/LdBE9Vte/8K3O6VcnpFd
ORvNV194etJBVt7+zMssLaGUTArYFSehgUfkLUL30kRJhCzsiDx0+AkV/wPFYeOecT/6xelISfDT
Adi2nsKg/cqgyMe/r8V5lxdVDDMC7X4hat/Dz4PgAa6OQGfOD8C8tnAhDuUy+xwJ9nTQRhfxMD26
OiP4saIWIdPR0P/SuPm1P06cUJt99Sk/myBuS/m9dmy4IYkTAN0QjtT4kFTD9mY/hZdMOzDCZWsE
rYA0nADVdcX65FjXj6QLyUUA/l2Tt5ccyMMEvJZVodyZWoEwtTWObsnNjI7+yj9nx1eZaYqwXCuK
HP1IIc9pomTUFlK154c7RIWhUtX6oeRhpaaNFPC1ccnSaB0uiA3YVlLdBjDRwk20Qma+6MFd1s/U
RlOPXzRQjUEGmDfKRXi6btG4RtcUDSO43oU7VAidBvn0y5LbT9qHNnR9CZhgDwBhnrqBQ0KYG8Su
aZCbAFliupkQXmwIsVTjxZA2wyDcAaHiCxmOWOjvMhemXC8epoZbsQvSIT0BPBGuzcWvTedAIHGq
5t9i6nv+L0NSTpw+aCbFu8JXo6JceacYTORjGpr8pFx17pBd4cPW7JLsA085xEL0/PlFYGX25JDJ
CS6lW89bGP7bpxgKq0E0Hw9kNaGZa3NZSLw2xmLMYrybtsF3xERHr3DVaDlzsmW+ntXGmIASaFEX
OkRI6GEf8/qT2TCm9oLKqelLL4DdvzzoF3iyASRad4audh7d9f6GauQWJFP4lS2iw4EA3w90lG+5
wfcwL8agIUw+v2CF+umM9ziNaHPGiHjskK9LZCJmdozRE2Kz4mDh/ijLsE4kRWgmZuvwWAA5eYDO
4IQemJdboRj08ihzelmQRZMmkDqbentJ7vuqlFTv+Ntpt3i82KYJMiTLJrpmjg3FPyzC3f+BfYDQ
b18keVaRsv5/uddoZoSViYs2mm6nfCpJDo2sFxMoLExsu58Z4rBEbXYgPLlqbcIfC83GPRqRG68O
w/R6KDSR1i9+W5GqKNT69AnwAPgGuwAAa3QrgF8mia85hWwCAfIcUYhpstG/fiNnl/N6epQh9k7C
H8npK4h+BagprfMy6Vp//8Nm6A266XqIJK1HT8dr5/5JFcS2bnLmqhLJ0rAp/UEGWrLCJs1BJ/+L
6i3lYJZyMGGhC2zjEIzWpaf+7MSXP5Y5HNdl+antJ0yjkitp15GEi7bUXIPHWh9pLsdayyhfaHId
hwtAiD8JoxHQunVlaTqt+fjmYjlLbBkcQYhi8TI0h/QYOMYuAiLO6HqTsNlNtqtqDduN6edRkYZP
Y6IFWAFR0vIu9RnuOntZnWllDRNWpiom/7Gb0NoLtEBHl33giOXZOM+jJHTaK21fym9qVtdC2Mm/
wlaKgEwUUiD1ZiFu0R5D+lSDBer0xs2uVXtjHQLcZWI3LdkRZbvVcRoJp/5442ts351vsjox9XRe
PLp+HASMAawqMaoRuuKN5wt8IkJ2RWjs3hDkMre/qdVLHSuQqoERP/dJFns2l7DrLKmsSH9MHqnT
kM7++GNc/zKZ05dpCbRfblaST1ijdlRlkyfFS9kx4k8i9WClJjl0a6RbYH1FH8BrWKEMWqIb0Z/2
pZ8EgHynFQq4GfF5Tw2fQcbJWKARFii7RyiIu8GYyfsujUiDsy1eadbcdVHHVnLc6QIgsAVMxqEb
KHHcJ0d/GUWtGzisFZk4u67L9pt7d4boHo4KXQ8diPP4dWZOrZzMzU9Gkzi300TxHrnkN1H9/OSp
4EGUKePnJ9aVsokNQsTAzTa0+jiIdH1J+6rZp2YICWDbJ2pXJXWM3ZXVq9LR2+Y0KnV9/71ksGzP
0fTfeisYPvkf0BFxzcFaaMtq0C/Vmwf6wqTfUYHouPWZnfmnP9uxgsz83PsdizLWAV1Jcfyp+hEj
2FtluLtWqcjLCSFLwpwHD4efrmqc+WW1WE6o50Q3+H9/KAyfv6UGardaX5/xB/3kRzUzg+i6afmF
5wwtrj5yZ4NURDblZNS4IkCa/McGnjX2CYcZGzioxF514ixAgRtasGtQ+HWR1z/KfEpfAIdfevHG
id1WVJri3GFIefAubGs7l5D4eyO5FHckTt5WkKHywoh6zMlSWVhX15Yfieu7ffPeyKMBwRIlYY9y
7eeqzcS/vFc0E61UxKCHc6+vBeVB7Mb+YiiZslqZDbN+pDOvnWLGpvGLZKY3jDxR16gqOStUewZ4
pCsH39WtcZzhSvnItVGHgKO3u3Auu+99ZS97D83ICgk7jcsIBbBSp6fiBV5GEYXHb4AoAfZPfIo2
Xch1WCUMfGhhtn5N1RSf2xqQaJbGrrO8bmI6CX6xuaxr2jUlH2HJlFEyyEQTZ0uUT978u5/SBiaR
jqn6i6Pd9COQVoAzm/63U09tZiAHcYy7PQ2I0ydaAJ0icpvgWpEcOSseoInRIaAWhtDsflfPB0Xw
8jizRwksf9da1JTNlRtiVuZx603Klsd2yQsTpkJmptsc1VDgR5elu6F2+S1eSBeGMiyvg94FLRcg
FWc7lBW0Iq6uRvl8I3T8GJ3KbgvlWMQ6dyuecvSsc8xSEjqHitfqBdwT5S1J0KrFrWdqGaF2Fpbb
008cC7jec3r5bpNH4ToTkUMyu4y1Us7no0MCx6Mxdu4nz6EhJvIRF+bF8cH4UuOHd/yrWfY0mXYQ
gaNItuHrxkTdVipBztEYtxWYsXBvK0+skyO4rMCW3oGV2iY6wmKfmnKBd7CbsS8nICATEGKHOsUc
sBZ3ZPGGOf5w4z6cvs2TgBgdCueNXjx67YkedD215efwS99Jb6LhCl3UqMaNTW8Xp87++NlZfBOZ
ote+a00maUWA6pWDGBWsdw+FtAgZq9WY0depd05XtdPnoeXo3XyQF6Eezbe03/koTYT3ew5WBojJ
vxh93FHs84DL47Ldn1HXnLx+EgHY+Y69SlyS5a3IMrVSyr4motKPQ2ByQsf198BEScv0gHqSZPWW
iCXniycVKUOqgvqfrJsFYcWXkYZIxrEapS3mLfEs4nc3fmgCvIWFuL+ceixui11FBYslML41msIm
R3i5SE8CfLWq7hphSxkJfhET0mZ7F6TZEat5fhxPOIoLFPiwAx3SUiHuFPM2odRLlruBg8k5jkeS
3VdFZH2g8aBo8dJn4UcrwMCqKDqTi9FabMO1SC/KR2gPp7OSNa6cD8G9Cq7SX825Qr5cLtm/JHTC
dPxIKHBWtuIGerL+4y9OWFrf2pJ3MSALdlk28JwAR9RAZYe27l+VATHThADNPO4IRSPhSLRKWFVC
8bx4SkN1z1tP4Esnf9Fw4eGgbt74mzk+Df6Hn+/36ufTo+6Kj8i1A5+L6nokvbk2YAdxIXh1X3FD
pr39dT0Y9N7bOC9qeBeWJdmqn8QrH14Cdq3pWGNmCQXOMaSfS8u9Vyldhidbgw8skNeOjO0LNIvf
Q9uM8nSoBgnStGfICSPHj5J0emtxqjyU6qdw6dWI1v/A9HLY/JOpr8i8z6hm2WkB7Orb/NhGlO2X
ZLD12ZRGeNXu/PxVjJTaFoUpUpHzShlCQQkSAlNCDa3MbQJ/VNy3q9fVli2Irk1jwfaQSPb4VzI7
Ie0CkFfcH38wkDJzsHpZ+AT9h9Gpgk9u6ViYawQ6S6D5gOBU5t3SlSxyDI96I9SynoZQrsBFddCe
0++WAXkQ1vaiRRySKCSEwDWdQUjG541USwcvkwx1Mf0vUuqSMgUhv6m7wKE3YMN35XE3JZtx2Wde
RR4XnUrXH/52SE0BewmuV+QPETE53zLVgvw5yKRvBpslj0COACbkpfn0CHp8lcSnO4nDLQCZEyLv
Ny7I8kgLJQBV1OGoVn3A3LXWEb3d6yLXTVLeRaOshBk05Oy6vmvqx7+fKwudd3X3kRHpYjyrp3ul
TXkVpPt+7mspkbSpdWgL1SoGVNNdpqArPbc4+HE8mZBEoj80kdfdrFvBhmzezT8/yM43cle+nNv5
CczsVB5WCAf6c/xUgVjdFhxUyjTX1KoU85eM+L9FwhPrejZ8G39fZWJRDVaG8GdfVG67Z6poysyt
xrdNIlatMenIf1hqzNOxkmVm3SlNSVpq9ij05rfjWPDQQ9WkIGQLBpdjZ/785zWy6tvC1PzREk9g
rkR/P3BAmgfJ9aWW8klcYPDqbWtdaUQ/zCHScV58kCzWxJHAXXAmx7yvWa8EqLKuMidsL5KZDC8u
d7mjul191G4dOFoBj4FJoOR+UEoZCQh0MANEMFqmG/2VyjHAtOoS9BkasGcN0YVLY/8gtVdPqxyD
hmURo/HNlrvU6ar2mHY5Uk9bC979+O5QmLGH28LLxC5IV32TA3wjvLOFYtlIc2jWlIW+8wwm3lZI
7jbNMX/3k0un6WrQ4h7WVlfR2FnWSOT+6NYbXE9zB7Fl9po+b/AZ3zzOHTzBTfIZo9UGA3CM2QX3
xiLJzzTIpg4E5cMB0NTVqedAienEMg7amSU7D0Mk2twgHkuEXdjclmu45iLaQZUzn6uYghTO23Xy
Qkrjt4A6LAN1tbnsMjPf/t7e3/ZWf4fFglBrtgqxQRZr6jzv8lKlJ9xQWut36E8LVQZ2ICqYAlli
QLDEHE9q9rbyArnVxHBcyCtSHLJUyRQqFxXnZh682RuyQPc0F00rFQ93JaAKFsTXu1Lur/wGDk3r
I78uXezHhaVayhxDlfmKCLWcZFLEbXMqwwMRVEHTnP5OWriLlRaGUWu3GUkZAGFm1Y4O3f7cQcsL
KKJqLbZHwN5ITS0QUyhwYB2ifQ5bj4PmV6xLwSrd3RhpmEuGlopzylk+k5eKNSlUWPKRaOYQrRJx
SuoKfoF51hBDjNDPh8vgi1KASJv+MkaaY71a6Q3PFMcLHuHO58cYPiGB0Tiw/nrhQPE+EtkAnATQ
cL8Zyg+EQoNGS1FCJuMy4RaoJREneSYlv5CAT0ArMhZlKeQ+nvlDZ5iPJ5yobXyWzSWCnCQ8hHfi
YR+x1p23m8PjfiAg9q0pxpuiZYTVnTv6vW9NOJ4T3rQyccYeFyQQhMQB5+qPRRgQWcH5BDPSA9V9
quWbQhO06t4XpcKLSC6WG80VtkAZnnELz5zXjoRcRLuFXF1ANffuwuVybdSxda9lhFW37yUyx88a
rUzFQgsrC0HurC6FSEv7PQAL5ppYOYK58yFrO/Kzftkk6mx0PowRZDz8p5xTN3vtmpu+4DJ95R9F
BuWtKE+ZcnnY7aVm30DDo1xpF8HUeDpN3WMayKrwlIhxVuL9nvwWfThKpiB9whbOfmmTq4Uk+kY4
HVDI2JiQztoHQUw7Ouincwo7vyPrVcKvcmFrPP78P8jNpV8weLkuAZD/BmyVjlIvbWd6LddZavoD
Z7SZDDaD4QVV+q12tKV2jWwEcV2XDteMNu1amIHfi2tZ7YzZV8t7XRbSzKBLsS8naVg/eB3L0XXo
3X0u5PB7TrSGXPwKYFrAssurVL4NXpzgRiQhPcfnh7mSsw8R8u9ZCaUjVEXMwrV74Qh+jXizCHGU
6ofBpcqV98OxB+ZHrGsSnnLYNbV7T2/pI3B5EKf09d0UsuIlnOWv3DWCWKXfbkmX82g5OqutueKd
5QaKrXQVXTCBvm2c8rMsbMr2S9jBUKTa42lOgIUfnwTiutP3w9UXqBLb747sCk/g1MdNrhuTeHnG
AQtmylANaZ+Q5K9ajLNchJ8BGIpth5vwyyZvTTctA8xTjqn7fjegEmryLrVOeljwlPzhp3LnFdOA
yK2Qe9qL9cE3krySKeM1zqsPYG6gIOnKHXFlIrKc2ip4L/itNj5czE+yexFADt2Iif9lV82D+fV9
xBv57sMtjeEwPSfOSeTL1q++v15zgvNyxC3uBA7WBs9n00WOJujFrHtnh3ZqZzUhILhyE/8dXfxX
tPiLbFwKtVqR6aSWOcvIl1RfqePyypZFAy1u3vTrTHWnu3s9Kdu1pOyzVmrLrjaKMUui0YfbU83Y
LY8P27g0u/GbUgwQDnWzJDrOnFn4rGaWtENMhrEH4KCzQt2juAh4hqlhl+8T4Pia/UKBmpKL2l+g
0l65L0z9MvbVNyWuHEMs9SrVj9tLXWg7oP6lCzhGRrehZR+wE85wlLLqmoSnPgt0k4IGMJcSAfzv
tVRcyN4x63b7qmY1C8L+0kcxxUfkqVReCuy5LIiuRHNjgc2OEDw9znAaQfuyVOI8rM4yql9wWzXJ
yZHhSmfwglLOHDRDHnpY8GuoR8YJd6lxBxwl8fFaH03IkhMO/pqq228BT626TBEMpOLsmUemlgOz
8ol2X80KtP8Ef5DHYp97VfbbLlDtml7K3zEAtjYpCF92I7JLjXIMYmXpkMZuX61KS5V2OdVgpaI1
duX6k/MaNnGdtZpU572K2C8j/F6ZP8MKPWiuqVdUzwl/1r1Z/aIp1RFTrOis90QgP4NvLSaY2EFw
gCm8QOf4XRiq/47GW4BaRCm9Pw9e8q/skFQsdeHROkfbYAj7xKGWFYO1fqk4nIAUV8ddFainU1c8
fQky8MiX0udLqQ8XyJmdHaxHcx9k6dyYzMOorhovF7sEltHsC2RvQuRiacoGBCdHTeWfEQzLo9ta
r98En5XLaUHMf1CteiOBA6PtbJhVOc1MCl0zCkAUApbG3KpzHRtVgDTImYWiGLgzzbnoTILCBrTd
eLcViwn/69pAriPTGBv6q5dxiwIA9FiqRL+Lo7K67heAqqZ/ts01swKIl6bEbc0DgWbPu9tz8qTa
PCjzHIChYvgGiBREtgLNj84VGk/4R8QkJ1TXi0mzC16ulhFl9X++Qj7V5KjT4hVxi3t+2gPxfMlJ
+8IjSbB8OQbC8A1Ii9AvWIXYOr7NRdLpQHbwZXc1UufSih5aT4NSj6ZHGCPWWshwAewaXJmeYt1f
HHfM4bOW2118G0bxddUYL8siKEnMlm5AlBwiy4SWBORSIdgTHel7dOeXdTwtVkg5znGn/IpFVYSA
H5POU1T7tGlpjS0OfRo2fUCAh9x9c+yMyckDPbHEBoCMdsiShnAReRoUc4H3VdwQLjJA8xh/L5FB
3yU5TNR/thVgZYd1JVGcbJgd9/mhj+OQXTKvE87mCLuue5eSJLiXugu4sKrxTvVdm+i9QzRNuuA7
ATjkzycGm4+AI/Se8oybGbyi4jpDywptfw0OZ7JPXvXseBo0HwK3lh1q+ZGzFRaE2R8FMPoN7nl9
oh9PvZp68DJFWEezRak/SMTJJXal+99A5cw4JB3BBDgzyzsz9ulD9HKZUOP9Dihvg7ggS5MBddvA
0IkYfUI95Rk9RMlcaWjUwH9P/riqenj9Ppme19WtGUFQ8wx52Zwg6+PeTSpJid56Tne2kCvI6UTc
3AGkmQkTyLoWpcuURwWsW6Pl13one77OYpcvfVfwcAHUycfTHp/315maT6aa8kLJUujzR1cNDjr2
3a6n2+jOYWGUi6hshOoH0uJODT6Vw4z/eEmI7aqsId//7M3abY6J8YnjMCzR+fJwJVRHMX4ivAw8
Nf24pMUkHYFdj67jNMxlz/uoyhCygDV5mN0YrrXZwjjpduRPyD+W5q3OBxjS/9EexbXAn4gdWNJH
fodD+SGKxmn+4aQt8HjUxoixBhDaw6/wW8DonMZmtxtdUzh0AOcY9brdfl0AR1xExKbeYzxO5VN+
jOUUrnNEOeZmbwqUVbWow/w6p2lW4sXeQJ0dk0OmeyBMnXl8945f/747iIgGA9lCSnfmqHA++P7K
V8k9IFqZutjBhDXRgeCbrpQTDRrcwQXRq5506fmF7dI23fqG51cZalOjZqwdCUVQRYeE3tGmQw3g
gRK88APZJnVyhfK7q9qKi4SV2jZCBUWGzGJpkUqhNjbJ4HGffYpmeVO9J/OQ4SZFAwVPFXfAtSjT
/cAirb52VUFpLS9DLzGIRM+MPUGpkAXTZXDy+zmfeElLdgQLciXioV0gjRcpzlz6F8ei2mdmiVbt
5B8xXC3Wa4up1iLET+puNa0SLnnzcnIR5UVXd5CaJYifdV3pKJo+CuaEwfK9rj2APqUdRAwLk5Hd
gmmd6bl8M/yDkMigNlH7GbTF2kEIiGr9VuqlFr1ChUsm/FXdLCt7g3Kne9rgW0TLdKUbsQ5NSoIH
JnF6K6kAJrkAW19LlS6tdNjXsu6WSlGJEO88WVWd0P0CY4QgAMFN3a7Kt647/es0lWb+oDZU70kM
hIn2FndD8Vqi2SCkwIZrZb3AfjW1aneBoe1j0IlQhlyWLVGbqSORnMBvfv/SQkViO+5SmMLQKIhK
q6H+i7WUWsygUr2N4NWsb0LJlOW3UYm5uh8Y/EZfYt62Po5J4rXdQplCrGmU23dJ2lhJPnVbm/Ei
OUo+nTDIxFz41//jVTwDOKnGgMz8lx+aNebUySmujmI/GNAJW0HWBlrrdcMTlSn7+Kmmu2NkKOzo
OWz/BGBO6/phXin3udBoHH2cIIHqVrvHMqIwuoG1JWqXPRfCxAbYElj+ppQbTG2B8gd3uoiG0pV0
b5Sjw4aBFJyTqFkenv2al29/VD2t/WtpDln1wwj1g6BjU0aWHQjSdfR1Z+DURWtHwNgFhi2dIfFO
tZNmQHGEILIcBnugdUoThjigMYV1KQfkMVwwBEmzH2eKIKWV8hc/LZgG6DiZY3FzoytLlGhdc0Lt
POx/tol+M02z7iyPXByxZRJlTsf6rSehkR8J178gd+jT+9y6f+7hrABVO0+ZKb2MVDfBNN6EhgSQ
t3r6aQd37C1Kfec/Y6BPUVqULFYR/Xa394rFB3y4xz2OKoTlbFexQoaJPXoDeie9jBpfC+nlR99v
0HJOJ+aWD7TM1mji+gweIeLJGniH5XSrGnKj0EdsiUVrBGzNV3+kX1HITzqx2071bMoWIcbLSzn4
/hV6eXroetKyoxsgcTfXI+pXUvrVS5H8n1RoQK6DlLGuon/i/WV2uCGnEDiDcx61xyr5qqeLEOwX
1g7ZAAsEMMk1ycC48lY4JxuvSR1zxgO81zoqf7D2Jpm4ME77p/AxUg6Q83VJlCqvL8jxdr8UIq/h
RTahER2rAmepFxRSPFKGGGyRr/QSIpY2Z+VM9PLZGsfhhTFdm3Ni4oCRmUpgyftQBh/iou35ulQO
e1reN0Sfdnn7mOUjIuv6RNSviNtV9LnO7FnkWlJK3TxEEKk1iLD9VI/uU4wbbXwEuflFq2PRHdDb
WcvOYXLAY+/JMqDDJVvi59vqxW67xZW4UEbsETlR6Zy0hZ9rlk63i7OIlJIAJTIxURBjWphOUy9Y
hWReWB9/vltbgPReZMve/vmhAoWgD4rztIKcsk5n9Us2YIaIJKgAejlTa3Ibb3ZIJtVAB7weleeR
tBzrk3TN1Mm1aItWOGMzV+0SEFixWKBwm+IVDYN/ANAF3UAM54I0L3jYZU14xcirIzt8bLiZno0r
5AM+L940J6tcGWXGLMyB81rOAUwEW0EdcZjqYIWTTiu+2guxXmJWG4a8SW9psNNV3QnJMAbYmI+o
vJKfd6KxgSUWAoBP3vLnHkaOjjU6hRCnsqmtaex710psDHJryfKcjqfMErxF00xT8+kbucPR9lKm
rIXHHYp3fDUuoLx+EGqIrnu2pRHqwIdBl79wGmQcVGNwsrv8j2WR14Jy7VWFjwWJvME1qBmPHXcl
p/+NNnZcD1JlVIjyVPWrjyYMq8KciV/ffxpDy7nbtZFciyFzchgIoDg0A50VzPtiFtQuFutlv+5V
gVp190pNV5E7zf0aW1zvP8w5QXXXZ+DJIUpDfuISQDjVOmngNuyAh9OLNFroy+/kBm5N1OInXGm/
LP5apWwPqIFa/hebtOaFAwtcxf4WKCjxXljPScNCaAm1OzAl8GNGsGAqAEdKdMnDJN77ubsh+/b7
cYhigIWfFl5paEImz2gvRIBtLXHSfufpii8XtSRsehfFYCuoMr+2ZmJ6cfcFdsOGOdatxpW+qrBo
DZBlia0fqUftcpiumOqGNvPd5CKpFkLj95RvZ4AD+d+M8U5CMpvzYRw5+go3UJeqqalv2M2L3xtU
cYTLmZ7EQVNrfWd2ud1KD0DrX9fk0m3a2gdtK98nn1e2OzPnVvg30MfO6BIDHMG+Rr5mlaMqtC0j
Cpei/cOt/hIouwyJy54LKW+d8UzlOg4djdW0thz6g1pBHAR4zlEPIF7ByeYOztDAxwPk7BBATv82
TINPyE2sRbXhYcGJdUvRu42RillLJgUI4S//bgBGE6HkRWZ8KDk/F3dsU5sE4+LHULwM0AoEo1JC
G04X08trsdOTD5bWr20kBCWVPHTkk6Fe80VCJ5qRNJqo243B7pm5JHjXKCtB41Qx7tLBn+u+zdAt
hLH61M++4HtOiXaBEHy+sIhgq3jBHpq4FvK1XwTVOq8j9q3c8KatNO0j3BMeSEyMHsdTyK7QYCRh
5JYis9eRG0cpE28GnfSeLumye47w8VN6oUkYlSgr49ulF0n4Y+W1j6GwDUjXaPfVwRlsRjX4dLA8
8hw+iUocuTkbMLiLPCflkDlRiluhzeFH2djZHLZVGo1u0jaVyyNPVB7/OhPTqVWjLv3+BxU7PvS5
5oce/9x9TfOqGao9S4TtHFKqTPO6MPwTGnijvhYo4EUBsw3PAiCVVwMngkb8i8lsB2nGEIFN9J83
gx2Kjp46qAoQXKGfKNDdzefb+R9F/zdaJpJ5Dqc6K4T9epOzOBuh/nI31taJcSmyFPk8PnTaIZrm
WT56PeixJTh0bhxLImf4B7DvNQkFkwMJTIsmhW0UvRd5kPkl+u72J+Id2HLe/StCZs88TMN9+fAQ
N82w2ggMoWJNTBByjJvRbw2QhVulp72mNCqIhjiWDexGepBgd0Ha9IpyVh4zG100wv2/ng8vbwTH
v8t2SABTbF9lFnFmabFYZ7pq5jNDpufRBQkDkztjficGZlCY5E6pJsJ6uX5X0dtDxOJSc/mBjW+p
axkMSbhGlZMI+z0kBqlIQ30HHK1exilN+e3xNfj1E1F+65rK3TVHlvzbcenGDOGhqxlmR5jzlbxH
nYBuEyEIdmjVnxJZgBaVRU03rsBDGxx0ZW/xc6HyzTn5qnoWrAsuH77PgDDYGH7ipl5ZJL0c5Wi6
c5fE56r0XTTCrAFnt2p2oNmM+EX+piI8/zEDBJZwuJSjTAdB3uWq2wbZOnhElc6jV+bxB5Am3WC2
vdk5m4QFcu23PSYCK/OPzulpLyzJqYsJveawGb8Zbj5YXsXbWKXmyuySVeMnYECaOe89+e9WzpGp
0XP/dIwXktdiFEnFQ/rCGtoKnsFonDVuU8JIdsc5yHSHQF8SWlCRBDlwVo89DkXY6XcK2iDhxP5G
yuDoiYb5LC30rAPpELalZi2rYSPetrVIaKBXEE3K7YHGsql81cW7cjOYoTtgOzdz3hu9BCuiJsZy
zngbGjMyBpWqK6/4GMGHMeuDawK/l+AalKRCnfHuRAJ/ev7rs8Xk/uca1SiIAW1ZJ9t7nwtNNLeW
A8GeiA2OeXB7c0SEPBDIT/EmCyHpJt1NW8draPG7t4GjGYaBNhVCHHwMVNijMre+PHPERrcZ0Dcm
l9N6Y6ePYmoxfkEk4d8DfvP9Wozt3xxQAdqDOEogWHTRz5364LRMI5RN9/gCUDh4b3vv9EwAc1g5
Zqt4BiGJfuQ6TzsCkeJLGtL8z2eY8WKJp/BLyQyxh8JE53KyiK/gyTr9X9qjTMU6exJReW0YceFl
DYExYwBoiDa5XZE3Qo4wWsVD6QPUOtrUfOEAMNcjfmJ0pc+5G7hRlzhsC62OslsIxW3029opoGRr
6Gj4QDYAT71aywPzzgv5wyMp/XZ8CwfFxwTutLQFMDIOauVmSsodsEwy/w+TC3MGZvI/v4CT0aAQ
5ce6IoSrHNCOrZLblSjx7BtRneEB7ZQTmFDHITkfIG1C0zsgCbF8PhsYBSIhdZ0rniDp90Mb5krS
clAfeJI69wLTdscCogVQNCz8sdw6gexQgIKtzi9rSvQQzJprc0GM02jN12wq7EzFRQuLCa4Sv6vp
vGfGiAAoxjR9qoKN5RyB7r/pKb9b7Jpwxsa23O4mfQKIvk0sT6rk4Y7uTfa6kioejVzcQDW0EWGP
qUmsU6HkLuRMFfMxSCy6Gl/iYedrU6k7gAllv9xNFK4ghpKIAZgAP70o9f7aOX4+flZO+UPUTeoB
bDYJCVsfuBJ36pHcteMx6mEEepK0aUAT4CY+b5Y4HpEw5dtUnH/oZwPp4BXePEGTlf23k/6WLD38
Q61Z4NZ2WGsWtS+3tPS2DLdOQFQZIiC8JxcoholVafs/GlODQy+2sWGfJqmyfEqM6otlsYeVTRm5
6zvjSNTK89BgQHtIYNcega2iopGVXLwmqfnGIh4Na7wgRh1KZXc4RMFpJ+q0tIQj+BMvxo8lTY30
8S1NcHJsx3Yk/MWs1FfbrHY+A/YmPKiSOCtwrDWLIUy4liJ/olwbfKP48uqBZIYWVaUn45HUW21O
xKdX/SPnUtSTiN+kPV2kRcu/5yiGtnTQK84ZPsXpPhC+faZFAu5D5/BXEoBhcex0fXOM9xMeB2Un
dTJsN/t86rPkRPCgIMvOTA7y5//JIF2yybYovYjl36PS9gswuNrGlp7MeUhGLfSIwZ57dAJhgKqR
AHDEVQJqi/ZzCRdfxZern6B/RW7/KyVYcg7XZYBzMWBM9HEKIVeuj35cMj+wku+e2w/oN4HerQPU
i1su9wlKMejOMgvDRH3BoaQVC3PVj3wr8YX/3SXHqp+9Swp+P/Soc7tFClCb14HnzNW/ZqfiofOa
eVXUZbhxgA9YSgO6Zxob3SIjNqeUEYYcMM9BJY1DUVcqmOBGezuRy2H7g79OvLI/SesV73S+voVw
tug9c4HWKSnhp13NIY/oOs/oJuYr9cnGUqRah/MExzgE4QJmAT2ea8sFIeB4r50gOztXuBhG9Kbr
ELXYFpyiYmSIGoa+GVwxReMjQqscherpqaDad4KidtCrpyvEZr9aeLzdhzk6RCWZ5PefEwDLMFo0
U3n5n1qiMnwt9409RpzvCsOpG1YBFr6/gmvPCZTKqngWprHFBjm5Aww4UBfs3bE3xB7ZBcM5yaGu
SmQ4QUFGuFW7ts2sZWzIzOzfd8Ws3plxRME8390ekxI6pwVm7Y/wst/0JnMogmi94KzBxzEnJTnF
EH1za29SEcGalk+nD0RkR3RguhShedcBk9mGQz+8RI0mEWdwbqOIzgmnsK6zFDX9q4mufWXeiHNm
b5bQMSCgQMPBTA/rw1E1fCmuR8i6Fnst8NvWUlhpBC9nY57HEKzkqtJAxcOsnySVOm+08Ou0kxCk
4RQQQadrl1aTUwPJnBjEGx39LNqwVshQ8fbH//+zu+I9RCndZ++3c81dq5uh+OpP9Jvonpd+S1m+
bj9LBijdxdHMTQSkhdc1odyKF62tfgk2N+eXKws1SXmndwA60jk9umM9oBr8soFaLzLI1Q1KAvSI
vHcFA6X7yxrTrV5m3Pe7ZhfVW+cJpX5D9m8hR4aFhzF85ww/jNoY2lpQYsejjfcNZYWH5tyB18hn
Irmy9aOI5Gs4ZDupMqpOnUayT2bEs/12fLEAM7IRhmdbZYOvr70hLyRM6X5+NIXXzhhLaEDSA1BU
fFwqT4vGlHBHj5n03iesFpETMMOEOjxuKc1ukEvjSE5Fjzp4O8KVLQ7Ho9Bf9mWBgMvg8te6KD0n
BwUKulIbkSV0ODAWipx3d1Z3eDamVDakpkkH8H7x0HeHejDpd7VjTSyt4iqJ2hL/1IQ+QNYSYRUG
H9uPQbZrRBmK7pVBLMXDS3X/XAJZCOdkbIY55/GLqHmJ4266DDgzQn8Fmb9GCYOpXUGBcUWtFlB3
WDHdTK080c/TjGX9zaKlD4ehrUPGIui434Thu/qLz8F55DAJVcmmTMPGqG9QuHDGNY99qcQybLli
tJXimaYkLI5AQn5E0++UqeHewxnSXhZhY36TTL6XKNjPcxNFY54D9cnVIs3n27jMmIzbRq134XTQ
gwFAfeds4Z8sGICIyaG1BK+SKPPmsJXVx6NzIe5CJ0aV11DMRq0apTE1fdGEGcSSHx1VYd53xyCG
SyaUyv7N86tWKyhhbkyLTfEMuyen+ULQ1RIw9KYRdiwVYJPYgPs+PmzKU5HsI+3+XTN8I+91mjCW
c7HImOOkfdTqGD1GVudfOOk7jJcwOv0InLq9H1Df/dGcLfR+rRr2S4Riadk08uAoVKRvJ+SpzLk1
X5bXgJaJYRyldPmdQlwzbm4KZJW8WoaIhaT2yfn+mObq+pbly7YfmkTSkyE7j0E2SrWDPxHg9zfM
aTIQ6Acz/Cyirx6f17ZunSfG72Tn6cSs+baAMrT9lKfUN5XxyOCf2OP8evO32JCOAt+XeJQjxBMA
/dKXBzwU83PxnA2keeZdlbgb+hUpsx8TdaFBahxECFI+GDv5rcUH0J5o0pgtY0zkC5JRA5oqPCl4
6HroJcq2M+WeEbxln9ayHZiWtD/za6lQJ+stS/MeIZaiTSh6HLS5TI9dcA4qO65tLzG3KCawCK3j
/1His7mMaJ3qffCRKO4XAsQ7jcl8NM0/1jYvc1kupS9yXqGL2IvdVDfen3IjAg2+H26LTy8hVras
UwjZ5MWhjKZbj0ZYQEyHdSVpt3FLmcBI0wMS8Y72SnC/V2TlTulBtHEEtT5oh2KPEbVg8lmG3t90
FsI2o8kf1ct+NdeaoohO93NUf7dP/WYt4N/BaPnHWXN1i4LLqBIA5vXTZFhO3D1BSRntar+26gof
E1i9Qi04XVUfUdGMGVDlOThw1fq4g8KJ90n8X8kDnLlFAS68KIYofU4EU/06fggvRcno6R/rwJYr
8VZyXh09leaW95D9Of4pWeqgEMdp4jCmu0jjNKJi5YvUjwJZNXAr//HKL+rcT3qqBw1h1+QsGgqB
rHhpdD+FKA30M43pkBjZ6hgDhqTD/qQDM7JtyNKMrrqBfFxYOahXRNsPJeDZ+Neg/w3xwPdKU4Um
zGRbDsIlUFOdeGpMfaT+ROKZAP0UYqcbZeikJZ4Us5c7mLNUnPwx3QHwJ+yYnkkAgtKg8tDX120c
1vE4hEbwcrCcuyRPsS3BOpjMIm0kHJx6pKty55JOn0opCxRWLJwyU6TkN3o+b7daUDfaHFLQ8o+G
ASEcV+0G69rMroq1GzccpPxEdXDqJXbPRKxL2cpr7eLqPPgp582+MaAAJ0goF7vicTARBLLFkMpu
LKdIzw+PBOFVm7gkM4e5E5nO1LqXvW7p2ek9EtcpQGz87WCNuzpPxiHKa28kqgGfb+QgT3M+IFfE
a74UtmtETFqxbhilaZzaDjpznBurmCp9LL/SGuzWDFXhYYatqaH62IeKklU+XmecqBQ1FdHfgX3/
fAY/y6maKqXZOTWXg5fx/gdRE6Bf0vA5/iUW5z5YborWBZGEcMU1x2ihSbeIYcB+jd+oE+tViJiz
Ti6ISKHA4a+I36SM8NyaMEn3ePBZM5X6EV1SYfgTo1BS8A3f+a5ra2LK6grnJq2/uPlP9nX6k2vK
1eAbVdec5jRAfUPdVBfnAcOzngYYHnKx/zy9FuGberLH9e89pi5ooOy6yluqI8XXi+JLdV88gfAr
JI2hXbmu28Pm3FPd1u7s7Phq9rKI/WfVm3MZQRJSZD09MsynkHRqJuxjxcls8hBnUQT7zy0bFZu5
ps1YBA1d7jEI6hmNBfxrixevKQ53nmqnfwFHWenFOWpQ7xTZQJVL7JStJ6w1rTT26Lw4sAHogAzI
GUZ4NacUq25i1VQgCzvovbAhRpbn97nmYk9aeXtt05ksq5/+0naXB3LLSvlRSCtY0IuRSqF6xSi7
2MlzXyqya1ICOOT9YDekAiOpFL6+1uvtFzgL6pfA5Yve64REw/thuUg1QkdoXL1oMeTohdLhWF2u
l4wWm0/WKlVKgeLDsfeSvbf/5h4LErOBFU1RScGE6ev3JxInfx8YFk0mI48HrcMnRJ7OnPX9jk7D
JtnYUbZ7E1kmsF95/nacM39T5ZnQOsxrdOvG8pB9KSNDcWkmsvVvXEq3d5JhKHZju0Vh+aJhGvuq
4s9CWluKRootPAvRX9BEGgDIDA/nry6nYzK1p60CNL+uLB+HjPdQePk262ilyEjM5Xat4libUisq
UjCceMv2YL8c1RZCwdV04T7kS/2jStE21z1fyey08wAUVu54dRd9YNyZdE1XSvzgxAyqhgsmr0o0
jw79B/o1mX0WHW1Ok+FSrWRVcAZI1NRzfWIWG96MnFRPIGrPpKddENK21xlw+YmjAWpsMV/9Vn1H
9cwojZIKUgBvCUpsP0WVQX2DIejde1MnM6/a+NIb+WNpQYDUZkv1wUlYj4y280ufKRCVA9NSfVqc
sEM/TSf4YXqP557+yLINrrjPt8ZshvomMDy3OPsdfbQsK/OumBzjponMWEvyhYob9SjTNtAu29TB
cikqobLH0ss44LBeHtiiTV+55FPZMp6QOSn6SSYps530Jn0dMcu6Zn/DUqMg57ynGJMIRFopZfHY
i5/qICOWMCYGKpl59ut8/IBd+mvaEMPODwPXgZw0WY8dp1kJFkJjnd+DU0AcYYBLJhRnfbsftIGx
8b/zYRUpcKeDFSZJPYyRJbI3mU6NBuCosnWPIre5KTQwNOiu+W9ODmH77aoEP3eWitsJ4s+lvjgT
rh6K7YbB8Q7Mt5rYiUAYwMGiymdju1DUDDA1RK3BGC5Ym44SGHOglje925jz5BwAH8sBM+4de401
FAfu9+NjwHOyLAwMTMBFFROdn9PH0Svl13huT4/GqWDJiIYEMRniSFZC7mZRr2hInlaPCj1ZidGd
YMZISADKNdIW9At1vXh2uQaH7TqBWA7H9b9gdGFepzSwqhS4K3IwwnZP3rsJReKqpOJQdQ2EdL9Z
ZxlBhPSpsPLKsSvaK5CTJcVoYp2x0FG/UlhBUU61VQ4sB+/EesIiD3ZUHHF2htuzrTatjVtJib1L
APLc7BylTuolnvLBJVOc3zjXgZLiA6/RT3qCi98QWq74u4+7bz6GPBoTHbUkDQXDq200rJgT/uCJ
DhGPXFFtvJpIB1gyEPa6ScE/qbeVwPqpOmSkn+8vjgJ2noE+vEbbRCBRVIr0cZSDNFcyiaLccKGS
UrZaJ4KbWBENBQ4M3NumrrlKFShYF79xlaiB8G/ruzykcyqRVgiplsSIhy2KC6zNrhaQ+x5VvGDk
qxe8P7+JvGRiUrcTDKTA1+gsYMJF+d3GUcf1lkM/I1XAs6TGeOnxVQe2cGomcxNyEhQvUTMtlJWP
MY2AmxMljGmYK1bC1NsM5rqLd4TWIZ5SsXVmJ/mqyFMSFdNl/XSQzt/c7dEgO7hSIbcTdcc42Sp7
OFqEfRPzF1mwegMNDOWHyf4qOsK5RwBVjqQlnETzMJcjtv6C1/k6pHSAPWsjXHkKITxAQJDtv8Sz
kMvc4VrY5wqoUUA4zz2U9lIWPR6i1NkGoJnw6fftHF+xePER0iCCVLkN0h1KeT96Q6IIAnJ8oA3N
CpDwnSBJRe7UhrS2ZFfoxXL94QgTMtm5HtCgprtc4NoIXVur/ZovGYsd7BE0dlkaAjLsh9QnMzbI
zA8EKEwF+EP3DeXzUj1Jm5V9f0psx0WWCTIV62PABmTPG0nlcnKR5Z2c90xP7Y0ZStcUYRSqNqUb
Jq3kGM5Xc7Y5zfZonCjLFFshIetbKEODcoh5+Yiq2OnETiUR2GVoPq0GP7FM/N1YQ2M4teWm035b
ksqYOBcxAJpIOFwPOB8KZ+EAf2r3DUk35WXgicve6IjtIcJW1Bmkh8U7wep1dVFXLDKCubcX4XSy
OSykCVnghJ7Mc+LtzubruwXcfhe52hOIloImyZ7I0kyp/InIoD09T5hL6D/rvnb+Cq6uu+jdXtkd
KFGXqTA4EQODgwEgYHHyLQnXJteGraW3T8WSOYzpv+4vX30bsKE5wwvnX6s0NJvtPaLhhjfx+r06
HHWY5ccViBWFhK3y1HuaiG4M7IlVFbV7AV4ki2DdOAwcC/Rkb+U/FrxRK8/nKriCC4quYc1shacR
/pMkF2TogcoRaGBBoPbvM+/753l4ikNEQoVdYnvYmNDfqaCeQIONaqazNjGi+hQT0TH6Am0HyKzd
rAh7oGXFyHnYxVB2hs1qj7e3hbCl9o8nS8b9xBbKzC359z9gaVSijxDzGxdrz1+pT2FjdRHEWt7j
XTTJztAVSyGd6/2PvnRd8QbnRbl6UY8pg9dH5294B3dxUTMxMa/O8x9x50VIQuYqvmrMGTduFAHX
UUUDKnwwo22jzf6eJfm4/KN8SMx/zvUrRPWbDtXOR/m2YSH/z2rd8sLHLwbDzOxM1cwkuIR6sDFQ
D5z8hP6SXlSCCzwfknSE0cwBwkl4vw4qzCohpcynjWx3EEnF9v4rdjOj6KItdYGHl43f3pYHk8Cz
eeml8HKSU+0uPdw39ocZhZMIjQcX4j47LZ+/D+Ys6yf+yWBnB2stj/zbX9spe4P/wxc+R3ILgKtO
mv79SE4CYtuVILcjXrH8v2qJckQaL7I5PpjvTkAmJOq0R+LAtYuaOKxFlQXm2U2CKjGZ8xbsFSFj
O+UjeDl8s0tSn0KpRDRBjUgLvKVgIbULqKulZ9qeyBrTQuqw32sqyMOoLXZmlNNPKyWKQWddE54x
2P32ke3/gSmtDDNtsrcBr6qGW5Jj8QH0o9K7O99Cktrp7AYh0b8VLJM9A0GSias10pEr1Av27rI+
WwfbkGKAUxiB/JDqhU5jEr8FMet6Y1fynVN3FzaVNKV2bK2pIdZJQwyf1V1hai3kkAKSMurrNO/X
tRvrZ4oxCfUeIj5FZsJMkCHMAEHexIwk4gc/jMXQRSTjqXp5DGiCPgOdVVtiCltxmvkzCQq17JDa
eD0QJyF6vH1HkcAlj810C3IZWIkl9HHjiDx1Sw0/xji1dptCiZKyJUIwfFZyMjyhIyafkLGfX6ci
CGZwa4nuHEhWEMLTMSy062A8Vwlud/EA9AsGi4LGGfT+BoTst3kzkBHGHL2qvox/wa3hNdy89kfS
XE/0GwAL9C3OO4LSM+7geb+0JOeG9wbsK84e2Jp5YUFV1tfXmpNqYfvOZpYBYp1j5cB5gX2P7K9T
N2Ygj1XujQIYqo1TQ/zUZ6on7WLpKKj1GiN6QfP00q9/2z+hLew2wdobWZPDG1a+MdRoIUgTc2iC
UH5BCk+lf8hPtNdepzDDmvkOYnC/uThL+krU9YwVKrw92fnh5qmgesVxNRjeSrHNknt1Nep40SOb
NPiuhKV6M1CJjgPkOh9lA37UEVwb/SdyuepRyZDiwT+xLfrDgjIXBgZdj9sEnF/pSxonAaEwcfPq
p3ZRzWAvc09zJWpR/58Mxhd04Y3TA1mj5bl9bv9PAut6oJ6Ab2QKXQnSNajzCR7RfEZZXaBOx3ye
2dGE/mfR5p/Wc+vqx0wvbwvyK6e33cQueEjyOWGIyE9WOYH09CQcSpMnwAiPCcW3FGFnLINdG3pd
PmEKdgcKAUpm3w+WFIWa+cvQerO2IbwIrLh2lTaFnNZQqzjINmvObzjsws682hZJz9JoA2Cl3CY5
TXDDbLKt1KNh7yp2poi/Y90lwho+dp7sJ9XjKj4X/Ls7GCdonDyQfZjUQmsI59y7TmNqlyPya5uG
LurL6D6L5CBp09xNgKtCmaSuHDiv5kcR8MwJqFLl/xflNzFkQbZBu56zKZiBFaSN3nuoO8YIclhV
G4s2fLjVO1Pu6EjiTL2T1kuTeU6ZAB0OKRii8quZuiRSikHkbDXC8CcPlmf1veWZkQzVIV4Pi1jn
eVLKxSvP3hEFvS62mjZRFO1l7PadY6jbliEFhD0/5Y1Bxn8RVeW4YPvkw0TNE9w0pFeVk55OEeUv
n8ING4XPAdyswqhKSJM7BeZnU+Dxs10/oZpsbTM1ngv3bqO08G37REn5XliaqVj6o0EoAwu9t8sY
AeWgCR/XiebASGSTVzJoMWuebNsakdGnsTLk5a+LNi2owANeM2424GN5+GJ0aO8A8RtA4coNHQlM
No44oByoVRf+rjZE9v+hovvKAmOQLU57WnVsaiVq0Ze5UNnugZ0SOWTy+itzPcYHhL1VhpM1HBG8
660MGszsSzj1utthyWpk+KPeLE27D3VnnLHFOxcmq/osFd28+FnZIOlhAMrLIx0No0LKCnVssZ5T
FIuWqZv0d7FVdPODUqnoiA2l1Y0DZUBQngxPhw+sKEprQVgemBBmhsj9qfli56Qj/gCfuFoFG9Hx
ZUcTq7U8De0ZvEjVbOc2EotgLoDEBER62lixi1u31XNvfAIgmVfyeoIXI/10jp0Pw1ZC9yaBAU71
v8TifWTX/aVtiURUmXTRbnJ/X+qi7EmiqlRdHPXKnpokjycTJ0giJTgoOUShcGyzCTLrxaH9eg1C
OSoxlOigTDRv9xWB/4kTqq/tDd4E2sg/c4X3mld5+hoNVlcRW2A2PzyLNdEebivfEsbvccoOLd6p
CpSUJR1Lk19+ebwKf23v9slAQ4edbl5KA8TF1kTbBPYuS6NUur+vsm2zB51ofDocsCHuPsC9IrCw
xAB8crxS0teoxysELtd9z4w8yJj9kX+K40AGkgVHQoHpZwlcOJY/NS02FXFq9zWVTfZU2hC8vhv/
XnDmCF86gMvdW8fVbbHKk+AoxivDX+OESRF/+eQX2DsrFkwJeqI+xlv6OInMDB6XOOzOlZsn5RYm
N8WcwrXFdxiAImVVPpG37mRXo8FBAzfqNQAtGDYJeP7m9xLRb3PMB9dKoSyxObrrO0+lTCQNTlUm
Sw9kBRi24WhSCD2fXpfg+ivE3FLWXGcp0FwCJKOggmsy8hiLaMXax5i4lAmqKVRxFS0woQcf0yop
lomPqjJDOSccQe6mami1NreHgJMFr2v7OB72MZx2ukft92RSHtVWc0N/lKm8sA24c3ZHLhMc2tfZ
1Qa3SmsqB2gmAHanN+qgLu0QE0kepD0DsLMHP9k7L0Lfr71IHoKbJlqdodtIvXr4MXYgobzTcLLY
K5MUyGKPnS4HAPndS5l/BU3m0m8JOW4V8Cmr9KSjEpZR/7CIpZ5FTlB08BLipfJoSm+kaPya1iet
Tsk3cqDClLSgf6HoewKzNqoLZ/sPvSZOfKL8iEu+CQmDWeVE5nNxkk24nFtr1+8U7CkA8a8xsnkl
4+D4gmgVsoK0CTf/ciSkCfMojdkcn7rCHRHQQdEcKEh4UUM3x+LoHwKsWMk445PE5yv/tw+mgODr
Hsnr7a0dYRb1UjiT33Q9qE7wLpf0lkv6KW2Svs2FOIJnyo3QnnN+Tu7gX7xu3km1zqLVaVHXhADs
EEjSNOq10TqguKlwXeWiNI4f3d5G66Ze5YIC4mu3SMFXRrKdwVbTt+jUYNWO6UVQkyPBe3lCnT99
pDMuSICk6j9dfWA+tPSdVh1WuyJJsggaHcUXbO3QyZyhaeZE9uQfnlvYwHURCcrryZDJT9QwSeRy
t6zLiE5XGpv9C54/fGLl3Px3K8elfeRxtXGGHMikhTEurXe1n1CBsCkntMGhnsaheOTIpRPqf5o7
sAwZMvdRvek5SoIh8qzJ7Toiq7pnguntvvAdQQvTh3FxqTFwwaqrYysWE8rirnWQtIY92NBs0Y5p
6JaEz3mLHvg8SBisjA1pi4Usf4C0ibsG7HSacktnHa7MZUX5Um7W7cKqRkwhPIN5QxbGptx2j+5f
ouS/HVECqWLrCcGQ/1nMAzDoK0y7OG6eT2Xh15A5VPGLSboBO31uWjn4nwKX0dJXVX8aDn59nApc
IMWyhfjV5OMzoG3V0yC9B3NIfDJcfHVqZ+StFGsafrZ9sC3HKSc0miJahpJCyIuujuHccOI9nE9f
GUIL95d0yvb57DescW8LH+bCLQquN46fqM6MaOPOnh3FHiig1WMk/JGAbGtDtQe2KOoFcvq0pws4
89bLkI60GjVf6XE9xSowLesgu6PqiR3EI326oh3/C0acrEeL9hxI7WbemjGWKYC1jJogUZE8Nr/a
C2wfd3ND8QORthB2031L9TcjZkV3ihlU8Mq2z9Xa6DPP63QTl8wbFxwEhqExeXkzY2ZC18vEy0t2
6oI9HQsBnOfanhYrERgrbv/b9vHCHYIqFCaxlCu8jJJBXymKjtUpcL6XmyVMXRwU34hoQB3r+Tum
dqnkEl3MQLS2+GOvhHDR9fNoBdw5UffSb8OOw1FFPutVwFQaqkAiANSrF2lHdr8svlEyiDObqOp2
Wl/aJNuFZojrMvDA9isHCCZAm2918Q6ZJ6QyWuQWh2zGzZ3bWH3wQoo5nnkd5sJna1U6qqdQwR1K
PiUIpFDc/OUAz+u7FlM8wbA86S2oX845k+k0CWxveRmUEOD00sl8GMypTCqrIHwfB2JMaq/SbBXs
RrQfkD7oT7UZ25i9aa2e/Cxk1NXawb1V0VXOifak9c9tZWtzTvAEiZTDecF12gwSRC0VwdjsiBIc
WLRqWH1xyf+kFf/450MLRhUbh9zHHN8T8G6TLiYkfhf+A9T2CDOG9laDsNjd3w1HSTX2/1/YJzhB
BO3jaGSjJeIDeH/aHuy80X+vemwwag1KztHs8kkyuNY8Z7c6vhfiYM0abG+OvD35eCmaLTr5L6c9
yHCBgy5ikp3Iao5m55C7UZmpeDRT4NHpfQTQrJVmYyyPrIcWr+3o+IZUJuEkgkEzjihDMvpjvkwo
vNeg2RFkHrICLR5dX5FjG94sFa4wNOSNT1bg4rBqYG3vCQH+QgdCulgMkOxXCU/skPETwmjAW7UU
gGu7hUjJIEMM/mPSwVwyWeSlqrg/LDVL9cE7PNrSUwnC8/DbVMIdl/BSijDV7vLlQWVal+nJ151t
pruQkrPkAjx4MazcRLxOKXxzGKlikNy+ufO7po9ZOINtbQBNMAFcLJn/tbuOjeKrJB4JB4q8Tl6G
bV7RgZoZ+LpD/Ma8J3F+0Ol4DaQpsax96acPA4Pmy/ofwKKWPIKjfND3holH3S9Wh90LeiQAIRcA
pgdy3X13vrvRJLMZqbqoB3tGeu8bzEFyzyIVDCaUAtNrnls6yXoEs1PML+CeGyfG5aunhy45LEsl
DBs7Lz0dtOO0aECbguin92ltXq684X8zTWIerCh2Q9eY3+cBFBgEvXm8LVHf6kzm/BgKYjpHHOdY
4fR68q+uvT0n7X5d+ZVlhEhIOuT3EPikXQQu50g1Tfv9Dk6XOPqMYwzUQPlh9XP0ZtFb1L8Q+jI9
JU6WxuK5E9r9Q08+spTu2Q3Rs006hAnL7mNgWhnl8KeFG5O5xMfYrh2ZeJfmjVV7OjO6DgFOGkBN
sifPXpDqj6GWQpk+yn95Dat3Hbxmk140+6Dli6qdsnek5nbh7UTBSqtTLTw8CACpeVfQFnTcB2uI
wB3H7D+cnRj8u47e6THIelrId/cgLy7k6NiL335lPbIZCGa9JTS2It4k9M4QC0sVf0C9hlctv/fE
YT3j1f3XTNEN1xZiep4bJ1FA4IeQ2dkonJHLKXyJm/lM5Kfd++tj6F3r5qPDdVhnS1kvhITR+GyI
OEKUNZEWyrdcBQYUP3x51n3+qaJDDlX5BbxAHCsP6jQxg3ULCvqOxUw/JijJiVKZiOET4/IsC4X0
l8+dbomF0XU4Gb02AD1Rd2/zU+RwqhiIBeKdD0WO+pjmNDvzWfCXS8vm2JvqQU29osNS0+HE1fKm
g7BrddnHPiLL17gDsHX8jirh4VAg84wzLX44IJu7ilcjxBfa1FlpoYZDN9qWWtWxO7AgAknJj+t3
AI9SmGZ1sRU3Dm6/IjStSrPTMaPMx6Bi3rWwxek/VtFp4AXMXz6Jem7Nm9UmrFaiOoK3AxA0pX40
8IfJnngg6CgwtsmdLq9hWIvNBmBv29YyQG+KX/G90+i48L9Cs7wjV4hcEQRv+EtZpdZwMW4iJjgp
w9hQ4XY4ubTQsi2DW3XT8aQk7OoXRTLGXVFweX6GT7BTZPRq3GdPCY9/jdlMCIftSjMYVRInOx+i
RifXW7PrUKg2Nk0CZqfZUnc028LQj3rwjL4zj/xrR2B1++HmjSvc1g8fi+zwuj/uYhp9bZe5JQlv
HQgpKIBII80yKZ1R1Ry3UeTMLgm4ZVHr/tAMORnJ659wd7gtythUsw0e+I36lCGXz8XM7FXFlayM
uTyZDex9pmbySCKu047ZbYtrS1EKAX374hZE8YZfbNV+irHBTo6rRDsgUkqKfVE0/wVVRA2Cwd6G
9QSX5Hv4egQuwDmXXEW9Le2VhPF9RcRg/scsLYobzFsAZhauOLre7hY//WVvXRuYUuR3PCn9Q35f
ClEhV62bQZUPaq/lbKVKBqMA8VxerLTGh1CDByXCgZ9Js8BVDKb5PEgGAcM79Q0Z6vvG5sIrT9Pv
GMfzTNxxMb2MbLy9IPaSoQy8lgrnmTP+GgmBfHOJHnsS8WXUBIqyTzTTapvMuRP9klH95zyA/l8c
6bDps3P6etvGnPcsuv60lWht5yqkYTuZEHNP/gT7vtFdZtEAqBoMeEOK4zGXTo8rSmfs2++PdkSh
LUQXc86doJCQaIb9dU+CWNBNHlgdfEUqeo9gp1AhDKnGgIKuH5DXTwtPxTlHZrJg7GV/WHyvv7wy
3lSaDwp2H7nK0LxdZyCczD1wuYp/ZDaqeHXgkyZKFSDIAWV1WsOmtiTAggP3iSmInJQw5kkv9T8u
rtINdYH5GAeoyT5ZPyqfo/s1iF2CgoCrWAw5IQdQ66Z0T0gRstlz6NKzs7kl5i4CdDvA6QrQVyQZ
twuaJpzeqmNUftV/xGCkeAtNYWR6qfX1HLpo6bOy6XfPQVMeLz97jsz7YGSQoSVjSHx+iz+T9aVd
/60xezrUoGrXonutXNtwE3nUNetzAcWqmQ4wFhLsGd03Ol1Hw6TQYd/8PTpQYM2tjNEEl9Hq8oNA
6ZD1AGR2H6iPPqGi0h9+ztCgfqJ7JVfCP8WnkmLqK4EKvo/AoFj4lnRutM/OEpSQgIX0/mF8hIqv
E5dNHemlpVkzEt8G45GowOxyIkT+IGv5xuDRmlIqNwmJi9BFWfTAKaLIBiU0TwQnPEUIwqJr8QYx
TEYuRw7bQtkMHlhJxpl95MoTWCpctLgmHAPl+2luczJ6MhP3/fOO/yajPY79SynoDUzBQgt+7xhd
WEnsaZgxtKdkmj79mfJOINxY3lI6iKzpdZDq23qFOMeh+Oo041q954rpSMGLAfHow240MHneXVpI
v84CqbLOODcwSGkObr/LZTBOv5mLMCO2Q7BvFk8V7Ho0DXUuv1MsNWljmxOqbfy4E0zA5PMdKKH4
LT4jyxjVSGzOSBivAckdKpr220JsQ2iT6Zh6GFp/aDALluseW5Xy+iXjz9aJlx/WBUNT5uoimvFx
NXzoWudoKeHIGNQR+/VvW7E+kHVGnwssuNVjYlvKQnWycg18MI5Lm2gXNfCRYyEPJ22jbLxP2Ekw
DdQ9SMRbdM3UbbGtljRiZTgy3NYwEo08hNXnF4ykiS9Mir7KCcThradkaBmNw6wDHz3505ak4anA
o+bFHHlRfby6SyJ3J1+l9RbcOzIHgtW2254rw6PH7DXtF67elwX955D3ex6jiD8IzKrt0GMd7M6k
1o5Mb+NH1Ex23YzVSW3/FOwAGRVpVDSso1YN//QUpgq5G1It4sOJzHZugoWwmHURwrZoH11l7hTD
2SWapDd1JkKdXH/GF+Kxuto/9Oqe0rjjRRMewcpNnKZBfDFQuNM9ltvIX9m9WSztxNhkOg9EAeVh
Rc2JmoioazZYwfGp5fjdELlQU+n1IvJ4i0OHcVmX9GfaBVTl6z70pF69SZSRdvjKCJPSzJlC8Oes
t2CSi8Wh5ITRSK26CuCE1Bhz/X8v4L/oi1UXQ1Y/2HN/QuYINiAHbQo1ZnoyJM10EtiQMp//ZXDl
Z46CUJ4za7NWf9EPsDpHVJwz0X5357nmetILeRZJhIpVBWeeoQYpMxwkOjoQocWjRb7USBi2Da0k
dL1aBV+do+S7FlZ9DlssoLaE7loAwE/eVIyvYEq+LwG/z5NOVRBMfDtPY49xJf8hyK7j6IXEvWJ/
kkcv56loAlfzgCr7Ey39pw6F81ntBzs/Dh3RhaYm8/+keuC4hxCvmlEy15gft7eRqiuqS1uesyuq
tuBd/wZyAmcpvYQGzxHjxqeXBgSOlXX9xAVg5ec3fbJd5h2QhLu3n42wqehu7ieDH6DIFE74hUqh
yY8P8zCV9JcwqwCzj4+pD/V3NEOpovP+/3KmaCj9U6xFC7hKXWxs1ISHCUM50JEwfRMyk22Ka0QQ
bQvaWSpnlrej87xqGEEPDMMEPoV5+plzsoA0ptXSjcyQFQqASPaUlL5oC7LpaTA4DkRT33vYsnbn
zZVYTE7cibPoLTfNKABE4gg60DrdBtzZAlJdHRMz2ZwGjUL81RvT0Sg2tkodNT38S02OU9npRgTl
LIKj2TYv23FDwWag47X4qhsgdXvP2gfcbjxQqGTZ0ufmeGxETTKeJFvZXxgNBVVtR8dfk4/iewCp
BXjWeF9kMQEZH7/wMH4fR5YO36cKPjNAbCO7Ct+hg3QyK1VLW3qbtMyPx6UbJcfxzoG53K1P9ul7
4heDV/O+4skGwMR+hUyDy4yq31OawXYpJRGWd30/GGOJBEGPzGlHEjoDedMplOHdUYuLFNfaPw/K
4tISGQCstf78eyHBze4dFoaV9/VrETaJZxZrX98QpO8ZmWjPfzaY7bbWVP8nbqp4L5Yg2o8+AHAT
UVIm0MMRSc/9zmo3T/5DP6Q5A+37yvg66ezDuLe8YU7+KoFzX0QC4GjkNeQrNwVmOByUvjj5+GgC
cXqosLBKbgvqQrwRNjzZFkVMD5pVgySzDTaiiwApyH8aRaAffQPTQvitHiMnjhegmg7BT3qZwamm
iIvpySI29rDIy070stkBtSvdrfeien63EpiLyMqpd2AkfKH7TgD+IlVlWPaKhiDh//7nrhirCdJz
zJ1DMcGp6R+TpZeFyovTy2Jisg97Mb86ZJSOhIF5AEvb/lBUdqgPFYVi9HZT6Aj+9esNwbUd3t9t
XeAu2hs5AZM9o6N4wbUa5QG0ODh+8/xSctklDSdHSgJJQiZ5bliBUFU5pSyTVLeXDERAXigITBXp
nXqpZAL+4ROIbQvVexrE9VTqmcU3cF0b0UslXXGJdm/s8O7hA/nJWPhb/hz3FRwhB+yOgSDODK/3
6zdjxpvVJOauu/wkA0W7ECXSOixDWT5rLvM+FtIuBo+VWSpdewrEaLywVkuRqTGGeveRfYuFZfXr
02fk3L474m62F3jpX8ostjYOTDSV+EmUd6WfrBqJXqH8d5RwXziGKKPZxvzBLvu3r69uUghnJEqU
ZvEgzmqaSCviYNIZ0VfGa4AJuUhUjbuI5K6UzXFdKNv58bq9kOB39gc3a5Hg42WNYErZXNJ2Em3f
G36JmMRmL30EV44wniYEQJBpDf0kdMUAnuy4d/y6gTTUDWMVLNbhSmwo2A4Ag4W1iiavUnWVq5xj
ox+V8Ip8FF+FPdxnEZXRmV5elNoG9fhP9UIXa6iwW5cZglpzEVh3wYYXS0zglvg1j8YTcdV3ZNE8
qC04r06MC1sFDxntj8dzWlPfx9/H8cn5R03tsbXPwajIaj6UPebG6p8aL7tVZ/qPJDAe/pwcM/yF
do323k3TIgi3XxHbM74igMOJBj3rVZdTOtDkWZQEFxIavE90n9yPruQT0zs2/LPrWFfQUSvS2xIL
WendP1D93lDMYqfqnjgm3wkRo2pGlpaj1538NzswgeKAgHPMemhJPsBxYhOyb/8fz6Xrma/CT1FS
JwdVGQcxCsnJsAyHb4kAAAGEtdLvXNdj3kvv/VDJto4J20XoGJ2E9Bs8HHf2CgF6jtcv9NuIe51N
C47KvIycZEo1vQTBqUzcMTDRDy87pz29v7RnjkS6zl+7fskscYmWfRlruAqIvNvfjUi9iYIycwUg
IzClUmZN9GVusuoPLP+JvWNnMKOzvdfu/VYTUDT1JcC99qAf8SWJMl5Bv7zxfqKSqFZCRb380Tgn
Ox+V5WycLWnF2fJ5teeJgGQzm8UgdYVtWll2uA6DQZ1ZEiSyTIn3BqeNds+846hwinq0oOo5wZ6f
tVcs2c4yPRPdrN/mDLP8XrHBK/oJEpB7e6/R4NCvw0gfGnYTinQEXlUfb3MPAvE4jS7zYSaSHZsM
r/usftOEksoCkPgMMBrn73dY/wzCrzoY8+L3TA2THUjkE40AOvkVSIMYKDFlzN+NVi9hdv9NFJcM
v3MmCPyK0ubBThtsjPY2b/j0lwVljS2UKnDMspQNqp4uZuK+iGyqKMdhuB8fGhKsh8ZNse7auE2e
lMi524R9n0dSagBGaX+021yTiBuonXaRhhXKnN4ckxcJu28STCBUo7AH+H81hphvpJgsSZIx0sFq
Fz3i2bikUDDkc3XPjjX6eobAoRPGG1guzodLcq6FqtwvvAMfbbZI91j82GGoxdTPTz4AnlYDWKva
5KFtTvzWYi+V1SoX7zDslQawwLVCQpvhmrunXbAoJeYsSrvuK2kJUPJXnKbJIFYRZ2biAc2fYV6p
cy/bnJKMu+rM/8mPizzK67qL2sRynB/39zEorvHXurIxY9Ugnnme0FRovkhNLd7GI8ajpeVcWbqr
CN8UjOgfHAbG4R9bOfWtrwhTFRmp8cs29wNPkedY8uFRViV/BcmSR8pNeNAC58n27zJ2oJd4ayMc
gvaxFQDXNItAA9XdPdrPIE7mXbITvwwwv8TcLpjgrTSPs2IxeR3rv1Mcud2dhw9sgFdWwMB7ftZN
zgOyzTHIjy3LukHioyB+s24452SAkSEf0aO5F8cj+bVKkTNGvNeOqQuuX8dq/04ueHtOXVP+sqUR
7JHaEtHoZlX9cjoEZMUPAG/WgVaPENzPCYgcT90ms7Pfh4cUHfd1TJTlw6UmH4cpL39Od3gqVbRV
ORD2ucgIa1IABTxTEIesjWQdPtbU0ADwuiqMpWYzA60RPS6Nw5emqWQj5Cizmn3NQyyY5ehsKQzR
ZRJdhJlCHRkKPLa8rU8j8E4BrTIP0TgSo2Byr68oR8Hp8ovojYqkmtAupVx56PW7u8A2jq6+X474
fO+ABHOtTxrvNGYCsZ45fP/7IvLiNMw84pwcy+uqA1rv1KxJa/MenUEU6rD6Ffzm3Wr5qjwufPJG
TeCQFBOMJt33WO1LFqd1qOa4Qdye2NOAQUTiw6V6UZOqScx0+muClABu1O7dkBb+6dAA4qHFRuws
DmF74c98rdFdfSskAVm9SsSvEoHnjsvWtlK47CglAfbaGHpJ+3TZ2tVoC5UR6phF9bf0lvjIKE03
rul9JiQOgbWdNoHmcZxXfFH4+zCXuKoObJeCIyrNwtDljvmXJbCctAGkNroKoPRWOEm4JnjlvtH4
dCeArzBiPVjgirxbazWhwUxsonfkH+Cc/r1XXON/JtO6hwFggldka+Bu8e8mOaVUUNZwOvcJqSjS
StWTW7eYAM7P9oTMnzmqWGSJ9W05KgPYL1mtaoh7ADdmLSjdWI+qwMH37ejAYVq1l3NgDtgKTBJR
hj5g66+PKJxtYr9txrHup6QLNlQdoISwPjZfwEyIphEWJJ1r1HP1tnLnvkBuhmHqMnFJjZc/wUuN
uRV+weENpt39CBmQqa9e5v6pXSEE4xKr4wF64Xqw3s6G6zadTdUuUXtPyKjb4Crf+426CRAPUtq4
nFlKcC2Ecs4K3GVL6xRRpilb3pgtsxqaAx63HXWhkSDJy9W40qYfyv0LrNwb+eKRc2VN8/SeMaNm
RmTY2ZlcxlKyaX0PNCYa/f6MMSIOhFBz4PIeEYw08UtUhAQ9nDa3jV6HC1ra2aD3g2jhyL8eUeHK
mvw1YRExH3Diioe+hsZGmfr7zzOanNZrnpIl0i3k7eM1I9DCaTds9wKCEr6xqWDUGvGNq1cenerG
GmXhK+J0CVHfMWs2oxTqAY0Hf/d+T9lqIB24AWk4w9nNvv3yYXsfes4PE7DwOSDya/US2nYvwcv2
b7KVTtdu87/LIQrSexFBZZq86gkyYPXuC6Va9OV7HYhMD+fXTnS8dPVvU+r/yL4r79iP0IasfZTv
3nMfjnilNPnk0LLuR3xPF5QqnNE6S7vnVysJiSy6kOPs9aEmXzT5WbiVbFpGR1hVfLfqqKSArWaX
M84sQAGAM5382YGZBw1nFw4FSZjHJqrTesLsEeFtyvr+wiPw0Ss/uZtVeBuMbAhLkFRmX9F5rrIl
D2zDij9Mcl8Br7KTsoUfEkyZoaVyAogmEMJmcRRyBvHcEJ1SyNZz5sNNVlp3ElHnfti6b5uqyjIM
6SZZDzRvHw/yHbwhjmXykqdoLYXCk9wLunzuroQ990fkbrYdHcKsezpnjHqSCBlEpBTDCvEQybel
YJqZOo+fRHLU93R+i+dM/LTgIxquoSh6nc4xiUT+iKI0b+ZGRh8nJ44nDDtzQHhXjmGuEf7MZmHA
q7kaOzGifTfbXbo5Jp1lZnjlm8FS2JmRjmMLz71hpNwFkLVvPW6zlVPQkLnDzUdHsbH9R2VxBHf9
abwKpqldxlmELxHohk21KR55ZTTPdSkVHEo2s8kMYonST6EslIlRIQ0lecxAhOXuM+otWn0NbBpS
FEvYAhGfTFYPbkv6Eff1uF9865rOAhg63Cq0VnOFKrh5VI9M7lbMw0STbySGADVxUfHPOwR1aIwj
4gN0iwq5prlwuuX+dWc6+QU0ukRhRxBPYLGfG21jwjHtJ2yEPu3KcMi9h7uee2Zs3hMLLT2OvPoN
LFdzAhPEYhEWf1qcSuIcdOXtXz5ufJvVCfkARIzTU62XmI3DP1BQ1ZRzTWsbkJctWSPWAVbfWQxv
wpQt49y2fEo8nXPITMKtN1C18U8FLM8NXi0JloQlKw4lbzOFZhINysj4hDa7UVU5p1U+Xi3P1d7x
DB2nVbhiZR4WSlqB3vECmgR+JnU5g8wx6d7SbtyOXNeI1A9GtOguIqGxrNzvs2tOSa+1Tiq6Thda
3bbZ6BQH9bKzHC00+zRpAd9wabIxKhYCSMdVAnxaRsx5PtFn6KTp5lqNuvIou3JxZZ39o8sKFmTp
yPczJ5TT6P0a7bNe5aR2sAgUPdU3i9lFTHJkqMGoXsIRKCdubTcA0LMi9ErRlxwIrFQ8pGSQoMwN
8SfDdq3+kJ+dj530ASqrEOEDxoKzA6PsRVT5bh4JIYkhOsaibXqXiGZu5bEVAdTY1rJrPdvOVhE9
E/ozSr9OVuQakj3V+3iL9Ss3MN4SFi76M03HOGtZhKl3+r4GOkwfTY5c82pnDuNnibZ78ytdNkw6
a0VaTdnc+S2or+JnEmmsC/Q303t/yseOYAiUhRCssAFFRBgH65/Yu5HODGSBbfniBik67M/UmuTP
mKuKK2kAw2KMHvZqHaShLhdcHp1sOTG8+iwIr/C1wXidXRlNbZnV1YhV5S3XhAxX4x63OOzi3snt
jFON+wlF9g+zy2vfNp3+xdNkdtPfr4/gZCsmyQzu9rT0t8VeW2PVS7y/okImLxH73IKhpKYDq6SB
wS3zok6pqpPxTVMTJ9LoMBJtmnfb9FogPs2x60NhZp1dne0Be/7iuce1gmnA5yOptO+zF6DikDzu
la6n2J8N1Sc9w2x9LVhy5/5Agzw3D9ed9M32v/f7W5T18Xw06A4AnRPyoyrpHZ8g2D/nZ8nD6Jhj
eDRSSe3MZxMlClOwAvhULN78vll4ac8XrrKIDZqL2pREVvIOOD/qPQmdLVNCA9GAlApfGvZL/vuy
pOJamlX33dr1RzYR+bLJMw5AbVlZ/RNqAvUr8YnYINocBIXzIrJa1jaGMgXu565xNBqubJYPY3Aq
uGFA1sBVYy4P6nMb80neRI7QJfcyJMyns1TplBB96lKQigS4zXkX13A1ZhjbogX+1ilvsp7g0xG5
rIdzTH6NgSy8MNPaJLRZFcFZBdQH1y6uG7uz1NKd+aApeEJwCYQc6bIO7uliecJEFCimk8pJAJoP
xXOFlOi7Op26FhV98Rcxi/aRyV8N4UauFAxVWhwhBq5Iay33cxPzb2ovej8FeERRq2VVDBio1lgZ
v9bpK+Q1WvWmttNYLxvo7ljW3p1hgOTNnQ9c1fuUXwcbIRkkPG1WvIyQp5fajO2AEfYgHIF4kIsw
rdbOPreNPEVjVJtmWvsMZXYQfwUtac/eUWc1K+IvnLkGtr+hM51LSHRoGnhqtp7emGMnRZwK3HNC
ARCoVDomptwmIF/TOOvO97nZe01pjgr1aUmD9JD7b+bl/9iQ5pV5mfRFZqsO+JzXPJTiQSP0Ox6x
Em0O0/psJiMkw6IbWdYhqgZmAuVmnMl0QLiLJ42kOFbMj08XYJ26G6uH610cLycMDaJFiohl+Hx0
1ulODnXZU4bC/az/J4PbUF9epk234wj5g6lXhSQUCq67fE58hsqGv46kZi+2MI4WNFge/n91csKI
wCc39cCfvzP2zVaYsPWO9CJ3xiIDiqwPT71Ics8oABOH9aQdlbzH8iaLuN/9NeKWNTR1ZnyMfUWG
xXjQ17LTa6Kx3gUXFEnpGpUHwovsmBlXiK85iRhJYA3iADLjMshC1U/v/Z/qZdfLiCefPZIpwoeg
g9+bT3qtDVIFjHvmcrrLECBVR7S1obf76ww3z4kq4IELoa1Jy3jL6iHrDKoJvwPi9N9COlZri8Wy
p+134fqeMfVlTNSvd42a9AXpg5foFFUTO3GCShcQVPo6TLpNBzbh3hNYu8TgSlGDbgBJIvc7jgy+
0cPoPM+H8LN8h92VTh+CSGGqY6aXirTO7vvzo+jIHJ9p4sTPQQDN5MzZPdEivjBqLpS0Omb9NA5u
qbI/Zl7HuF9MXcx+0mYPqKZklXFcZOuaW7enQVXMzuwIpVwADLTwxoLmMAXMxdBfafPRIShOLAo3
gG9A1Vkw/rOySUs/spbDm3pT0q+IcW9L1bmpGoEOxV0rS0kpvUxO4/4BHlsdkb7bzWB1A/xIb/ZT
Q3N8SZZ3zjzFt64OU8T9WdPm/RGk73kRsn0BINx7tVQYHF9YqUcaShJ6gVIC8bPZMvq5h5vPFVYV
mPqazj1pgnIeDcx4rZKP/C9ik6gjNlFn8MiNdoxx1RXzgW8xy0uNv7SGYJX6mI61c3CEoAA6OHPq
eJJ/93/6FnqGzEnaG0nz8Bcz8HD3ewneyjofxk+4UR7GzO99LJNLb12qr9gsw4dRpIezONXpNAZ9
Uaj0fjDdfNzBAhd3UcO2Adm6Cilw4TEzdJc7Fl+W65TtmCMpBSWcm0ipWrOYnoVCgg60/l78OTDx
5iPvxvJWH/5uljtZ191TODWLbTXJN+xw5CJt4+O2bxGuCwv+eC1DRISqpe5/fZFMQqiVcxOp1Qy8
5RG5ehbpNeOl06cVQ/4jySZuvoCCEu2Y1zB3BNjlwaiO9aZGzveZwaf0lZ/mFTcOpz5RZlqQ2/kV
p0nCIlpglAiUKJXBZxTOSA4Ng/HAJneg8WM1crYFn/2COFD7rqcGSLoBRtJgl/ddI/VUkyyjTxhd
UAxnh3zddDJeL3g8s9KozeEeEsaf4XqrlkHCowfI5VAZpcYWTdoeF2Ry6mvfibWbLNKkOPOKhVVG
jb4jGLDr7maVrwh8J9e9Oz5H8K2xUqcqVu9emjtNTcFrIv1oVzLb8LjEL/2ZRZRsXqTlTKdxdp8i
D9cxbLGVu5GXOqWnGbDW1q/Kghn1imrSqFeiSy4f/skVc5BMSiSngH2vR4s2lAgDsZxjGBUAgKwn
l+HPiP8QC509gHidl1/txDZscsRCD2EynC69qK2OHu9JPuJPt+n12h+qNvNkXhfOTUsYUF9HFnrg
W5qZQEgPIOtexJhH75uaRuXxdwTHYDKUTbscSt3cXMTiTSeJxwVQYvUtN1yJ3vX8ZGFzD4R2i6Sp
JuXSZmEaHUYvDSQfKBIctoDq3U3v1IJ8vELZgdpS/lNUFoNV8Au6svne5vTg7xw7lhdoO71bbKYb
BVo2TjWddR2ctAgczMvNMjfz3dfPFpkXHNddhVqgZtU6vk+ugpS2oeZgEwrxQdYJSaU50uw2Uraw
JA6KKjBpvX6/EBQ+RmBIsjgypy0l5XNOjZ8JsFU+Y7W5zhzLK6Q2qzLluATPEDxW3N2UGfsich7B
Qwy8D8a2LAXEd74mQ7HnFEVqmJ9XwqnOFiCBGbZPzaG9tE1+lxPqj0Mv0Xm5jnBAM/w3YQubPU4h
NZb6iz8joJ4b9iakLSaq6gFN7R+g8ooCcBogaYAyR/uvmIMkj9D2uyl+evF7AIWpFDBoZQJ3WVtt
u7IBawl259JglMX8T9wkUiruv4hIm2gtHQUnot0OqJSG2BtKhb5uLDTMax1Q+glvZDizotVTTGWN
uvaAqGRYBwM9KHP1L8NCUtDyTukssdSayVsDH8VXobGZ/Xpx1lCtXx/PiRAg9W5kcJfbDlaWVSfc
V1/NNe+jyYZUuVGC5fzAVHMmbTb8HcosqS8S9JQfhM3Qx6/XGsrrl1hElLzvdOXPUQREGQHSvQ2j
iJnq3Vru/atJ0N+fIoUmTJI1brg4u+FPDdAi+QSDlqO48aMfBegUH6FhG5SQSey1Kl2pw23SsYjB
biunGhkralmf2HVdaGNDXohQN9pZKbpiBnBWnUq9fMp8F35ZSIrUUdtc9SNGcFYyhxTJdzCt1wGw
r6d+BwpOB4sDeh4kcshIw4eLeQDb0Byhj5HTDCyiON0x7o7DmoRfUF2ctSNVDkXZFYbQf6oFvyIU
iN+6CI/jjQdWzkNVtnQ1IdYgk7+Mo/efUQGRBrNWOT5/mIPB3kKVioKNiVQRUYJo5m7G+W4irNiW
/5UDwShinCTqEMpNaM51CAusgi+yRnEH4yoYSdfiYAjyL0s1YJ9QIuY6r/vgehO8aaKOur7k72ce
hfivsh56XqkCMHiRne3micV+Qol4dAWfH4mPqpFT9TkSe+gr/ujgCKwtcd8Z3TyNsXgBd7w0N94y
QB+1vi4u/rchRQ/RSag9XE4kVqYtPyT465pdde+Mn21LOc4OiLUKngPmlZdjyI9a5zI1UnaYN+xS
3i9WHjBZ3VtCqy896S92UErMhhff4rC+lL5BEmrxNj24W/bgZrMZiuKbQHagnhaAItMzQDKOcUFJ
yl9qGKA4sHSE2aVeXGi/zfM8swC1PMlOd7ddww30mzt+hFOEXcWku1eLqd8VnxrAcN55VtTmVs04
i2f0CocmQRX+abLSirSjQTl4YherkPEQQEbnN9T8slTo1nhRpX5M7HyN7PJw1ztZtcD29VG6QKWV
ulWp5Wr/QVtoe/v5tDm4IiY6qPk/vPOXYiHCvWx10TNCCPEikLDrOqyxibgPHyDQgCO68Vu1AEG0
kycO+tmEL0BqrJJ5PBPJFX0CzIaYA9a7oFwkLahUmeK6dfpkBCuCSwlwJNGXRwkQUlup9EwyLbCc
VfQ4Tl7Z3nBPkEHWfGn3qdnOJEdwvmPTLFGWxe0Om+KBAFpZ+sFIlhPe703U729dDMBB5Fi5yyQI
9O1D3C4o2Aox9cmR9wqpklb7kfkh0kgQLTna9HE+l+r4sEpKx6ea1JKNI1tSpYXcNriQzLRFvktP
H9Wsy6D8V7iOrXSTDuMcSs6nP5dLHYZNavIdKKbl83xNsc41ltSB2HHhYksohbCy5cYDgkSqFWx8
8JQhTMIU4eK8oNLDGkPFrV0K6Atyd/uxZXQ/XI0S2BD2FxJ1dCm5IxFYukPuMSYUR34bbnHt/Fbd
hW8Hf6pn4pa4W0PsOB2j4S78wBGGUC9Ff5Nj0YjflZZjjFT53IR2uHtCrgWXKbjYFwRZfrzTe1xl
wgui30+Dae1E9M2NGUTmzbevfwz5Lw+bO+ualfvFTioPoYBuFr+7cWcLipXsKh52L8swmYsHScvF
7zXtT/Qqec9/CKNSY9cNAfoFXwRUn+uodkFLZYKgu9mfrzKLR1LAEL1VEIaGtYDLrMs/CqpM3QhY
Ipw5mfcKthDg2gAmLHZUL8bV7ddT0yy+178coBezj8p1B6OeMOePdH9IEEZJkiukvhdf3uiYXXaD
3Y637mBElgksBqvzvM4vM3osPEQ7lZCBgdKT9QgNNyhEItReN3rGAoaGFXnEvdMRh4LleGL6CwoA
ghLcOzCEbooKJFG4XDqLWIfoZyqZ/OW1spiIEqyck/bRiSrQIfdZT9T8SFKAd/8f6qxv6GVUSGkH
+IrotOwgkbWDlg2F7gZyqQ5F6u2rA+RkSXQkcCimZLhgITEnCt0Sd5zcr/v1dwVD8CLp+ZJ5CAzY
wV5k+w8Z9uLTr3boi6vrzcp6LuD+wry6v5evZ1a779L6NbQXCrWbYz1Xr4MNztaTpSyp0z/1Ftkg
kEvIp3Oc0cLKVY49/CXq9j+GR26tE84Y7iRCIEhgCw3ff4WHdxwE8HxPGpeKpaTctXYkSi9G8If8
ANjfCACR3vhcSbl68LtemSwmVXmy6l+6SyEsKRl0jdejmD4W7gNLW9q/6lujTWFq2pm6Vdp6FKXU
mkyabMpL7M6BzjexpFHytjxSEl6/hXrW9R+QGeFTHWGz9HL+MnH83iNCnyNBJFAIyvImPCWc74KT
GU7sMetDnkfmKXtAU1a/qnRsgtSRoOvVk4gKGiA/g64YRONl4z5Q+znPJCJ8l4StvtcSxO07D0fV
k20MqsLY7T2IH3w2cm8YHC2F+1nq67g9GDqpjlaGecp5t0UjNVG7tPnOWeSGnUHmITIEwqt30eNE
Q+mL7p951L+suKXC9jtLAD4laCUrGRVE9rWxyF5ScaUsb8w13xzidTc2B3cw/o+1GJN/H3OqU9TP
oPOdHcqW0ApcmxCELt3XZecT7nzO0HTX0p99BR4v2V4h0PRpJGXe2WQPmDo7GH1/grJDsjaTsC14
7wErhJ40P3Peqv2C49sC4YgB8FpCUYrw6is3KLS0904ZOPDRL9KtunEKpBMlcm4PKSKb153dwTnH
wpdT+poRP/EN0U2MXiuvzG4zLtA2rVlyISubJY+a9K9e00Aoy2HH8pkxo/OqzvwLUZJ4eubwsCH4
6uzdxVPbhIfrtCe8nzS8/TIpAOaZVTM8KDuJVNN8VsXzo89oVsOR7dEJ1J7+VH4/RbvIXORfWrdk
Xcay91cklc/9lSmxw15lRWB7Q+k8aAzPeGLBLYU53a03z6fEcQlGVf6AF0hjalKLeR8H8aqu2H2/
2sjCEyqfD2cJvwj8zVoIEyhPJ54cZS8Xfinpvj48ps2cgZDdwzBUhBxnX9RW1TL16Yx0CkwPVtif
RkwUAdhfWWkjNQxsnrdThhg5t+UrLYgEUcGy+yFq5fB6Q3zxpsbZZ/7hxF0Aw9Oy+ZVi5CsJ/ir1
VPXRzHzUpasoi+6JGqsnQaSMsAoGE9sphjGm6xOqvdb8/7TwH89pnwFWZHKi0Ak6Lo7Oboc1qdyY
N8OKy6u9AhqHmQ3EnwgVAA3bCNIB80FlZIgIGAfcsefrL7OR8uvf4vr6wUCQ9Vc0LMvNgIVzlZYe
GXfJV17HovrkAr09hocJ7shwdkn+UComQUO/7B6/Mf8KtXrtcfmZ4UeFLb05+fTBZKwmNO7mbjdK
66Xe2XE56oIcwdUqbu23DLtpyyN1VkLGDtUCLdp68F/X96dwxJXzH9UkmCapV1Qz6t3YopSW5BXM
9S26dbqvJh4VBIYWzdK6l9aX4r8hrLyITSaj+IQB8k0o0tz3muyyK4WIpKAoeUo+54GpD2FdWEyw
fqSL4P6iqDrC6SB7FJR1CJDu2EfCu3ryFNHkGCm73mMA229CX9gqSUEgmaalYlL1H5iKEIvorYQc
x6motwDfdvoAO0S+dOdI9WS34+PjwGkwtZ38fq6yHYwb+Rc+fJQ9IM3YcX18RwPN0ZRbvlIUNMYv
FXsmknIVMSR8HL/ZV5pnrf4YmaB84Gj6TJec5tq9ccCSvWjQzfmfF817ZK+49bGLx1TkB/6jUez5
ATpJGxYNT2HRXvagJTrD2NX7o11Z0FtfWZxqVvuX5FN5+GG5hBJNz+m51QEUo5gaHeowzbT7to60
qZjxC1ym/hczGINi4mVSsqO6SMXH0agJjciiDbunPite0FRql6HjYXKKFXdo6h+hlkqouD7M8DWY
9AqTNOeZgQ2RRc0/a5RxR8Fz2SS8b8if7ps3/u7cCoHYaT2/MsF+ju/bLg/VAPhbUGLmuEZWintN
rF6ZgCfO32gdTMbGNzLpCPMaF1B0y3WkH8oOoDldxnjNiYXxC5wzrtKE7O6g8goWz1tQAUp3Ze99
dXWJ0VheQGBfHxyc5F55Y0PhD286jG5xHyRxm6/pibrRFaGcfP74Fd20OqKorF1wr5qjIErUnB8g
THx/q9dHyeJibtePsAr/oY/JCsqqWezmNdfa3jAiHp1z1eq2FGrErf42e5va6aYDoSzrLHPDcVAL
tWacqmruFHk8DRUG4rBhUb3rLqvwPHm2kYh2O8z6z04n2uLSK/d7o8kYArCUtf1ZmCT0ZbIhPBAV
VNZmRG6XhMg3wmSJ1aHPuHH2j42p1QZHhEib/A5FQF3vmoSTz0gdK+tIjhrK6A3f/fDo3ys/NrmH
Sx/9OogFs5q8C96tckeJ3mQoXMgPFqZFsyc4bunkB+3PX+Ve2VYOPfHsP0YkRfxE2A1r944KBH6z
/GwenJUaLtwCdwSXtLqAV0wZY/BiJ6QCi6h1rtpjoYGm+jsN/0AX+8U98zmQ7COpR6MX27lgPff5
rW7ic0XILfjnf1wUb0tKWtNGdiD155//WXLw76FvY+i7ggd/pFliWHvtT6ll1qQu+08kAkf7plVh
yyO8OXCPkanSsInrBrPwH8gKPVVSpnwCcBud9Sy9U00v4KWuSZykDg0GkiRHYNUBRI0g3czthhcf
Mj7ypn2IXLwEfATvF3tshf7HnbrJ8FNkB7NrY9hTrEUPpQ7La0aW4SBU2MuvlJPOGgdf6FBp3hT9
vunlZoDFFvyj/97pMJzjgedfqzj37CQHoHPgCYzqYommM5H0oteG6jIxnWkHeVQLKNGHz6PC0odX
ywkulQdAkJu6obQ/mFgTQFttU4O8Jk52nlvfw/IqhdPILW05fYA5urhDU5kyBnlfVV9bdnLZHvrR
AdlMZpaCKLM+qidOh/Xg8lalHSIpmIGq0OGVsSSoPZ6R2ipz3H2Slfdy1RmkIGGnfz4FLOOSg9aq
Z+kG8WHhLP6KXJY1QqNcjhJHKCRDTPOB3Oxv1jjDNpZbWgYb+8UPalxSOyLr6wNykLjrrLHVSrNz
+uHSnv5pVdYFT1zllQ02h+CgMsIT7/ocKMsq8FUMqqaaNPCXJl0D1t11u/jkHEw9YrMS3Q65F9zV
g7y/LgMvB1Uh0UVx5dP5BvNWIkpFC//rCSZ35npLSB93jcCJSsTGXiC4nnEaeZpJLLyY4z+JUbB0
HoOv2RNwIwgnmGDUXCcOPlN2Ug2c7fkHfKO3espxEYA8asprcFGFm2F6urHYwGHTdXDzwsEVmzHr
jz7hvpRECnP9g43Oq5LByDZ6NKHuLKIAR8ZzF81kDYYYGlET6Q5Hd/NyDioApsNgomchh0lyj1qQ
K48BOEgfR8nS8kiMYMhI5p59NtSq7nlK57nZlSPraW1bSHyiBZueDNqvxGcfy3cWw/CSA8dmfpvo
8YPVPN+XQItFuYXmga2ZTQ+r7ZoXvdZj34XFXQ6PMDDzeHK0kS+zo3YZ3YFRYvL+RMuUfgwqAmcz
TG97cINOuFvQxIlzAclI34iuDYsQSHM3a7yKgqA5ut1rVABdvo/3CMlLnKz+DjPM03MNkgx9p0VI
x4MO7xqW2GNddKLgIXxkoUZyaGqanPamokdadKgfKwA4zxFMBYyIeuej0kaE2KnQr1bRbARauV9k
YOKzD9ckhKWPsS8e5lvzDFSC7mz31XntFy0k3JHPmNZgwSZRy9cfPgeUwCBHK9d0c8QBp+Rma9kk
8y4paLkWcuj5tPKKgvzi5sISyRrzKJOKyuiFGxEsuufc+rfvN2IhmZrKSsdnv0urhtixsHN3OCl0
fNIc/DSqQzmJ26zpu7cHh9IfFff0ag0ukpXGlDk7opT8M/45iZzShmikK59eJ2rEIdqL+b8x9AZz
Cg4tUPxhlcM2eL8RscZaJMJe6yrD31geCbjal5pABDeX9aRV3/gbA8qTaaYxaIVrSC/Ap2Hluy6c
PYkbC9KB+V+/lEGn6ke8w7zXUJzrmIQdKhFOQdFwC1u+SkXIi0Q7yyCh2Jz2uJP1e/p6RkSvkk/3
6DqjKir/yNKwRUScA5bSOgPSrMWtb88RCc8UNf93s4eMkP6We4xsudKsT3QKVzJ/feu7nkJGLJIG
sKDIHdpg8u+v1SmDPEDascZApkUuVn/5rn6m6Z9fbDfBfOmcrCHSphK5tXyIg3nsT+7ioq9XW88m
q+ixP/sudg+MAD2vCE1tk3R26jP4Lk6FdJq5lephjj9VAVDb61DHcT9wHx3uwPYLXxclAz4NDxqa
G1ZIPPY75DTwvXcVbF1gf0l6tItDg2PN78NXPHzT6GTWs0seiU+F520+EO1c/qNNFWve2qRMRmih
t0iI6UKTP/dXw3Z2xkPnb0p7l2nloA3TpJF4FjCcjYi1yP7AX42fXejlhaqqWOenj+PDYHQzmS8F
NNHTjgswYll5Q7WO4qPUY9AowDVMfousu6Ac+xESGaIT+7OzmR7PaImlWHcBHojQRrsAJwEjdVu2
3Sa3pBiB2Famkjdv5szlfMr8MzzkLXh/0XoCk2B8X5IUmireBwBZGOc0LYf0YykqTjDnjNvVd/Bx
iSXxYExm6VqQoCjXLyb6QPgfAgoHjaX+sal+8tBYClSBgNZ7JH2eEaCiDglHAjRYGchCYtqMqtKZ
0QjkTiVB2VZ5ypKWBrTivnMSTETSYfWj1yww7V7Gj4mnPzyNNH5jdd3vYrGJnJSp552mqtZFesLb
D7zWqMbjQtGEYEE7Vb0GeVC83Ytoxg8bIsycqu/r3naSi6cX2eVSkpSzwf9T/BwIgZVbCOx8KrIS
Dcpf8Ux+DH68mAgbNePsN/smfiDqpRL9cPYR37BPQLcIV6IpA9BukKK282hZLb8QmRHpqky4RTlM
BxXlo3LFIe3K0m3JHqvEPN9axEZTm6un1hjlPOq671vjRDl1tXSG1A9uDWXBi25cnT4CELJAOkyZ
J4WQ3kszylcwqhrqcuNKcpq/P66IDJNWO6imQZ+t8J3tr+7vd2S2sIxp0K1uNkT4AgiDPW+KWE6x
4geomiuGd91uYmcxLtGMe2/TibF5YVfO4Xi7XYdiEI3GlkK0dDNsDJ36yV8BvURH4DBgbm9fGRgG
gwrm2XE+/jKO6f5vMRP6R/9B7Im1xj3q/wfloamcoqnoZnblOCD4iLRgTVHYaNpd3OKt8AaZOd/J
b9AUsZ8IlxDmRLVsO0EFJLohEREO+Z1fUvoKSiZ5weOdPSIT1M0L+VuPvuFk8CfcAJGtoPMtk1DL
d8U+BEj0XEm29QNJN1wogjop2xFM2aNq9vpEZp3AU6S/EFPwKyf4S2i7orIaLglnNGggfzURamrh
tfVnxqPXE4u91Ru9/EekIXfiMqi2A4C+dXDnTEBglNz+A2JHAff51W25OXF3xLgX5dxeKVqzZTCs
UfFcLPYFl2bv664B8/B2QDULI2r5jg8RQE6oG6jjG9iabpEln/m43ct17peudmSl1iawzbTq2hGJ
6vu8VTVFTECTWPsK5qc8s5hbk8Q9GPlV8k+QMO4Hrpq0FwqBYk1NMRnABVOrj6+b3+SQpIg2/VQy
4v3bTdJ7X/mposjJmaCo03GXBsH7V6OYz2VYGrb81sX5uSjJtmTe8mL1xzkM3eWlFRnrI1o2o1vu
MeDQneQKv1K8HbOKZpkUIa6k38MMdl4SDRgQO3YE7oQ1KVCpUD2k18psuiTYy3gFii8LFK6mnitu
2IIICOZnVxUpjubZDYkkljA4TnPmrXZ6SJ4kgAy5J+4WcFrK0hWP0bZOImu/oCu030b56AAvP8vh
mIoFfNv1ZXXNZbU7cmtuf8BA6Am2onOtxFc7JyZbziflR4WJbqkpQqjUHx8piWZOCxdSZXKuqAfi
2/XyFvGhT6Py3rp2GwokGlYr1qmxsC0VlhcNImDKtqMKLqlU0o+gb2g0qCUViLYSRJ1rAS5BwBwJ
R41gYrbn+Hn3p3mojkC6xwImS2aGqhtwh7r4/hI1g/vC8VLib5ZIPEwmMQQkmask6pl5wcUgG4j2
ccpO1mf4nbplX94T8S72WpUVV1rtnaP5Y8shSi3PgO7bs6JXWZUlgLDptOp8J4U3V2LJp2SGPv5B
8PWIMjklI3xhuKZxJikkZmhCC9SsfdtuCMe1Z+qUapqM1IrwIiJGRrSyQg7EZEHaAryrHwljlAhx
3XnTf6CyJXr8ImmWKNRhv2w8z5lwiEN/7xrEPwV0uFS79pRCEJBcPVGYvRIqfVBdrRjV8VCJeQbd
qHMlDg/FdgfJooz5jKHJ9lAxt+GYh/W59UR9BoCtckeGeyyh+uCGn/cXtcvUJ+R+dygMkvv9n3cO
yrP3K5RpEeorFr9ixhYh0uPTaAn3RFZobZ3TyN/o+yeTfI0MJ8e0IbbV0YhLa1rSn3Na1CwYg7LS
tdgxPf/80T7Yk8ba+NrGeDLtZsazNbpYgokT4E3aGHFhzd8gyoMBlFJ/tPpiBtE/d2AO2PY2YzH9
CndLJz7gerUoSoE1JcOWeUvACQZl+qqVBEdZyqPRSdrBEFXZDay7NHsQZFPhygbzLe+cOP23ZNIk
D1GV2cPm9QIpyy+utOeOTq/bkNpgMHm3ix2NakZS0cHg+1xwhq/DZdPlfzXIjUxtrLui9Iz1+YZo
XI9P+EeyEaV4iLxYgxOBW9kFSjnDVZS10yI0lNnWf/8hXukKO32Q3lH7LMzW5J/VJHlRQTDMptr4
DiWxdj0mM+TKdGKekeX/vf/CIIeJg8Do2FR6yXGi8I9rcnXOeZhr2iYwnCLrIa+dQJIjkrtqkC+A
M/Wif46INHCrRh5rI5Z0+MYCT0Rvv9W/ZC681HonE1ZV3sEZr3YLsFnZdarEGJs7Ra+d7mP7LTNj
kgGfK9oAuVgtnNrpc7vdtdQv1MtzUymYYjN2W3QqblGAvAp7/L1m//vNP4JGO4YcuayM6wh2cB3n
+1FEcNEqbAwSbdEhowcU6ZydbC6j6lm6T+/aD0W/FBGwDZiDV1JipIjANI851QW8z7PHQBRRkRos
i08vzIcOxishuZX6pLVOXXepvVPFQOsNOosSLPKMZPRDAty8Mf8Xg3LeLoOSJ7rg5Bsxah6RJPx9
77FT20ZGxX+4uh8+PHRPISul0oHvLWvMXJGy7c4o+VuPAsFYb+XyTQAOEY490wCHdkiZkw41In2F
GT8FI3aygd8au+zC0f+LX2s9Qy6yz5lrClhH1I2x8A6NjgAhOJo0GyumrNzVG6NJWWUD6kT3AqAX
Ab9K4c9XIfAAOK5rLul3xNsi3JLRC1fvnMRFowZGsZChcBkJ+iLHoh7AmjhRlvSIEk5ilrsk1gkX
fyr0pQWhRCV1CbmAufDPq902FBXuDLq8eTknsi/n1T3hze5ZTW/pXRwQmeiEJOp6/YgYsSx719r1
JS1QlIZ2UjJumfeZrsQeGjujcE8/k3YwzCRGXWCd3MD/WTW+vPoQmIPCSuzpigmUrKe6MNx2OXJX
Cwm2A1Egm8jbcglukV2UCXOs4mGhP7KpAWrd4ZORSpekU/lilbBNYrdIi1R/vvSwDOUUWpm2infF
WBZbfGqVQQPWTsaAuf8LE75imL4o7b7XbR+Z8F9tSpzv89D37AhJnDtufQzfpaWyJWLh30f/Sl3f
cMUtJotk+Mcn8+DmW2flKyCs7OyKNMVjgz1iKfeE1jz0W+fpW8+k60ZEJx2hbnwqQpLKFfLXxLtJ
8s3Bwmu4ENycwCvY1j5mtPvYYzvBqo2Ncc0kcb4M8HTwnJKbdi8fQBjtAjfVwSqaY1TGuFu3qWeJ
mfGvDDyW8Ev/NC/F6LqiAvYZl6X3z2iF2EjMpjCyBL9PdvyyIAcAycATadL1XaM2et0nqLcOt5hz
NZ6etwXWem5Un2FwDg3pLMs5C2/vfLYLQM57SOkce/r9N0xJUc7P+AepwMF+Z9p0S9pRNZS1IKz5
0sONx2ere+bjrsYfBM/KqgRFhlKhD/VXoNF69tiRap4j5XmmLhx7ygLSeH0M75Jw5ossRhQ2yyFA
W9dr7JQmfn9dAqDgVBROKgGI4awzmainqDrdECMETJtHjLQ9tDlFlp3fcqz6KGf9V0LUwao/GYce
xkZY6DuJ8LwESYfDHZRYIbOW8nSleX54Md//W9yhYc3N3T2hcvCyrh8ARRKYSehKIjgQkUpKqkVr
WOlaqTIuayt4NoJ/JRkPX5IOE4V5Bb62JBUXTTGf03gg7fn9HkJgVrxn/g4G+2nx5vDQvP3ZE7B8
pPutDtynuSUdUxmtYH0gHNTBPHvabUKbfI1nKMoq9z/fzJcbTdB1QDjBwBEmAB+YXpyCixRJFk37
eero2XvFppsj1mJC59ysl9v96/OT+IljmDsNoppdUQnaJN2BkB0lRyJ7D0IW172jXWvtseZmo+oh
TFdtd3xLfj3aSUIg5QWWYgbpcRznLLgZIGxkP3ND8gkVNfsj1sQXmIUkWxEsmePEkTmq/LzaKA7B
DvU4ICTqRcglgiKtgKhMXMIiANKBq/xTlmB/bCoItEOw/yHtxhT+7nUmi5C6JRSpUCfZY1606ApX
3MYREstx6J9KENo4JXwtZvzsQ+AmRkKkyTrZF4ZtqpSf4jLBwEM/yiv1O3IyR+sRCj94Z8VqiX2a
jgoT+SNIEVCcPL21+hU8fWxw7BY77frsHWWDZjxpn7mgnL/O9fopJWD3DJK2XmUJdZnJB9oFHJZP
y9VYoOwIGJV9uIlQANgAeBVSWIuyXujYyPMK5D4dBDgTxlpRQJQLsevvk7HOwrW+doIpKq8hW572
Z2AJeWrZUh3AVuL3RyR2G9jB5W7l4WBy8p8dc4mqKtuJ5Z3DFsLWQPUGQcjIBYg6IRo307PntKus
Py+fqpHdoPfn3aAhko0kOid+mTOMG8xZu0ZipHDxA/Bi7KxOzAjfMTeYRd6wdwuCO1qUvLaWfIZi
VDPkFkYt+skuIms10sr+G+raJMCvLunSQ0C70iUHmQKTPHmOr1lzLfdk3yp+lIvEGTLOR2ELULnH
wCEvEwmgeUUTo+2+NuvrtrZotP98ek92C30/bNDVhu54mA+67EjFF7MjcHDLnkGP3V+Iu2ZfKz1K
dsA7DCpI266bjzjhCJTo93TY3HqmDVdgqlSW5ewhGcWJoOKbpN7N9HuSUG3Lt6t1lNJeRE9mMOUp
V7nKP+p/vKDwGIn5/cbVwkQE9aVUvYrIDo7RLLjjM1618B5c/qhjUldx79rIjCDfU9n2tMfgSKGi
04zX2H1gVLEBwN8HBlyKH3OeSDQEGy0fWT63mMvHoqKqThoVgTMUbCOgIVHvAAnh7pYM+0FdXdFd
wWlxHVuDGBI0012WmOoRakn9lJKii0c+Z3CRpJ9MI8a1Erg1Fmg6zGr4bldP41lCJ+F5BZWkr65k
LPpczvWk0aZ7AcejGHpmXQfPz7Ic9vOYaovsyhubjaiXsl4e2Vvkxt9bHvPR2+lanyD7Bkc8kYZQ
l5TW+7TgiubxRR0vHItO8RgoiUdHoKlHNG0HQCCjiQkvnM0v9y6o1xyb3QzgrITNKV0RYx+GgWOV
KObFBLLb5O9RTzAg5dt/FNW2mkFaGTEkgnOrej1Nce89e6HJGF2sLV2Tqku6vAolFr5yvFlVOmGB
xBSJzNrWuq8NB+Ja2xRDmuiOmawjHuezD9H9kfCgHRTZUj4THAVsVE1a8+95orJO5qdmnSO8MJgP
NyG4SNCcsL9KHXZD/zAZ+JqkiFYlIBqXVqba/6k+1eTcmbn6qJFRtwXY//+/ZTMtQDuJWNFYeyBJ
lC48v29K2lrYUxvZMxxT8drpg/p41Sf20KnzTOQSRz91s0qDZpdAYUukJPOkelV8hdXOjLbdcjaY
RAykA7TRrpi0Ubl3DWHxjoK/3/UsxsYV1qxfQJdflvNNn/zKfeIWIueW0TuF4cbov2Mwqb2rMr8L
fJtnhPyq7g7zn/SvApp7gHwaCfqeC1eGn5B/EVDfZZpRP4YJKpl8wmn/hxzEY900oDsOHZOlhh2j
FSM4sJlKzyAMnoW3+iAK4L3rZYkcvrT17fl+AA7t2V2RzOXHZToC3KxEa/xpnbCTgWdAdCHCaomm
NOpL9xQAF/P9ZLGjpUTkZ0WWGzlynY1tvetU8XYW8oQApIdfDtqjKBNp5fm42GCYrtd/r6ZokRxB
Xovs6Vj1CdbepmJuZNe6fe6ZrVevxuoDeNlHEurKs0sXpfef1SJKWoNzemIugWOT4IRkQpu0s+ic
vK0b9OhRaLbSYojz+VH8Tv2RKzbBMQqHSMfiSxTi85TtUPHgKw6N869lz/OSZ2AiVRswY+BS65Bl
cPAmj49dWDgmRil5A3byxCeX6XgETD+35as/zGzEGTVbDqB+vq7x9nJLmHvEiWzcSpD8S0ceArDH
02YiUxekM19+DJTxZwcVCR69tz5Hl5xt0oONZudg0puME3ElY7JNVCinjFOxdyXXmAzRki4TpVW3
2nHoRX+AisMB0dB2uV2e6wVpjgkVmCQpExpVpD4Zwpckqs+Fv/7fiyjFeVjcy6fspHLWLIitKQow
cvb30ZAsllT3hssrweu57VqTBs7wd3jQ0wjJmHTpMq+5zImfRl022ovvU5UNh8qYW3B52zDGy9fA
9tWWtHrp2qMju8WiddVGL6SW9EkzM3iIbw+IEhC1Qio9w70sYVLaDG4Z1xMUTUQrPIQ3/x1rkQyD
KknH0eeTlUQ+hQw9FGJjGYwzTS90fN/kJw9/Rpr+UdXrCA7V58h69BLrIRw6TVSmIzspBRaX6m32
kI4zsmSqsUCzFky3Q968ySQOf1L00hVRQgeg4TdHmDXCbs8tyltHARmkcPivg3wVTpmmic9gNdys
s88g+QFJVQj1fNhlQcxLmFIlcUUikbiq/Z/uMTuuPgXWuei6I6BhV11/uY+N0I3BjTk23nPKvn9B
pqh4Z4thP0YVhhOV8hC3noX8tSbjZ98b/WJQb4n2E91rBkPUcPkGCKrsLXosGzTudApTqB0zmPGC
QXqPYfvR9ZYKYDy3kGhnmALmhpLUQI/3uXdgAGqyIMT2YIOEWLF06ChqkJcRd3Ch41cHHbjWjIBJ
LUwoDifXN71I2BwSVlhiUtFqGCM2E+1dvbs32KyNGM/UNOMfRB7h5sGsaLpoOigk2ypxCqe/Kbvi
ThDEdqEzIH+8j5a0KdQZNq/0vyON8XvMwP9GWQlV88Uu5wj3LruAwDiYS0l5Am5/zhsCkwPFqVfv
Ljq+keMAM3BydvaI6fd+0HGin78jpJcBh+Tu8NU1Z3ig6kj53rS5XGgQRg6DTl93hI/UI+ODAlYZ
CusOyJG5FZ6tT05OBDwlOR9Nkx1AjnG/G6B/H2Eoj+u4zeFoEEIPRxwkRaEwOmDHJiRnU9FUB4GW
gJKhyLluZhkhoKj8VT18wTcNYXPt2pe9JxWRXvzCQvLx8QtMT689ZIY+LkKmuWFF/4O6gOhfhVMh
/hpU6DsZM5HRoHtjP53kHbp5hKJkZo1j4RsAUhzs/DgfzFs/Ram29ytj190g8iP422x4t11IZUAF
yLr0oob8uPOOZGXFOEg4Hlg4XQL6sQmYjRaw+yij5NCTMzYV3DyOZ+S1ZaZItuPMfT17bSUtwnsR
5PX6jSNRSq2FKj8OjkorODjHm/GF2VZvHgLuNiq2q53VLG0t6JtbFsUauqWtjiA+GP6YAKe9KHKL
bBowGwQt1Z9uP/URQRryyH6GVUuKqUg2/8/bghscLQPE0GnDg+4QoJNHEqqrxOQYFEWb2Es1o3aa
yCzCDNQJYeW07Bz+KkdSFo2ZkAojPfoFKT0xgX1T7OCxtIYyRzOq97hOiUGDDePVioo7kL0JHye1
qihhMl6lgUeA3eB3rlN2gq5hiJq9OFy8PNdCtMvo4wiAM9mGWPi/prv+9ISpAMFsxr+QFACBed8n
+s+5tUGnhl5kWH942g9UV5kNHP0oWOXh3y6ILfsavn8SUQzSHB+8gbT2/wu6aSOycRJsl/xEJsFf
yNXPXajP7zxiZJfUdc9RS28TIeHR1zS2UCkiFA5WEu/4TrTJO9gBKpo0vS6fOI1JNaqrWxiYzpaW
fBMb7jkY6YaPHWg7hyOnNqc+/gXwOf67RjkS2PbK30b6B2kmfXhHlrNRH8rN97n3s3ERExgk4zC7
Ul+2byHxwXS8JMXhSFPlBDNgz6p9rhLqkpHkd/rviLFpR6HcGCp29h5iPpL+nqDn+x5nCDsCtLTY
MAnG3sJGX0TgvmwnNdawO0oavUqz7Eh3wHfsoqng0uWK5kj4Rx6UVimeyNNjYdaA8qxQ4j29E9t5
Ms8mfS3H3PMKp6Fj/b/Zc/Wq9TY1mbq3yygRT3Yu+VwppJ/XXBtKdabL70XGWEuQYoB5c9mFEMHg
RAayu28VsDoKEjQ/LUbHkyhM+mE8kO0NAhV3Sza5M4vQWC2NuGdOf966ztbL14iIscgA5tQzJbgQ
WGYCrP2InEGwzZTPCA3SiSVXX/uWuNX9gR1b4yif4yfsvMUqouUA9ZZ2shiTosD/2vSu+oDLtqCg
6YSdIZhtjSOo+ztpMFU9S/Z/7QdwbTCHjJ+x9AC9VN3N2ID3J1vWvo6o7LLWkQf9WX2YJJ1eTZw6
j4gHYabYH+dluatKibqoKrKIklh4i8Jr5f2Nfr4h2nGqGIVnWqUD76qBrpmiG1fH7c/3alp4fVMA
Ny77kXHnbIpdSB0Lz8/v09qPyhK9TKUOTAXdFpPzHj1cCH2oXksigktNgJFIftWv083CpbPb9kwp
xhGYVsamzILvito0kjDc5T9krXJRzGjydb5PWnG1sC/6l/KMSUYhYj2phy3OqajqQaI77l002tFJ
GD/ZkXZVOQNuHFXRxr5rzJbHMEM37jKG8DAIyWQjywyItKwINgvBBQdWd3wsjiN1K/FCZ7UFVgDX
TkVamaD4wcjJ6GdbzTUX28cnSfAGgfk/7Hwj6jSK+oxexEbL/u2XDXfeITng1c4Kb7LWXhNGUwqr
qkxOK+xjD3nfjEVe6HaIiYAtXuMnCOaQxlnxZzH5J97t3Kz8Umaig5YmXLiGIsoEuxm8fX+geHHK
sOp5JCreP2esj65jc953v3dTJwId5eNs5F2Bdb7ngxDGQagYizECJt+viKc+d+zsDYngn/kL1EcL
quFTpKk9O4zD3pGnuBkVvIyj9XBFjke7rPR6hyKvnjXbg7y0Jp2DlrKeFrAo0SRJrpl0hAwlfgMw
T1amciDWwe8kK35F5yLLjaZnJIDxXCMIFtPzYVnQ/y2Y90kwTsYRs3kTzOVMJy23OoUwoRvZ5/I4
854INSmunSLVizOJfDQ/5YsioUH69l3e38C1kz1y9zOnFxXxPEkVRDTof3mV96DzuBJGgwys6v/S
ZAsG/fgx7bbCNpMo6gSr/DEGLcum3l6KQJ24dwXRFinyFdRkLIPyXfpUoh9mTXqwESkqu1PkG9z3
fGe1fACphfEX1OH+Fj7SPIPTiYs8Fv7CGwfe2IPB8Jht0gp7j0hHkF70U+WHwPrO7+c4F6a0JyVu
dTAUjVdfO/cdcJ+xHzd3KrRXFu9z9VqqRfPVcZ2xGL0VigU8bXXB2JuPM2Klc4O4tC800UfSLS1Z
504HcQ7m7zVdnpKLyAdmVyySMRbFupBZGry7V+100in3YjTn5zDhLe0PJ1mC/NPDZKu2aHqm+3cy
quaw/cv94zt0QhtKBF2PsbX+yemq46If8iEo5Wn+6o13nyuaJhRAmaYAFI5LdMaMdbBVb1kg8umb
Jpd1OoDMnGKA+FqhiXtdnWQbVp48LuTuTDeFgNVR2pxSsVW265oKv3MUKgqAekktZlKTSm37H+7i
s+0PoU8yyGsx4dWc+PZ/AfcLiMKpO/vynGeumDZLwGsY5fFeBpuiffVYGCaYc1wV1MbNpv11arkD
AJLfUgX9R/JdEVfB0+PzNl0Ge22//1KBDRDwwhUvFTJWAcwhOWVtymHTEECEjiZ4rEnPEwP7W7RM
/pl8OaiWUAJhMewK0/ptEj9zCcWT0nNmdONDY7umVGSYZpeknFQ0mP8n3iHo29rHvbnlm469nrLx
kfBCJS8ydj3iRRhKKfZRbmFC+FgaQU+xeIDKWWig5pDWYmvUMtx6Ml25zrCFeVxVdsv3HlucQtfS
35fuYWYdld6GI1E2nNy82oaNnkrWNRnlODo69lEBTuzEIM0oojmTllUgIoE74uH61aJ4TQfgqVAr
GvMCmRjuQdhfgb6hIRnkgwEjIXOkoRnOE2Tqh8Z9Jbe+iiBiBnVeD/RtyRZ5NAfGRWGT9RME56uq
zE//nz1+I6JtjGwqWAesh7vgRU4Fd8462KL6p36gHspMk202FlyFn0/QAJuuEPwEt+llTM9sgKh0
ey3XMNPKXRWRvJMIeC8NsRFrwYtRFXEp5xFs2yN6PsjwDum/dUmeERMKx3YuJQYgVxPJIjQB6a1k
OKHVVsfDButrEWN+zhW1JvLWNNoq9kKge3/IrDI01/uFmU1I8DT490oJLRINR6q1N+BvO2gXsuAy
Ajxaz8doO4Ls19JR8qnOB/oJCDbR2O8KJVyXMRbvxGBywVVyWpNV3pV0J9otEl/1e1X8+U8WJS7x
YZE3D2ZOdGQraZY7eqJHXOQwYLhoPsYVc98WBSKd3/EimVJdhZsAkHrGpx4aY+K/tYoDeIbp2kZF
m2BYgzQ0pNi67INlKDzMs9zTiRmQEPLnppmU5h2tyCtGx/ffLqHfTTYAMd9kT52lv/nB8gnmFL9P
+nQ60Kx8zH70p3ud6uemapd6bYF+18aacVTiPejqPg9S0Mdn4Yxg+JVQ5hXuGf3UeK8Z98WeVda9
J1zPJ9Z07y2WFsZ2zuC7XB37Tmy5vnuRSvO2MiJQPh8Rw+hhm2DO1e5dLJoTZGl+2DQ/v7RBGuS1
ajPA+n9K+DiDz4a0V1aX66JXGLQtsG2xwta/zNk7snW6sp9M1yRC2CKXvPrCbkRDLOC/MgZ65/hp
mdJb6ndNpUl6orBrckuSGVvwiMsXxlWpARWVoJu6MgjuqHeGB9Qo/j1rBRSx1YR1Cwhs9uXPVqmq
+uCW/qyEU0c4P/pIF+NaBIFdstTQyBn2EPC2auH/9NqCsojBdkyl1+bQxqjMzvTWXXW5bmLlCB/p
QpmRDvT1u09YjkV653eFCrbhwjkXFGMBidviDg2jr9vgas65gln88eou7wxTp/fksJD2N7AbO7lU
Mxiq10xCeVez80v/4QyODdomjoG+E3Or4Ipsz971v7bwtT/zPhuc0P6WC7DeuGRSLfvuAQOA5an9
H1HkpmTibBTZArDZAsQ1QnjXyGorUnwTmgiSCRamD/IGV5Yq3i7KtIpKw9OARHQdysQP4QJQv/qV
9PoliBQN1S8tOZV/ydCFk9VVQwzXQmDJVN5Z+HgnNmJnGaYg4RdVJthf1BEOLvHj3LA0gVkxIQXh
sKOWReLvojRt8WiGePVmohwwZqBU+8AboFx0mDQnTSLWhaVArTdsB+fWXxYkfOzzQanc0xwofFKr
rkC1MSHGzUe061dtKeNNvspmziCcusSsuv3TTuJcvnV9GBjB69nqJbxygVlBUo4syjkOdykn+x0Z
Ckf86WhuJcYefEdW6sqVHKjvSVU3D8oSNxlvEotB918qjIuVA0pIq4EgAQnAdtZK+i136TYnnS7z
GF+Z8ceuiwjSQa0V6yfCjlAZd7/Z+qESOOwmMSXz5se+8QsdAdLweMbreP9JylfmC2eKrYPcYOvI
I5K6RZ9SFbBgIDFN1Lr7Ot40tWenZffp+j/GVbdf1UXSGUDh/P/3RbLtNhI0EfaNdvMdFpc4LEmE
Ay+xbxUIVgEg3G8+R9nYUW68TlO9iO7WW+58aZXDeAIN9S05sjeuwxS5wBkj/KT6fVKLoFmY72X5
lmunKsW1MRmRPuTJkh09L6Nb9ZdQ/+NNEt9dYzhp2VvtkoMi8UyE4Clc48HwO9nbNtSSFNGyXsm1
v/gH2Y//QlqHZTASa4MH9Xo8cNjis/fS375HivFIPN3g7UjYR+F2s29rOctrv04UotC7nYEjkD+w
6f+bOPsbKmN9aGFGqua2x6rwzidS9BjRtIim9AgMHKfvCCretvAcnTxsOMFukuTIkol2Fzs69fEO
17BY5+JPLSp9BX+edizRLIB5jok+L+czm0r/iR2hJEtJt+gMli2E6xSTn+ohybuMFoLoXKyQIMXI
Wq8N3tSrIi9LX8QH5XCjoppd9I/L0Hzr0ay6XuuJ8P5BpeAlyn7ZMkEOE7NZR7OFjwJV55rCsa8B
w6M98+PXoXd+h5RKjGn81WcNfNlyYjGssn6qMpHcRqFNi27yTIHdAbD3UXRUMaAI3cf2oThzrIXq
1VP1TDJ6p9cvTheKFYLoHdy2jcSiQUoGpzWpOR+ooWeC6mG47OtROvTPzhJWj+HrG+uzLDaRhBbD
MvUixbOtRJYMdYD2cEyOuW1+VmAMFzdEKbIndzWnzoRwglXX0vj9UX+GWuS/AgiKCHV72QRcCaNk
BrzpuPAJceQvbsGnPvgrp1QwIxbw/tiQ5Vf+NdpPDGG1bXvb9GJhSZRfjIfTFnKeDXQZrTsZgtcl
+TvVgJLtGdM9rJyNHseHCGtptg4W7eKsF218eQRPY1/JudHwvUp38SyvmfhG6swHdHw48lweQ/2h
YEEPWsOixxsbpHjFjgXPCGO/kqDqsWZHd6SGOknlwnAvto9odOEpXGHvmEgKFHwijaKDRHMkilLG
fcsNV9JdMeQT6C7ZH6GtGNqdZG/cpp0RFJCWJReUU/cHKFQ30iUH4aUQJYMdi5LNyAj94riyjbbo
WT6QfQtJwMNsrja6eb2SAwngpPllTAROtHDeFhcI2gPWUw3fMdEdpea8hQdrZh3CUtX5pFvIXpcY
eMvnnqB5np0dy0loLrOd/X6X5nl8NitWAtjG3TJMQ4c3ustm1FCBMNYcnCBVuS+gLUvHlbsCATrh
+Rq6q0Q3xr02Jj73BoVLnHqy2qRmBDzmJr8HEDVc98E0kvtV7nLAVJ19RqRuDxJQXbEPRi/aGqzb
04qoMyw3O98xqdKJ3HkzNPu1+fdwWrdM3jBgFaSUopcQXcb/6xvnGYIpX57qqRrIBmCKK5FusqYS
IBn27B6zpSxwt1LSSuaBorOio6Fl5rjDFJqNIzdrJ1GOfJdGyacTYQiOoY7NvGmdRoJLO1EGIM9v
wr0ZRKjlBO3x1D7w+MH/mZbomYrioX25CR3m31+3sRcVW6yA95PFrOvvB4ANSp3BtzOardxenNal
2ODjwd3nJ8qA8AlvvE/r7kbg8zB2N/znSvCLb6CwVCYasD+qxoG7l8Qj6R8+P06OTBd8ZFELsDBt
P6YQaI4J91N4t9KBy4LVFFe4YpJvCuAYtGZnZ3DDa3daBGicv2IubcwY4N6VdYEhKyKxV95yUr5f
8a2Bpu6WmZmgr3Gz4OdgP0TtyqACYasY8z/0QWlWDg4ejVwAxZgZnwhF42ase7jPaUZ4Vk8HDMtI
5s2novbd+0zwK4xbGV+tvRhmpS8o2hiVw/bjo77a718qWNebes1ng5hYHm/MWioKT+psvHxvhCct
Dmfh693Ct2sdUxGx6nHk7c8n3EFV28KDW8V8boVF5zotjQBQb+BXI+zU4208eVMi6eHY6/l16tBW
2RSJMKSg9j0JMzqtg7Rd04HniAE+4G2/OAPEx1Udf4ZFM2pA1MxoI5ky98ONJ0KVjkaesjL+zMZo
xcut5PVn0a//wJNEaWHIcF0Q3Bh1lG0aPavTyd7aA3dcuoUnxsfeC3QogKI64ruUOAi/cnr8gUWX
/IWcF+chUgRIV23XZCaSg3XlCk1l+o3XUv6x3XKreMNbiHJ0ik2is4WZsYY9ymoXBMsCxEHQWAQ+
iOyxWosU8wKaB36GX+hWrmuuJ0xptJ8IWxuhxp5SJoxwQzCodDk6Zs6r4lZjoH3ArxYSZ0vgMiJU
ASJgGNikY6zxRdWDwYleUcvUZ73I/+TM4WKfDMo8Jw64fy6oLFsC2NegZeG4KV9Q/BbEPNGs40/H
40zuoHQLzXTU8fdd5zhN8SGksDmmM3hKBQwEBYvYfOnqTSKdz8VrcxX8RW//vRnLHV1hbLXXuuBk
PacbW935mAs6FJ+/EI/4rohY5nfXTjC9BBU2A3gr0TK1W3HwkWBswXCdB39llrBKLQnOuHaA2Fqt
OQqid1ZOtbOeulpb2UjkH99fV+M71U1UqTBd/lb04UdB77yaq0acrqAyOs86yElsOS8rzdd/kTrr
gW7EglZQA5aKj88jyAwEJ0HW8GeF677o533AGHV4hIXxqJnpK8CbqabvMspS1aABdZYKDXwXcL4J
YW/dUJ63lskLRczYWj/D03eNPJ3az0V9giiqt9F9MFkHuHzbGfihhi+6SdRO5fmbPFydrh80IeGD
mUChDC+TWGRw0jWqtBthog3JCOTeKf8Hytg6AcWRrFer75y7w//sZQe9m/uU3jNcDQe+BkmR+n5Q
eJBNVWcZ3mukLxUgd1UI6ZiSYeQ3fjBH7Xdl+NX/OH9dMgo22l1blnUt7bkkYCQ1X8M/in6UxGlf
1J43/Wq2QO+0bper8r1QancWEi3mQEnvXXE0EEDpQIzJISesyXNYVt8bGRBdDlvl+tFbTPqr+dWp
1hrbS1MINyfEE4uEwz2CIEg6Pag8b23nztfPov8CkTLNOgHlJVESWZfS7Io0H7NsLwmTLK+45PTp
Xr5Cbr4U0BBm6hxy4EoxneUngfQaaP4LZPr1t4CtVAq9wxToZ0w/x7NVLUscuMUjZoYiPxKH5D1E
7F1DEGgCizuKCt0jINrvZORJmR050htE+UnhFAiyAJWrdNpGQ1KYqkIHO3Pv/IovIlilLv0fsQR+
bcJZ5OxhVrbjqYHEbr2Kt/V65LV0YeKCI1+1oEdY3Dh63bWPzeqbjYg5aDtUxFLPVbeAjs1eMDR1
yhBKTSy1K2OQiSF0MjPW4nGp0te4R+FHHwgMO0RIxRbMQuweOLBCNGhtjA09TvvR7dH9xDglTLo/
O4CX4a7zBKUl5FDgz2ZfS/iUYx9RSV23ZaHm9ZMPbOqMMzWg1wmKEmOvoSo8OZUchSLJi2qXLf2K
on06ewW6c7zBkvgKKGmDR0clhZke4P0KEtTew8UakxMpw364oCICXER5tOt2NPlQ/LAPWjC22Rxc
tp0kaNfEwqnCxspYykQzRKxVPW6UqwaR+guLWKxkcFI0eyJlJgIeCa9LX53pmX0wBoANPEW/B7J0
qooVw1RSWM4z22ho77mXOWZsK57VLLEud6VpOWL35ol5Ky3GPA/7/tI0mi9QgRSscPerSRBTQWnk
AYudj+SZdzRcSqyFOT26D8iXt0s7sBw99yTZiomYuJ6zRGx4R5Rqw5vBPGiskS3doeRujAAoBtu8
GH3JTn5ySWNO0arxhP04FBwcgaEwCEfz8yKwmK5HMG2qGfSUC9cHZcXymSWxpMmj2DAX8KKJ0Tjz
yDXuXBWRG+6TU+v1cQ76+TwN8hFgyJH1WgXNcGiKUw05RPBhEif4+Z4xFNX1C5i0XQUTVkHILOKU
Y53jmM1NESnYl34PiB9Kcr/RSxXqgomH0frh3ybkWkyYjZkOZUKDWe6dS7BJgQdwTQCo5e8Dvkhr
UhSjgJl62p4hUgdwVgvT0tkOtowgvtzPFfiYvnHPuFHIFG6NnQRRGPao1vVOBGbBUpOd+0slo8FS
2afhbdLplnjfbsAtizG4z2k52jxVoiCWb8T5BEVn8tcL8KgOTD2LZy+zEGP+feZt09gIVDZgUvT5
biw/gaJErVpvwp4f9s8d5DYVkCfsxd0vz5Z2Xy8wraV5ziw0oWHNW0587bmxRkSiySu/RUs1+0nh
WtDWtFZsXfGcYioa+xaCkwYG5LgvU70WCJN6+HnQWR2SNEtyDN5EWphGk0Gzzpyru9zlgQ1ir5DY
csDuO7hmT3fUM9Eb1lBK7XrjhXKePc2TVI6DdNQ6GQXe6evj+qyv8IGyrp6B2fj4q46Gle0+WFVk
xVZdledJfF1LG75BqH6Lz3ReHj4sz9yCe0ECw5guXDs8byfUDe4hyQ2EfD7BZQe8pcfTzJl3O9o2
gY40UvYeMRWofV8sTmlR/QmB/VCAtrGRvpno8VMnHWsAu3daeqFajQ4LpimVaCfOr9RMRQchImAU
u3VidegPE97aeYGgLs9rQR7GijijoOp27jTEswH5fVmVjMwVvw6Sfp/vIeYbWyUZLQZNdBTieoeS
yqC+o2V5B3mKUv/ivmWErqpkk4VKoVbtFi+ZOjSSyS72thbl96HO0l1uLUe1YCurI8qh+mqdF5g6
DLJMsDn3QcvCK0dJuPYew+sIPcydH48C2YM6Vf6MA30yOkxrRXL/JDRLGZj2wo98wjHtunntRoOf
HFQtophW1u5AmxScM4Zpgt8m7x4e+UzlB09Vy1yDPgcC6y6GvPyHTq1kc8YR3s19uIOFs6LRafve
SMAviSeDlypM+y40mlKPbRS3wF/LtgXzNtBhhUE6OZpb8dl2j/+xnVDTrz9DfvcsDZiQF9wJCwtk
jkMRNQGXXVTHNk5HcxdB+Nkom94B6R3hm/S2xO48W0X5rTYLwGvXklpSq3GeUaQY3u6rVm28Qe/L
gjVA3LP5qYmH1p6S5mzZqDWiBOwTfME+PCp9qdyC2t4uDldI0xx4FBpiUbI/VqUkP5G8iNepvurw
P+bm41FgivZznzgGZSQ+bX8a0Vr99ZO7Z9pCGV08s8aUkimW+TmxxAirhyRIZ5Lb6SF7re6vw/Pl
z9GLjrHe4ups8tY9qZo49la0BODdOeL1fuUbkECQ/Nd+5gbdBIvBKC8w7ioS/NYqsjmHpDiwS8qC
CMKDoD1YyLR63Wu9CBTWIQiIy1KrBS0ytYrWuyEN8zIBVenEew34UsljBvFre5ovTph+1+f99937
zOQFnlx8X7RDagzxAQibm+LSFcIh/qqtnRfDAJbY7fwQYKK+AusAeiQppc6Wa7WSoND2uFcFbR6G
Ik+zPavKFD++cM2+qt6iN+ZzqfXlZ/sYwIWnY/QNgTQVA8DUzv93/ugIImifKyy92ssvI8+3Uof+
qYpj11eGube2pxKJ4buOGstFQTPJDF4f2sr6eT6egd+8AIQ67/dwmsFkVq/LQW5QGJTI2E6WWfNm
mfRICq1zgseoToKltxisWHwP0x7JFYjPmcPgGwAYSTP8zM1mVMBncB/3jQhyULd0ezr5YMTWGImj
ZkYXWqbommh5jF7Se6mGSxaJVNaWWJ+bDYzsjBe/1r5PEcUMRax+6tlxYDcwsYShLpzS5AKFzUhP
KtBub+hQ14sEt4v9Jom0slMQgkfQlO6NVbAden33lP5hoGoWbysIhk3Ek1uYPM2Z5dTLlI0erBl1
D+JCXhFbg6ZH2EEkPuPQcxC7TdsBLHKCcgfFbx0LpIH3N8GJxOwkBHNDn3/Nya2ahImU5khdAoxc
HXeTAce9WDOML55ntJS1SjFITUHdhuXJlM7PURW08ToM0eXwoIkkTa45A6FjPPVJXQYgKG1dNQ78
arfz1Ox1kOX7UlrgaWeNZXtFxpJHktOpikrEwFifUk3/HixoikSDJ96vqCL2mm3EhnbOpogncH0/
R6TGBzd66CCXk9LR4siu7zFWU+wbezBwLM4XNR3I1zjLlNkHWlJllihNLe9IUUG8G5xG5ww9W1nD
gMqs6Y1TmAQ81TvnhUybp8I8BQghFS8GgqKSeWO9R5LGDOInNije5U9zIAtpvS7Lnz/5T+Vl2N8J
6W9nj3iWsuCHc0jO4PDVYqMQOiFqYY9kP5lo2RmmK+KLxQW2rFiDgY0p6rnxoTnIHAKD02Smaqal
txWVejKKLMJCwPuas88b/+11q9mRghkZLo+PP27qLoaTWi9mNDENyxTw3orP4AF+nwrmMWb2rNEQ
3yz9g+DiGgE4MH3OpnwLZZdfdL4r0tl6gz4/WygayuJ6Zp1xHHTgCmspcqa6R7pCGXjEvDbXpcrP
FBs7acW9gi8x0rTfAEqSehh0ntaW+hN1lPLtoCA8WppoFKg6OxpGB0+5Tvv9rAK1FUtaBHBTGVSM
1aNWEd62EE0Q9ZoOqHQnZ2E8IMAjMwdvwHjg8ymoFxIZugXXUJK3Gs29/I4S1yiStFG45fLmmqbP
cj1gwrDQBnpu8IUro7krvXAlwIqYBAlfqYpipwLhrhqaoO8PTPGVjEFXgAhiwHajDSpO28LghlGt
M4QNPZwf622KlpP3gg16bFw1wNMJ5hqRZh/+LH07En4jrcOcp/1HVuSuuEboEOQESn2IT/gtQnK/
xpFCvAKNs2OMuaN5p4kWhgNj12E3EaOGLuyYqQpfhgQC/H+66Q2QEfsKDvR7PPl89RjnX2Hlh6Lb
VEQDPvxXnAkioPPqTUqFUL3KVBx+Qu9vGjNB7M6UCDq1unZHxJ3vL6k4p42U1NnU9KwLW3d6+tij
bTpbQQpe4tjoRCs4rLQnkqsE09nwX7m296jGBJEiiPvcCgxH99xh7WSohs6rm5Bb58b7wp1iip+3
byPxrafp+Sr4no4J5QLAbghxn5rJeSTDKxZoX35OkMNON64u11e4bKTbUsZ40xSkVUrw63GPJkZ1
BOr2vgybJ4UhSw1E3ec+tqtKtmsOFyq+AzFJ9Nfnm0NjvY+9XqVA0jWIh5ewHcFcRVmdFIejv4O1
iiTTgH4D4uSKVP2fQJwIV3UWMnobM8A2m/c865mHhOeidM/MtE49NlzgXnt/csr6i8UwzFvI/5T2
bhOgK//yxHuxuvR59dWNdNzjcjxcmiDjIc3l0Ubj331/NBMj7455TNQjMDrLmbdwlB82Uhlk32E7
cSDS33usV8lg2vmWYT48vRNGZYqs4ZDZxzeJhLbzErU16M5NVWnymiPda6mPACMDlPo4s/Z+Bqgl
+DNViaiPGA6XLV9oZejobdJikupzw8Mteocjo7LHxUSm3fgHYy9MYsUqVQ+oJQgyNjLX/zvr/0J7
LrijAdGGasYK+0lAbFmBq0TN73qdsL2WR3SaVxuMHT6wCLvWTsggt2eLQ7jqBHTw8vnMWUsm1ISJ
8ths6kbiMJw9kWeklkKYu5pDjmV/rKr6TajIxl57LU2s/olbnpLDhUbbyFEamQAQOSNd0QtK8eWP
F/Pa52/kykCgCQ3vFwQYCGlQ7usoHdATywy76OgE/Eqn+fIu6wUF2gFvyXGV5U8xn53PB51/C/eM
1zv7CTEQ9VqLqjgyxScrHaioYultBJvoZ5/smK2Yk5vCdpKxxFXAnvObziVlwcr52LA3F3jhnf9x
HrE9FO58sYd4c+bMVyyfEtEOtdyCR72tLmksL7BL/YLaJDUFnmZv4JD2Y2N9aXfNI8JNt2zWNUwv
PWl7eiKBsjdgPC6Gw2tS4OLfH6OeEwXpKLpontGKfVVRp1wBrLPsye5+AxZENWi2n9ZyR0QWyZQ+
bpuzenBy7DqV4BomusOQDKU5kvRzoiIg9lKNwtWFUTapcCPXHxbCyNX8mbIa3XRNA3A4t1FPH4vm
fm/LyhOnSxz+n235oXcX0kQuYPCASarMBYhvSs4EjnHmoeXaIuCBstc09vQ+DICXXB0DvPbjsiA3
9o3b32HokCF7Rc1o7diNz9kaLgWpIPcVbDSFIQ9y2ayha/jszk2R+oOGzLq0rXdcQl6Sl97qewbf
yWmPH3YrxzLNiSK3TOeirBHMGZ/GljXZBlLQmhyudJ3VdvUuj8bHV0Ft4JsTqFHZorxqP1xS7MV2
76ZuDU3itmjFGYURfuhoHn9gdcE4AgabApCfDFfFxPoVLJuXqSxBVDpdp9oPg6/Y6ic42rulXk6j
L439osmmp7lQeSwly94CDMKSyv/I+KyGGrIQv9ovxlPLaUfGK9lXDf9yELGcQs0F7pdakEzRrpBZ
KQY/p0eOE+lCCKvwOIy7bSZOtiVZRoWMtTSjIyIJ1uvjbWRR07Dm5v6rpsbr8dQToCk94EWoarTF
ezOpTohq+M2DGvlaJDbZxsyM2poMAvfMWTMqPP7HO4cazL44Ue7ocu/OPQnKqZW4A9i50bNtddEa
tSrrBBcOSflaenVEJYvYbObiFrUYLFUVNWKLB4MwdHrv39kM4twDvSpM1VqFWVTahnOk3RHbri7B
BsIj8NliCZbKMMYf4mbJifYqxliOwO5/ckIDDSN8u51WUw5dCU/JDO8M4aELcsObYsrkKJjzTDft
ZYB6svXgL5zk9KEtVmyQZlyjiG/LRmbWfqnDUCNuMZc9JkS2Ga8JL2jYOvBe2rDP/yL8TbMIUSLx
xvBQrkfAvkpNyc06OXnJ5pV97Jn2ZZR96HxZLqqxbzLum5TOS/RtF2hm0TDQujzSiXCcH6XAVzOH
yCjdnd0HbvNixybBbjnyoZ9UEwHcS7+Wf8bb8In8SDB0L6Z0DyAWLccIo2DUhjNC6q6uDrWnCO/Q
899FQoOEU/u18Y1T6GimubyiibwGUicGsOLgZwtymrxCkDHhBMJVvLWVuR3q/0G0Qy8Uic5nLiCV
OGohAC4RWApkJDqKnuJdBehJ6EsNoxRlOzKm1CBrT6F3LJopWMT8RcIhAZFKVhDofnkc203dOVMI
/Q3eYZs4jDxPts5n66RLIegra2B36Pu1lB4yrfdYsNKSbP8iRFlF8bj6ZWEeYHGVmWvU5qaeatLW
86DCkChPt7AGwEUWdbl3GAt3FJVoCswAraD9e5vjGXYa44id3M6O48VRFnVvPqOlO6UI7Vbp9HoE
Bl0rd0nCFiUHNKAoMbsY/oXIRVbRMoYvtUfbx7aCAI5AFgjUhoBs20vIR1DLL8zQn6KST0DJSlfW
rc9yLqlZSQJo0PeYkcgvSAliCYRm5o/lltFOnqqNvHI5CyQswxgeV7LH/6py/2m1OULQkwtG3C2M
a3ATFutVsxYfnBinpfzyYruIf3jBNTa/eFdBICLeuno29Ixw7NGdYg7U5xbfLiTe2Ov6/s2GoH1j
BUN7gBfhB+GGk+NrIWRVVO+Lwetglj65NWC/bWj8dFj7qO1QMjeHHNP4PQauswD2TuyRTwtAb2QQ
lg04m9FfFAk7DINdwVlDCRWa/UZi5mLkrcok0rOdEJKxmKgI0GLa7T6bZ8GccvVAYFUlny22W0Xi
x3gNzTbwLafcS43uF+ppFn2zBiNTQGTFAXi8W8E1oDHBX+VWMJ/McbLUIjFOoPtDjUUUuIsan8Og
XRHwIoyqqZbkHtTXtNDi3Nu97WeBkzCkPttqSkvO9wPm5rRdPI8dV3FS/yNkgjgS2kJu3RDLV5t4
9AMwbfoge0zD+Yr/cKNjPv7CrQTJyEqw1MBhYlcZUM/8df4GF7SMiIzP7eKZIK7MA0vVzeQrpX3H
izs3bc+lVsf9M6wa+A7Wvh2Rtzc40kc1V+cNxCVC1mwgbARvJD0pFnc9NVKz5zBUHdfPLiEkCWl6
4fmBHdHYMW+BUEYX9Ij4zeA8fMWqKxc6shcAsGNJLv0X+dE2bnnUmrHJmcEsk/UX1NsN9YW4/dTY
EqLrx1fMzENu8YZ5/XbwEOPvf5CsB77Ez4SFG6RPnVvZktpldi1FZRR9HbtINEYE0GEmhThc3srm
zsEk5OxVLaXErNYXdtFqKPSTyEYWUih1lQoYxErS9IJbnqYzt5gz2SHTxER/q0qMLGKqkcavbniP
RZtW3f5NLu+CoDPJrtqUIDz4fONoiugBtJlQjubiv4bJ17zH/6dqdMDaBjLW4gEHEurPVueRWhLa
CZVrMvH3iqJZP6ujiCNAFbgBx5rdyj5I7Qr+xlikDJO2tqRnaMEZm2VgGpQnbu9L4AZF6sl8XLkd
Wfu9B4F3xURVzofzNqw0TMypB0lLfU2+2nINehDKue4khIIPcYD/clyoo5MSMx7rldCQ8tTE+2Uc
dp1VqiIPz6GHJp+SYbv/IBT49AxUKY0LxvTR9S4qqiAFsayoGGr6iREE6OyFPjjkHuK1964Fh/pX
VViNlOTvzTGPm6SpEV66Z87budAONll8ojqucFrabKLVDazeTF+Mh6pj274qCi7uLyLc1TjesuiD
cqtxCQe/nmX5b5Sw7KzSAFhXNPxdP5ROomyn65487hwA8YbYvnfka/Xo9ZzQLIMVGMqZVcChNiq8
mHIbaBu1TXZRwCnIODIZQBe/jbGf2/keiJQQTrqLMDi0fg3YwUlpehw+f0ei/RLvgLZ8czTdCLCX
oI8gF1zJvTkdN9JccAi5M8u+Rmi9vtirttBCWw/S2abMIBY40E2Ws/fjLvhd76p0Ekx18OlpWeAX
P5G/66KI+/Rj0L6ZY7d8R3qPOtnFOLMbuBOJcfh9CVsJxNvz1WGB68oinPWtRQgpVpyGM0kE12pD
elotRyCbiRnVALWWJNm+0oJfMbN74VMFfXEpPpjRebvr/LwZ7ihCjl3NbqcMTGiKqGlMTJCD0LGE
htPDtSvvgI7c/YBNugXgI6uXwPTkR24qZf6PPOoS/4CUjSN779gs+9F47LxygUy2IEEG9wg2FUkL
tnmofvxaYHUriuoLUpKzAyUP00Y0SMf/Ygc+jDGljIIx05X0jYoOOFltTout7sJXKbr7bEOqGMY4
E7yJRrdIxW0Y1x7L1e7ur1u+f+LkTThMARtXJ2Soym/bm3hAuYaHYWCF/zhdwlog8L7y+Qf2B5DM
Lry8UX7oE30WieqC1SJvN+bcBHGcCM3jpEeyk+QwNJcslrIz2bGOBL4CDnGJeitTLoHHabYzPAmM
m2RFoRSiFqQmsov3PokMF5k43kWS2M598+ScEFuGn8PniqdrPsG6WaCvSFWw2MB1E8QhVUQG1/wJ
JzrU4XsBIjxHvDnZWOSqTMJYaAmhIZGPz6kEteELZ7SQ590l73XloZ/3yxalF1GXAkD0Y8LB9kzs
Oqqal8Tso0w//PD+ZKOCLj5ache8+jzV7W8nu+KvXbGn+Pjz77c4/6kI42jH1L4snayqXCdUNkQG
5uebpRJLLztLe0HbwpHUYfa56InQ33ceP/huW8xPzSN9VB1M0mEn167Q/NPKf7kzobcuxIG6STl5
u8QnD4YYLd20R7ohv5hZa2D4+DurAXSwfaD8imTMqlprHYzWJ3Tit4KJvIMQ6QnJcj8tPvoGU0S5
oabXV5TDmRok6Tim7cTN+Vb149BHF9Gt5a6z0GW6/MmcV59dDxgnTVlkf/KUadFLm7eoEch+BmU+
uqMI1/Tn1ALvfC+kUnlsgcPRXz4DXHnUJCLbnnbLSLUt/HRZF0I0aoZjuSt3CLn9qQ8UAuHCfoVN
6yhlhghUZF6SYgaKWEQx55TzPQLD/q99Nhk299+Ed2OaccuSEVPB+/nLux3JZMqLBk5q/1Ffq2OV
fFA5sg+/nPbVPFUwhq9epsmXFPguDqsOjj8hR8kWzHXkKMpbctrkxhEr2TrYD+XPmBQzY/CwhZGz
KX/siucDFMlNnVLl/uWuIVFOzZyCvmyPpk00OgcWNQBb4u+V2QycPJ7IjXlB/RQsFMi2hreBoPrk
hPKynDupP1BXZwkev3jtUOLGflVykNg0j5SB7b5L2QZ/fb5cNpMnPAcjZfl5jQkaBIvmUBShzJJs
DXul4d5cQCJO83r3mBaucDlG6A7DdOY7HA2cVSHhOvj6YsqwltVpFEQN3+DxgTF72v3EqYEC1JIT
U0IzvjomcBe+1pt2a35PHYNc7FZvoxftayKVKNJTywt9Nkj22arx4Pt1lPpwogN6kePPFAryNOSC
tijrhgNwK+3Qq13RvHBHRuHAh3KZ2ih1okbO5T5HGZKzIAFAyCvukonR5lp0LPexO0g5v9QI1Xf8
3eqQOORvOWHt1HNQWGsv5Yvgt3tcd7JcLGpBiIcsCLi90glZXAA0JI1rGxDyVz9PnmJA/Mf9kdUX
HADLPrTgmcYfpyTvH2ZLrspM3heF0braoKbt2GpqjtZVD2oTDS0crddScHJBfvUEB5gm11+RDdg7
QhLJVAJBl6blVBBspKG4Q4w3GuT/Ynlew84Q6neFLjPOymW6KM2Qs7KYY813UKKxqQ+bYG2VFwwM
KF3k/EH7qyudv/0prlJ14CuYSkBwaVX+xtOB8INuf0az8SOHtznsOFIUu8Jq3fpLgQHuz4v3hFw6
PAU3R5hhen8hJUIPLCREOxCilsIMBLIYbKGLlKaPnA8QS6HcMEP4Z0akmxdxGDpgNbO63MC1hryC
5uWE4nyfenHKk1jwyGyrAmEUCvXC24dBgeKT612q5zTlpTG66MzRk63eLt7jB4GAdzVpWuTtFA0C
o7OyOAIgx3EVCIYP6FIdrdo0yg78+JFnidl8E5jYMCjyvMLMVESo3+gE9RdYo4mjFp2qBzM+G0Tr
G2hrTtb8HnwgvX/KEeybwzFRfLmnuCyWUB8/j160DqLRZGntKJ6tx572VqRZieV+mL20wIroeZZ+
Y2RC06qNvlMT1fk0TZNH3HYC4+pnjp+nCLUaRXHoqwokfdsneSfZBePq13bUQwn9CbZlzN4PW4AD
j1dF6sTYRV/KP2sIj/bl7e/K4irZj+BMMds46NPZa2NCqn1DaJAADcnBgv5a3LJi9bQoE7mgF8m1
sZeYCYo8gZ6k7Jb0Zeu8EBbWKAUinL4DA/q1oslHA5Hz++ZSxhppI0HqN5w4nWPZdkIbKW9Xl5/A
bxvraMUzGUZUKYfhq3F3HtLGgdGj7kK4Wo1ocWelDdFWub7rDDz0b0J6UVv4nY/Db8ka2yNdNP4E
Lt4BwSWb1c+ljHV+8eVhco5w13M5F1rfo7EoMrBJg9jKnrllr+IpeK40hHJkiMEbOpkrcKi/ogEX
rYrxlkQ3XOagYeAOwJsqfdJmh+9oAkiLtdU0YluM+LUbt5zc+jSYOUxtoK6uTSrHkqEbCLX4ouOB
9nQDHmZ00C/MFWAT5O5BAm6sb1jdbsTG7wxvK4n6NTSI3oKMQrSxeP108TkOK/yRhp9edk7/E6Ch
qhzJrGZySfoBfixd0PYGqAtmmbTw9Wnj4jfeVq7CCYabT1egoTbuvrAWp0gclOzOwg2KcN/yeknR
N+bxXiimiVkP26biHa4Zo7AZa2GfHymfC1rZcUtcLKehroM8+H3FjIknDyzAuJmJrHZmYYbJlme8
oY0x5m2XoKsXIIzjbPDq+D2lkYaFodLlklIHmi0/217jDRcSkzLG4Se4gTfhPAss1Ho0sl/RyxiP
d2DYzQuPhpbkhe1MWquB//4zqXAz79twpWJyTWEntTIGz66HBfRxDBsCHRsljd+WqeBxTeZnIhGf
Fp+ckUZ29kCk69cF+fkLDB3ZqXTmLw6wJbxunr0T3rv8kxPnyJhaC7uNg9xbb+teU7wf4uSLui9A
q2b8vd8tnqD2kZ2wIgIIwTbXWYkYVPUG4e2OEXvuLPJduyZxR1bufze+ObUb8w/WSBsHxi2EkQ0k
KCEIGkWxJrV0szsjndKG++EYjpjRdJ7Mq7g9G3oxz2xb+S3/179RikShlKke8CkQLYkHakw76V2R
d8Dkl44xmnzcTmceUv4GCQk+bIBm+bmRYZ8qtaSekvqFzWLJVCzpGy8seHmTfLJSQnhy/NuL8GQk
myYPRt2s3pBZfalhkfo3CSuoektxZR86fukXs60LZeW516b9XkTSYhPPUkTakMcAgIFqvqmy+dFd
cc1oHor6LHXHo5+ywxQdsaENEIaFjWfVfGx1nVXeYAZg+bowh7Gv/Jh1EZR9gOQu/ndDHcF0MdY2
weu9Wy7RXCJ4SfHaHeDjxmqda7+yG3wx5QmsDFwmyoMaV9431e9CL7+MQsDVd8ac5Z2b2CKnASax
taFZho+ebgS9ttF0oDYJQv4vr8RCWmVsfTlN8KD8ovzVvSSBVHxCdmVYhtH1Xw/2NkgrnWqg//fl
jw7MfFFUDkBaHF2zcj2yjvVEc4Kthi80r7QWLYFmUeKM+zT1ghkuzG2YWRjaxtL5wsHo1lloS2Wq
as7PLpoBtaARy1IVsAKvnbObrltmA8mk7nWQhkgbORdprHBVkvZsyb7te1QjGhZJdKWSVethLX0o
73UsCf/7XwkM8GlGJ4To5Gj+6OMXRVHy3AcfdP0xp61wB+QrPXUQWSG1dX5MGmeSHJ3nIls/I/4n
fxLeamY3XMScPj5Vq/9lluemv2DRS3KSLQS7M6RrBEQzoyFFAu5ZHXf/meqRyXFD/zKEnXuOyZjT
lOcOLSfIrB6QZR+PzryGtXUjKVuT4cbqfxMjeQF6XZAuYJjMUa+RZvwDzzCrRI1PStLZbvug84+C
/AbT8IwtZv6xZfQ4QT4yytUt56ZrcHs6FKLXVbKI84LuhAWidcvoewlP/sz1Q8RX65TM0hWfyGIe
2q2PHuuc5gtP5S5ZqvXAP4I98wr+qKxF0Y8IuicshL+p8c8tcKijQlv0kUxybk1e/KtCGMaaegXK
NnyDohG6TMyhEk8HiD4btjTCxueUwpmWSU99BbDZ/d0v1UUb19s30W+iyPONDGRc0GDjMVsW8U2L
oNqdWYJW67Zuj0x4zj9Xf298YzII9wW6ruYcpJZhz+DR2mPzrtvpDDwOSPIr44BIJqoGE+VuERoX
/db1HO3qkJRw9k2kQ7l06nYcUP59Xxr4RJ8tEqW64T8PZFj+q5+Upp0q0ZGeuvUg6aLnk6IZ+MMU
8rTtGwrDhqzYmu4MS7rGJUnVr123fiJHcQXNqn+uPB8EF/ni4eLigsdq/0uA2pntkVtT9RybvDff
HJYXaVgGKECcCWm6PWk3d1h5oTwHb/cC/2EFboHZJNFLzbv+sBdtR6SNg+BqORHL7l5dp8fW8Jpi
TlrF9y9zGD+l5b2QuJwqVzeFqTIjBjx8fyA68p29HcHpwDDBj4UCofRfUZan3AO43GRsR2dC/4t1
Z+dW1eoBDLnKq3KFD1pv02b3Yf+q0Sov5wkgPE08JRudakfFIpFt+6/m65RXOtDHA0Sv9V1V2Uah
9OizHBCkDlxNjD6GnTh7V1H3Us3oMKFgihDukgqy9uvd9/HukcaAHJ+dzopJlqQ0RvLg35+vxmVY
0zW4lbzdUuU/jp/IUdTMXBQJR0ybaM49C4tSOJJoiz/xTFs8pEsgJOxYXGQ5Ufw8GaHfytsSy2DK
gWqTqM16iH80TFku57TO9rdrnMDmQsGHdt/YsR+h1l/UX7uBbUpHJ+F+v5cYzWSIwO4D6GufcSYe
oRuoxwAiEPQxArClj4ynZfasHX1ZmTTPUTQP6+O8vxcLyGYGndbZOphgadM3eExCLv4YwQxTq3DV
aEdkEgpIVhACVsDaaVyl3u5ljbobA/LZOJQhqGHdZ4eC5dDTrlCr25GbR3KpL+03KV80gZiYzLrC
k+Aw1yt+qUq1/DhAq+Jx8gf8ix3uH/T3cLorAP0rIG9U3ywuRaBy571djK9jj20H83JYYc2ECUzz
erUe77bMHWSIh25wNmljwr/r/4wRH9k1PC6XCy4q6HAYazCkyeIhDAu9vuDqqAnsMzKK/cv+3GJi
k3LLX8uV+0K9691KROM8bVvydlRaaAmEp1v7Hk97JLBJEtKOZmC8bFUbsbpLpx8T8///pLfKBltI
TdybhfEmpyFT221xV/JUj5i8eMcvIC0n7UhcpZT52mSo7lz3/AXqMe+/D80RWVeQTD7EBlav1XRu
17EHrxOV0PDEXLHqlJ+ui5jumPwMCDhxRX67vmJtD/8nZN6BFORTsbtYt11/Jigi7zPcKa6/ZFCl
6pBbHz99IstMEEBEie3QfNJbI/5LRlO1YEOKE1YZ0uLu2IybsgfPgcFhXSBMCfU0c0830rH95q7R
ewDBWxJS8uxrm21wRsanM/c3WsIU/fCZZAk5SYNBTj6OqFN/Erm+QQ5pD20GbUtY1T/8K+ajm4+1
qSZjxQdOo1e8rzgdY9Sg4VlY78UP49jA5+tUKZSf9Rc6ApfpC+SbHARAwgFZ/czy/ogkEupt7XAb
SKFUUwNADBT6dagdWRxC64jZsY7WfYCAizjkUXorfjFGZfsufkYRvaSbvcd8iwShYHug7o7iVbne
ea98pFzI1tntOXQil0sUG0vD196vk9mPaf2hlcSTusojBAG30TE12SrhPqbxrXXCP6bisG0cnpDV
IOO+zAWlRLFTLBrTtoLECM7mUBKf8NM1LRA8A1V4PsWSoo062rZ3jSsDZ7PEW/XFxfi+fcyHJ16f
gWWNt7HSaMRjvcEdkVjRaeeCmRWvapq7gNBaQfZ5iJUHW3Teo/uVESQkYUZ5BsnBH86CR0V4eRJT
cOXsmwlQML/I11g9auWgpivnbfBtjH+WZh4nlPF39iOMKQ9kaLU9wHNOavk+r5gR44Mg65fH5/X/
8clIK0Kvlfov6IRuHvUoFYtFT28IO+a5GpnNo86eWz6OnAsDmKP4o2/JZ4SVrwr0qmBXWA/brW51
z/6JkKYmj7kJbk4seajlYNunHjf0YWcMIO4ogkwu4l6d9kHgDg9Uy6OIaPfePzqKdzxjmm7I6QrS
d6Pc1AzW4gepPnRVveMDlUOHKTLbAmeBcIOONHLLfl7kJDn5ZG24sjD4FfTVwX5b9a0rCEyJhUrB
O8rAdapUsQC1uTx2Lqm+G+Cb8xdtB6cDZm2POuSG/eXwKWkjICpCGCshSEyxoIY9j7bAFJOtgYUm
2dmKc7Ejt3erfHK1Ix9turD1yK5+Iq6ao+m81/C6RSozMHHpMvN3UncuGu3NLHEIj1x8koE25Lic
wtA7jfSN6ZA19/37JkY32FjUcMK5EZdkSC//KVNLuGY+BjxWdhkcgYVse0R8Qv0+8+6dWGdUWfjx
7vSUBGtb4fobdZNKUiWdKdAdcQes+sbI0cydCMmM481fBELVIeN5XHXoA/CmL07ZcCCl2r3JGNhZ
5z2C/+qqSGUMLPhRLaQLdn2pTWe+5k+e6hNK3lx+/d+Ot20oXQVH2TveHZE7JZ6ft5irqLynePG8
E4yZsrqNhUGFvgokmTfP9GTNha2ldN9HoZS91h5/+CHwsWXDSqYq6kl6crXpk5rezpHaWkvQj2k3
2pIDyjYA8tbRQc1lC6i9SYDhT7MsvN9lm4cYmpDp1yV78oaCuqPz3hgHqAtwGCjjNGj/2/jlZmdR
frkDOoEvtdRyl6XMtWJ/sb7ZWEkvQy0zG/JX9cxEho38ZTgzqYyVkbBDpcF0U/1dX5NKDg5Is1kg
dWlafWREngGuT4wMrPpKUFijoA+E9EOopi79Vr+GaYnl7GagnOksxWrJ5wF24IaVSoKa7pINFxsI
sbjae2pNv2Mkk0odKgtSbdpXLBWV/iidteUcdtej55vrJEQnKK9xSg9c/wUNwb6YnheVghKGZ/IJ
FVovRzcPeWrxJz/y/yTqUrlrmTcRpZf1LndqKvok35bTlb1O1GygMW6NFF+YMH+IN/Yr+JZOVYoq
F38RuPvabQvx6/28INSWGnhW7o02eZGUci96S5Hk8Mnd4AtUiWIN0S9bLwvZRuTICw6NA8kY14V9
EFKRSvK+a694gF7zsuzYCFVV31bSSJ7lDD4CFL0dtpzbfzp6N+VuMR0WgWjI1zTlPpDfNkiwxglP
6nRzAyyb+eu9tqd4Gf39f2Sdp5KwevdNZArMwSmkgEW5qez2pDou1iVeYMfqFi+D4gO+UEOrLdBU
e1v730sJ0qmNbC6FhVsJA51hOQISFzcCuL0l7QmoKl7TrAjnJwo7MuMbe4ZE/1C0jGsSzH62sokd
lW7GbrH6D5M3G7jaSnnXTUM/ms7vpatvbyN/EuXbiA8Vq+2mo29MeY/3+YG/a44vzu/y4Qve0//G
VkVXdeXkinrxBzeeh7fyNZd/r7X/oJlYZW51digqJ3Crpob9YImvkyZzf00o9GOBeSsBJqS1cdbW
hfS02265P/MBivsU2eylc/SAd9Hiezi7cOvvpMEqmXjrtC1VKZWEqTkM5d2dD5Kis+DRT+sXq3DD
W3W4WRwcjLgMZlMSJ65Yq5K2I/8pZIVZRjDZ9FpqMq3rVWZCpui/KDfq9Madt3IK13nD0BeDmHqX
uyLopppqXVo3H3hFtdaDtECH0zmzPEGjptjljxNKzDfam2aIcRZmHwULi0PtXcHCvyYoNOxN1DOP
Uw6reo0ILsmGhtVo1HTpe2QNGTlqjrmmr/9qGpZJNUFzRsyJKR8zX5msnuEToArY/6n2oGovReeg
psbU2b6oeLyWcBhIavstVETIsBwlZiR3prpGyHPdYVqCDUj1HjL/S2WXFa8Edl1qP4+amV+goMog
g9xGQm95440Muo0fuLbndBn9qTmpFb+h7D2HoDw0i6+coFvonbIlaPdA7BQDsdg988XhGhSiRd7C
hPS/ZeFfCOJqhya6GjhatDAkT1+VbLjCnv03WeWdi0zMhx4c+M1UYFDxtsp3sxG1dh86OvybUaKH
oJB3jQ4P+/v+VuPDsKoo2IQih5B1W84fpqg8xYKhA7cipIzMo6+kphxqJVfmmRCxWQ0eeeN9xERT
KcsBLQigKsg956geer5CuHT8B0LfXSucGmW8Dqu4H/8OPFNo9zDHyH2KxzfcMk4IAeFskJDLMxv0
K6Fc8T04Qg6NatoH9Mnvlq/MbwbbHFydGF1EBpL4eFCgRFlSu8xdhY1+ronJBCLes6i1u3Y/UIAM
0kULDSN766xFr4CvDowc3y2CrWmX0kXJdGpfDHuXU06hH6ad8hPDKGmtuXAjYn4L8ZFar6uovyyd
A20PXnYSE5Heqno2SBV/f6GMAP2zyF/NNtq71i7GOFP5nx1c+66Ss+JYUgKlX2a++zJTuMNX/fwI
I4QYftvko1ItVfUEO9U9GZWw2oS6WhExxJi6lkl9ezN0xI9eAliI9zkpwN5qKTHJKkxydSncGfgg
J3Pp7SUNbr5cvHWmhV0Eiv7PrSFxkfqAaxbGBXk4/V9mqZi0rKJCA7L2+RQpDhOnBVoMMSbsvNr4
bYLgfpnVTqSLfs3gsN2dsV/jrDZFyfF7rmKsEE46Yo7V6UPANGqGw6kTDms1cMMq6igrBt2g0Tbn
XWddXDJ7Un+Qe1FutCZK/F9ztf5fHAV8UdmjboqbZbc5fLUcnHexo1d45hWvpop6oQQYop0O1vTp
9cSdjwLg3dPrF2H/jZyt52wTHWUcWmQ8jsuTaCrXxyMb78Zi7XHqoOg9QVmLvnbaHMON4oNw4SM2
/R0EwYcy4vVCQvvRnnksLDaCx+3nRdS2/9u0YF0wMBM+WSq0ClXgrKwrB/Y/B93xif8621IjPoio
Z9DUFhouL6yyrOJNysYj40JR/WbjFqaI0L388TIAY4V2EDrrGjQlc2KGx7o2rsOpli89GGGgrgCl
T0QWsqEDRiXmYk8F2cWNHpMXZfOdRjxIblnW+FTnuE6aU2byn2Jm2LoK4eti83DUtN7AdOU8cIJX
jER2gY9O9bKcfH+0MWbe7mx8agRyY/KwBgwYACXCRckshIwcddrvbVQ/8OoWRvDq71oDx7hQdCaa
tuUiITqhYWU2bgOEOSvV2RdSDu6TUv0+btIP8oQ4TnjHUuH4hZDmB4cZqePpS3+j7eISsDn07Xbt
f5MunpeTbNy/P0QJkoTeyAlxyjIHgwIqXfGWxMEfHG0SDSWNrpD3SU1dbMYUAxd/FuyWramABveb
QlDik4HuWSZDEE40xg9WQJbmutB4dm3fvLLp3EZuMfry/740iSpBh8skye+JBJ8CgDfS5g+qRchp
fUYle7zfZlTcJotxzqVQqSdkh5JXuB4Xm+mkShzx+pVAR+IiSt349VJ8l+hMa35Rr/qWxY5ONpZ+
muC+gYZ+Xv0nN3lZxQunREe4a74Qg6qTJoNZrF3WiKyLEyNCYXBZfVfVlUlNQ0ceoIX8vt0geMWH
0RNlesHo69oryXSaJss5uA71XdbuvSoJPZB8GU0OAPoBLIe5OLs/cXi4kJIybhJ9xFtYbnxnGbkv
SyniUN8fJtNwf8cJeNkEU2UjYro8xZZ2ZLPLrDacV4m+IYHPU2+9yu75uGFbbZxg18MxpnSZMyE2
1yTMelWjKe1RIY4xVTUYcOb5Az8rPtCIpntOcJSWcBe/PU6DYE5sQ8VU9YRmIFaoncZxCEBQJ0Sl
ylxXZhQwqrOt1jtawfCdaBSnsZy4WujGkrmi5Ys2TsOYkLpUuUzNtRGm+85kUREdd0FA+Lo3WmZ7
zOHvmrZpYqTt4yI9xk3aqTFvBTt8cvLlTCosQbdoPRBXJFYPSrNwaB9TTnk7ElPlIme2aOX+lyf0
MzkRiblDZHQ1YB1NQKU+1swyP/DB8zOPNs4aWb51bwgxr+sHn5sZVf+GZWjmeDFyU/Rqs+PI8suq
D2jbgDkJMqvgeiJhX1TIw0ICvHoKhqSyzWgNak7JJAaJoMDtjue/lgiv0CpsaHVKwwFX5brecDiZ
ATUD4UPeTQlCs1m/gK26J2jbQWJNP9i5RYVvXiDrCEGGqWBgHQjjCP8Fqo5rImC70Co1b56FnJBQ
xsxj8slROJtWIZGlBkwhicVqwRafsnd2CNkj3HVQ4FdlaQ4s7PNI7NIow9z5z17dp+G8TZYQraO7
XljnEh/W77JXpFcsbCEkZbpWoWQ7dvHokJLK8S2mi2ojiW09WDGvFPeqyGSNU1w/b/6LhEhCy9zZ
DRIJ/VSuUM12w4HmAK+JOi3l40PpYFaLdMMLoF22xAitQbG149LobxABlAQUbtqI6gEZnf8K0chh
3tmnThGUq24MgFHPO2GFeAsy9X+RSSpz47ZcYoCjxCOvaU5ccxn9fHET5hoOexkZ9Xdr8eBIDfLR
49JorU+uSQ4OU4OjHTz8+J5/QwQKwdYm1/e2fmYbIT5ECw5E/xjDcxzVYGVmL3YYawWt4/omuYQk
+LBSLyLerwB7lWzAzTcmK17qrVU0hxBVy3fJXtsLTvKzm/1fFN8BtV308RiYZvFxjgP0xT4fjvpx
+V2XphLK8iP0ncWsQdRykIoAuWTectPefpRyiLtFqQGTFH4rvoICtRYJ5MjuQYZ0ibXbGwzRLGsQ
SHIJ4HT1nk2SNs/HD9J5/assEtJewY3d7F7NTaitU7+u+EFmK+pakPWS+/nJG+pgzex4Rj8hhy2G
+x776rGFmPtY6ot2ekFAUBmEYHSFxGsXJ4xTF0IsHN55XiBg8GMROKYwekdaAbcxbRD6pAlyQj2E
ku+rtLE24fKxmg69JAi7zmOndElf3Gp/bENWlnTAvjCbYVzDN413NNZxFiY82eih5rxoR/Tqg17k
JDXH2Oc0vmzexv4tcdiE+ogkBvehabFl0PaLOEkSR6gsUyI2B373d9QFF9moUGgk/Gcbk+QOybi+
gHiPPb9Iu5WaFoVul8/lnO6LriDE7YyGfoh9beGG0uKMUW9w07JyvQGnMlU5yeWYGNgu0ZlgrMr6
IQ8rVuY/6wZQBqMt9HtVmP5+xNUK+b8RHIuQ3EtkHPe76JlO4FOdMLo9G26dM0NfWSmKUFe0CrSt
ShtaP872ECYpy9pfxKnJ8KYH2YgMS7t64pb84AO0WaM7lnQjxjxKLDHGGFCfFYV53uTYs5msqhBZ
GrMzMpH4LqLbDtcdB//BfkCY6flH/g4OI+Rzx0mkpnjVaewHNxcE1klcS+8Zh3l1fhLWGpuCyje4
Jm/vos0DHF11+MPaLmGUe34MPshZfYubhX8kg5BcZ3xcR9ZUmFKG3CcjcTVIr3cIHn8QAD4kfmrP
/qcjwiTr+vYwG+Fu1hfnqIiBoEE/7mLAbKdP+GyCYQmJQAGFscv43XKI1eu8+Gu6+FeCF/iE7wls
8/+Q4g84aB6GIIsjaZtYP8cDpk+0Wm4p/R+052Yo5X049cX1ecr1A5G4JhgFnMcdx+O60NJ1GNP6
lBqFUKMW3JQxumC9vjkoQfXMQ05tTxibTqKCy4MNO4/jQW9sBM8znt2r66xo9l2RI80E/mFj4V+y
+d55bXaswy6REqO4n+DMd3Ox6iljGpyMFQG+UEQsyiEUQm4lNOcswh48fYjEsrDq4uQgKSJUeMua
TtDfxvZ9sSbAagFnPqU7K3wjykIRRviqk8zr7BESca+J/McTaHTrhRaz2Gcl7EvJOR4/i5Aa67Hd
wktizOm4HEk7EWV7idjniVlBJFeBFdGSxJ00IT+lFXKFlXXAlYE8Q0mSvqpBe1r0nhRkTYiPA/Bv
twqLRHOzqqESOL2Ygg2el1hCqMo9oZ7V4xqcHeSLsyvQ165kNL9gk2vb/nVFxJ0N1XoYlAzsgHJU
IzoZQxWPi2D8FiAVscv9akQufTLddUNb85SCLSxpLbe9dRFTNSCP3tQdeHElfmI0dNDjSsjRH5j8
bFuVNKMRhqblwYHm7oYadCzRwuTrGewKtqb99WYUEUYXPyLaws1jNftH+tFCGIyD4hUVuC6t/CXd
NjQM4yPMaNWVDZXvTImO/AxIlQxyBQB9CdEwncsvUubwczM+imEhr83bn9Wpr6Q+DazRd+ut5gtm
5PfZFnzDKr38e8/Ansq7LCoWAyheB1MIhGfIfz6MLC/oTFcu8Sh2vyZ58/qdGlJRZgGQEyOQRsLX
DLJZ8MjyT8cBD6/pTFLDrCrf70wwBnGcoc0r6PFTss1mplYjoIEmOXht8nGN13GLPfW8GUzcaIYz
7nMQgTLQT81eeiVcPTvzHAlS5XS8Sfif/8KJ5VsgF2ikdC5JHbWGbR7iNLbPslz+7ZopAj3DR/l/
saIQ5YswMMqcjQkBjpdI8aNRI4tAotG3bgxtR1OxxgbnGTX65RxHoMF2jF+31+BE15q3hC3WCU7D
lai4WvCH9iCg5L7r1KHX4zUB3NgrFmp3ffWxQxSviy8xY9FjA7LrS8yPKGBO8SBBUg1WL2xG+yjj
YNe4LxiwHf64/6E+6DX7LFNpshQmgD18Dp8NbCtF0D+/x9KFvOEsAMAcjCG65QO+xv2mLYr9tFGi
EWXm9mXBX5XSe3cRonZMTbPdyFpuCa7iYv9iWgInddA/ur+vf/QbXkwuIQ3WREXToQ+e/uELC0Io
pSP6KO6g7dP1Yfs0/kyD3XUDUChQfN8guK+MKmcIClM8WrPyCD0+08NLNsjP+EX3OHgEpnjuM0Ob
ofPfCsdPTnjDq7e3ViLbLoTXHy5GgjyWK3K6ooF0fEHmxKAPkypPkUyligNPjtrz4JhhjuUTRPCV
3O6/lEhW28jB1QozCh/xEzL6CGY2/s0/0qCGhvz7Sm4zM34dxa5k/wY5XHLP+8ZAqYaaH4Utt3HF
5GaQLGdggP+LGoe5IfPZG/QN5lFcPFZ8ovsSJxWuQa0Q/8T0gf1IOxHMyLiMJXsyMlkbL9ftJXRq
ZunDYnMMBNNjSTJbSMjg480ecrziYemjn3Y5XAG2PUuesz7CKOehA2XFYbsNo1eukymcmK6ULOrT
PlfbfckDBoQrIcF19SFUfQkhYt1hxK6+pYq1S2B45iRHKfhZJrHltfCCHye1zEjTiPxP0qapGyR0
NC8z42Oig14X0TWNuhKZK+P9s6wDUrnZTQLc/zbDwhuXhkJzSikiTSm0fidGZigzHjjERuVlG0Ya
teVvxbL3Kq0hiefKrdmKszBY9liI/uBDdYsTgiFm2kQzukmrwWedcWwcATgMBnND1Wf7Vcb85D8r
9xO30hxeF+Kqg/cIDhHnNYnOFZ+rnsENof6tMD1zp+Iwv7z7H1TDkAH5JvqOA0zNcrI0NZp2/tvU
Pr4QBVm5giR3E3NLHtUDwSBGrkSxpxwN/2EURkGdcmE1LZpK8SJTqjCzshIzlH0ItXVnE0dIBkDU
rsx7tL1Y8oABsJ6snPCzzyOFPpiTC091F3QT//qgu2984JYiO/qtQW9GKXmcqN7KCRacggInPIaE
5ms7DYN7yaqoWG2esXP7KsyjV42U8I/6zo4GOg/kV74E1IM+1pEEYZ9wpMZr3j2pPBotAxVdfDVD
9aoahnXeKFn69YOLfMFvTdQeCMBSgEYNoXVMoMM3YMPEcFg4XVxpOVx0xLAuSRkqSRe+wBCKwlEz
1n5Itqca4AusZosIoO4+eWTaPzg5+7TEgniKTGz1R6DwsKd+KDyE25KfN4AIFLs0MjAbHFphO1wQ
qSWFJ/DYuczR2dmdGEUylq+k2n5KVpWUXqiBdLHYEdYrGDkb47eNxxjsmr//Wr0w6+kdtPtGhI/0
aL+Fr4HMGnoWIFMWx1SEL/7XcOuRdIonnmj91UoJF/sTdHmIc9bCscnZVwDMTSHQOk+1NVy4sDE4
GsotdCnWCkvgtgNePiQkEUccwo6L4mZU2jqRK7T1FOuXmGRVV65B2FTgYak41jgRJcSZSELEwGpW
uJ/8q20XYyFsoR+lXDeAZSjawWaqgfzSsYLFYZ2k9ww8vmTz0ojyI9MpyP4Y4rlFWgcaHiPFBNLY
4bJZGNoJHZqp7BtLcNLwk0hpDDsjTHiuW/FypGUhMEPg0krQV/c8g8KjxMo9bmYmyg7z/y/MJj6r
gkK9ox03unrGRA7NP1R24PAnxtQXrzOQpLFq39aXejISa5lsBUVu+FKrNKkZIsbLnusPN4tQnzGC
NIMAJwInZifD5idIQZ2ArXk7noV5da/4Grif/bffKxcX8ZPpRmh1nr0jeibNQCF53bpX/DfQjM0O
SyO8snffI81UvyPbIGrfh77uqBWkph2o5F7b13E6U/s69wdqWDr8hltW4eRRw08Y9Az7e9h3DhUu
rToH1jnCF0XnOMk/tXouEwvPaB3wSpbK+ms+IcnZXuMZAUXSkEIdBaxcqgoWeHASdMR9PwEpV1u2
rk9aVqn5r6Z4Cn6RpDq3ZUICjmD6wp6XYx6425R6lH9J58j7KkKxJ1iR0UKhjB9eWNef90O9jeDo
j9qIikoDxtpoOgu7x6PACELUoFR5jSSkHamOhoudaKZjreaQobQXaSxkhDXzSHdg6nuyZq+ud3h5
YLKIW8fPFqdTbSXyDWWglDr1TcIRXCp5emf9vRIpxx4wTHuE9/Xe+5Bn5XUFlzJJ31rDRwss6yjG
50b8QDC39WMyycKDzjgtT2WeQ6CXSJYHCBr1QUE/sbJWvA6qhqbcV651RZLnc2k2JPanxCMr14D5
SZQ+MaFZUkEeNOoYmB39lRQSWzKu6Jbzgp85shyoPEZSQ5uryLgLU+K5K8kzHCzf9FsVKBRA2k6w
KKpr2ASZZtS5J1kWsDdNm4UBdo1dWpTOZE7Z0/LQoyUnW48PUC/QIOB6RT/u912lGesmg0iNE7dY
2azeM6RZ8ODE+vGNRGLtkg7VpCzAyui/fEDJL4olAxFN5CIJDcnlw8iux/KoYtPbbcL/GzFJJGgK
vW29T/txxCLAiCwUajClprFZtsBIarPLfS9axbUmmNIy7lRM9WIuN48lC67sFZAoOQvG2mJiol3e
1E1ij2Jc938/YbgKRNmX+6PWZY+TJQSeHDtiYfwlXGjOUKlP5IlxY4VxUDCWQtY7CJwCXnrEVyWh
4Hl335StI70wOhsAHvYeTXONOY9jVwplds1v6wu0xSSNritXJiSGk/6oB5BLf5ORjpiy2CfOAkH8
sGfbRqDpFeiOsV3zgvac3Ew27vPW174y+GviefdNIycSDVy8pIK9hfSxviXIaTUu22trUjRsOtFK
UrBGwoIxv+c45p8Mqy3VuGys1TwmnO3Wcs/e/yqWl2Q1RTNBNUII0OEjnjMId2M0jRjJjA0FqGp3
IdsanfUdb+o40ZYR2LyzEzdwg3ZKm72inQ2oTNwhByKwwtgWdKxdfYVbtFP+G31AbsBo840cFTQn
zW77VFEXSs6YghkaRh2lsCqdZssnLOwiCoS+/5mB8CdL3HiGS92IH7rNhA12hJTcwOseUWVPi/Na
0ju7hoS90+ZUz938mF1yOw2k7TWUGHXsZLIX1FhymZeEi6ovByRBuRBcDA4WSrNTOE/lx/LhMTV4
0DZteNXbNJX7zrkDVyGTFI1fy9s5uTuWex4qTKsMtff0Itw3ChPxWeksid3lMThWPXgbBAaZhgpi
azajbYoN+UpAHn8CXURmc0cYY05p9l+Oa6qr0lBEtt9cAmmwmrgEhr3E0Qknvb03mJijQg731j49
IP3T4wKsGyrhNfvVnA6D8/AwNlv1qBtvkikk9+p5A/Sg+rwY4aPICvfN5t25Ma3wcBBMWBoRfBj+
iSOsa/P986A7339isLmcymwcOVXXuhHY0AbMDRicB3Xfpxixhn9Iw5CSm8Cf54wo4wlxD0JiP3gx
uuYWSsIsYqXjV43xxn1YTwxcydGFJHcKpIkanudmNq+Xa5ebGpwwvbeXy4XOPP4wO/K66RVmrm3c
Kshzu0PBaBT2gXK7vvz8zPYv+u+GtMUUm499BQlndhY6fhbbOKvW7o6PmpDLL+QsFhmzZanJQiK/
lqKtsLPryRkD1nsDB9zu7n6eCf1JVk2q8js8OEOUeAlGkVPRMJblOhdEPtSmFSU5CJXYA70QdJXO
JuGbY+p7Q4zUPFC4mgff4TL+HagMINotLHVeuovU9gN/CNapwMKDaE4L81Er08nqCvKuo6goQ+uq
Qge5QzSt0zOxsx41bKhsJUFpcKg6fGNUcBfIk3suq+H+5bPyq/FpP1qkvvxa6m+SLp6TXI4efry0
JI19Y+vEanmXWPUnLKVH38pnGf7jj6v6h8pzOoJTY9OVdRCh38ku4CPVRbHWeQzzcoASTX/oVUTj
5XW+JoVSbyCOKy8A42cZPWPKgKfb5Q7EWcQ3VIuPmswF53VoWPu1gLYQVkrkcFpmlgA3WNzgLyK/
IY057DW/Pzno/AgqjrO6Q/Lj2tRrWd5zEyTsLxHufVgm8UGp+zbJcJxy9/uNQC0OZt6mAElcjsAH
fTc21bqdPLLKJRrE2tZh0KSINFI6K0anAeVeCjqZVTBr/TMWmLRawmLvf5U7l69JrpWwq/+HM58Y
VbVIUbrlAoKB30zqQe1rxZ4bOW1Ab4yjjxYaFXchxbcaZvJYfnK4cvv3UwUTcm8bKk/PnA3+N/NF
iQzevsH0fS7vm3APDn7hzpqoU1C0ESoD9+Z5m1MNdJVfRmQ8x59pP0jjxusfyFIKmrkEeto9gxAG
e3IjWA/H1yHAhQDQg57ocryNNYkSN9nJYVUWTzBCfoS+FxNzkMweF7zTb3LQM5qPPVzQMVDXLQ1o
xpQDAqvVZ4lLWWAZ5mbNRY1B/v/eza/56w0ikcYyiUdauRWEEA95YuZ7ChTipS+IgGVW7i0PJ+hN
mq4Q72GNDeypkSnT/tJjSwiaFl4Y3Uvkg96LsdwjK7JbF/QrBitA9qJQwdqqZ6C5fN01BrAfMhBl
31+8yS50pdAia+Oljy9p4HXYejFbTN4B+s2TQOoRHaYp5Sp4bvkAdDTSLeogGXXzVuwk5hpCBH2P
50hjvrhajZT6Q90uAtD6+wWLy8DQR4tBVCWCW/L5YpxLD4qc2n3WHk9ecWnahuQXq1IX3hPeCE9D
tueIGvezW8tQl1HOVfSj33wCGIYDz6S+XXoiJwbtQZyL1U+vd6Jqw1QdawU+oNlWhvpLH9e5esXa
e5SzzBy/ub8BFKLhZVIQT2ckK9fITksU0eRY1hZ87VXP7ZrOgQwG2p8P+eiPm7NBRYk/pkQwGutH
qiDQRNTzR01mDF+b1ltygIwAxqwu39tIT2s02rByCp1Neewt0a1mq0rumlb8zARg4KBsGhjBfNto
JtKP0bDQObvfKKXAk0J+fDJxa5NZwBuuj2NeiLMyFcwEOZHEtn+WhReiBJiS9scaz+u0be/Xk5O5
nfN0OKw8Jeh1A80uFIKjUjAS28nPxaslEai5lZdx6Sw+4lJ9bhWCkG4X4E4znPfwpKYSFARPSjQA
Tl7BFREMIWzjZc/izD7IuiuQLSw4TqC+x0x8wOIC9UxywnTXoWYP+5TeESX8Peg/PqaysvNILLCx
bRnVFsiPPPK49gtCtTy+dc4x5fx/SAi7VXJi3Gpg0kYeKa4PvgQaaebeysIOfU9vArcUp0hCGkGx
dTyS6YqZ+lyN8Z8+BIJqud1PCabr7ZUSC1fZXGll4UbbHsIimJDixwdaqi59BvhaYv4kkygDwHmx
uEtV/jeJIw06LVQjMEsHdGnG7HYLSlsPqU7ULBMErxkQouaAi/FXCLDviCUbqmrTcQr2c+otzKPd
P4/AC/FmOBwvpFxZVX6ya/Taux27nFdyMQhu4ucgD76LPa26lp1J5pJ3IBbZFRlDZhWQqI6ENla2
q1TMZiYaxFIy976oL1Wk7qmFlHKGna+mmjf0CiFiGMDwkf/R3Q91uCSr7LazfgTUTn7bg0U+5Ocj
rCBGKOUeeutMnve86FlZyPmEcLEJrLFV9kbXpfo0qwPdfRiTPCvhXL0lXZj5HSGVCcOWee83qEsC
IgHOcyh8eDxpb7h7RNIf3fn3c6syE5bwtMKTgl7+toI5riFQTauiB55tjNKN45inPVNPoDBHjSyv
hG/FHLVsNDQBWGP+S4mnTo0bL7t7vPygiVeP0bHpG+mjRX74UuuUznItMFjKxnQwBsc1ooMm/G1t
TY9/t1ckP3V35S7/LZgBeKOZVHIjbmFBs0ynSYhSKmcyiYAQQrKGYYePvDfgsUNyL1hIm8YFBUc8
8To3iTdWfuMqKw6b3WJufMc4Pw0/G/Dpd0epu5DTNPScLahQCuvKq1+vxVQgQ1hklach52aQlscj
VlDHn73+IdK+RtfB6qUWmliEcSqTOPvaEW1JKky4l4IKzlfJip0cFc6zBMtFUfZJhKR6TONSGnZC
N3JnYsOh+BqzZ7vJRsQ5MjXCo5NIOoN21SldMX7x1C85Y2J/CbMZHI9jha00IcM819U4LQCVKrT8
2AYsEXCnR7tBBi3BsQXIaFQFNHro33v6R/Imsf9yJQg39MBBhPpvoCv5xkSR5t1WweV/UuarUVM0
RXc6LSooyozD0nECdtcTUfUOqdD5Kt657AVb8YkWQHfRrTST4YC1gAI1WgNokOFEjD9QBcV+5BNq
PHmCRRLiD8IAyIjpwqcDr++8eg7AcUAfFO0LvH8SrTS6RcoFuz5jUHpk+cYEzy4m6UwhJbt84Pxr
keIUUhXJA98zyiVKpdjEOiRaQs05MGqkJeRK5B3hhYieMj4/YUWvC4GX+1RyCKpHyGiS7yf3Cerr
gMGKScimmXiq79JfzevLyEHBg+0B27r/M7Ydcn8EKsGj3HbtVYwhzxbMcczWIBGkYFVzKOUEOFVl
pJ4Grcu66Mm2y0V9SYRgI58FW4Ep5hLP1J9nyjdHtpPov3188lRaz2oBBgGxzKz75gCNwgWbneAt
ViypdwNFRAQtW8BP6rEe1OtCjmqnyEIUFOVAcFyNHwEAgy9CYSJXR2Hz/VcmVPWivl5tz4uIkXOT
yzS2G8ah68hNYmQ29Q3bUQjxZt8UuhvpBbeCPmEzFRycYBUO73xMD0OgqiglHryqbPNYWF0Ditqy
te62WnHPfJo7SNzLNFYz7bEmciw0GP9wzK3JoCkGL+ULwa/Bxqi+x/pZo1D4m9+CRz9WCclIT8qi
cqCPnz/33LLmkYgyA7iMZiqV8ijmTNVQ3CEz1t5D9BVY/9nJ7i+b50LGfmGQhDJTMGR6T+a7i8Pb
XJMlyWoTyr57VnHy7jDZeDWteBtWPzYuc02w1B/ewmR08QVm9uyKt9wouYuESJJ5FoE1l9F6QZ0h
psawxkejgZ1GeZTm8Z/0gdxJWf3MypX9wUKJ4Kh0OHj42hKxt08rtvlkEDn2w6TMYWJQzdwbh4Ry
uauXTwLk75nTCvmc5zQ1PwnMFWokJ0ZXF/GCqzPmSL0T3pEZy0vF0Gad3cTcVDyfDg+PXCywdQ8o
Ut1i04akodvn04Gr8khnQIIm3OF9umtbcn2yizYOQJtGIBBSNngi3OGYFFToog9IUghmegnUNkIT
sq8nvxGs3Z7xT1FhhIcpumv5mB5K2fH0lpqNestkKX4W8n/WEkNdpHUAdzBoggNTZ3mLnG7H2HEF
SdvoDMQ44/mqiUx+xSmq0spnZ0si9bS7s26WPRSINNM+ZyU4sqP+zKghkTWdGJSlklyO2kpeaMTq
Dx7zLjRAfSQf94JNVP6fffbDV92SqMwqIruERxBryM6aq8IKr4gwmr9ph8njzhIrVs79Sp+Kl799
5PEND+oh7HkmzjawbDJgn942MVQ7F0JhMOi1gpss+YlmYUAN+4F7B1vYZGgoL91ooTlyyCUb+U0s
CT3CfGZhNqqrI2DyBIsLNj0NtNqv7JOpkFcF4Jxn30BT1s/dAnIqMYWgUmasULzi/zxC5rwC7LtX
ueI8M9NH88d50o2GxS7gmhYkc1fAzwYgfpaQGH8JjOCClAezo9D02ODqB7KuMsKtHINHoAkHGY0/
/ZTvl9UoFlZNHTMB2FKyAunJOvK/g4HTjCZtYpiwPLh6OaT2hNDTc24A2i5dM2TgvO/pr9XaK4OU
t/tWKoYv4UkW69OEXdg29BVtD+QbLsy7PXlQ2OWj7tEv+XQK8Zk5dh+IGqQSlJ3OcE6FfNf+xAVV
hcGjdOP4g2ajj1fRq0YjPcAkfbyy5l3Yw3rMulE+5EjfB9KT0IfcJb9YcL17U0oKw6r8Z9xFianv
VqyVLvGdk5pBJ/VHIoxOwkN6gYEKp2iQvvNde0r6lHuVHZ+PVQIXKZCtTtXcpW/8B4hEGC0cNnY4
sOnrvAo55glBm0s3SXhoB1oHsdry92Yx83Y0wwZh+p2JWM3/c/+0eGR1BvtARvcaZP0Gh19zT+O0
rubnfvS/UHrAGcC97p8pt4fEfPWIS0YbXxjlpFXZYgMdu9+Vq27ptb19gPOEt2kgvjksAR4qa990
d4g3+zT4O1VfwZlWtKQSMXbRh+UcE8gXJ71bLKoN9h1BkNHD0Ppl0rQ65tmDbOShz6ZxxV+1LgVi
lAVpKQdORzpEx/4O0PrUzqt8CoEwmkoCPDlFUlyOx4r2DuSFkpK9uHOtoDodPc9xjZCDsy0LnnNm
aQ3UzixLRs8y2VwJtKfAcv0YcMUwd9kCNhmLdssKPa7lVJuD+mPyIwqCNIlNW1XeixY47g/tR+YZ
H41gNtmGSgdS5WSdIv4QFytx7rOrALDMvWCege3PUWix3FG159NCmQ+0EQEHeJ5DzNDfnPUr+4WO
c1JzYQSAQhLoU7eYnR+mmo4G1zUUhnSPnXN42aGa0EbXKZeKbUMAGWICLlstEb4hLfM37A3+4/D1
lGK7q38HUvYD6QTRhbjnbNpWyJ9FTPxZTQa8YYMXYRwGF6bg4akAHujuwzzH8ihr0b1KAEUwzSqL
KHqrhPq3e3t2xvbPN6qx7q1jVM9MNf9EWhd6hM8y+WcBv7kmeq+qHKj6nBRxXXsPm3L6wFucc369
MXmIaxjg68WJ4uo+gUb6Yaq7OmWGJthgI/tjv4r+fuM5OkiFviKP/8ueOT3NTbF7QEWghnHB3mvO
VjmxoyurRFEwr2cpM7pE1jaMb5zxPu66/RMN3K3i+XltHUVJEBt97IFuWcY3acbZ5+cxCy7XIe+l
eV5qPZIW7CDdbQP9NAwGNuX1rxj24bJThhj0WE1WppD7512jc0OyUIkUrgTrbGmmeFlNbhPHI3tB
bL+02lUv924tbY+wr/wOn1v6tRxLZG/uR8lWjqeWaQe0Ud1LOjzhhsNkmgIiBS2e6HwR1E7QjOhS
GaSJh1H66V8a0PXaorDr2GjDcEd3+wP5JNdtPdCsAFRFx9SKmkCS+B1/WLroiN6D/ZbLy1hDSHQ5
dz+hCHNHko87VWTgOdnZtMKW+qmJMF+RLy0udaSBsUmC9exkhs+1sQPV60PY2aC911lJVroRKyG5
KjF4tkN9uQ53nU65aDeAWIzGyDMpP46upl5uytUK1N2urqfJjTio3CCa/ayMCOVxKQOUHOxN5PeP
RTUThSgimcZbyCe+3wu1QotAmulG3mXJlsJoB8QW9QQYEDO0VB07Sr2Dhy+oClK+wZvtRt86odKF
J7WIbE5bquesk11gPj4W0vrLoxqVC4otGq60gywM0XjU8KPHm2jUn6rVZ38pU5NZdSaenp1e0K+B
1gw3jIkAJPuu72rV5AQlMGI1v1nnigiV7mlerJuSeEXjB6+QVum25WIkQMfn6mclRCG3V4uDrReU
KTSsP8nnGqP3g6TNT5Jv4VJ0zfBdLiQvOP3UfA9k626SZPv9eO8Tuq+sV6L6ECBpEESb4njAKLDK
86LLIuFqWnws79W+SgHPCedRWR1Kkh9EIYyDGKnLPmwoK9u47b94EgWkGYkq5gycw7sZssK768pr
E5ribDlBz3ZkjnIprmwb7EcNBUPWCc8fEJtf3qEXsa4K8cwabDC3ZYDMqa1xUcyuOpoDP7Tl/PvD
90t+7ZGYvTfKh44iyLUaZmIMVUdQ1cN+CX+2LIrdDr8ygJwOc7p09ccBDSFZpkar6YOF0+k6rONE
pB/HSNieLgq/ITMYp2hfzcmNi/cre7I2dN4gTqJ5tC6IzIbFJiaMnhsHeLSbMb2F/27F3h21iy9J
dGZaeyiAfq9o05lWt5FGw5Dgud0bO/cK3HQStzm9dclsCJR1pKxBMRYME/JX8ZA3x8BE6XlMnVTl
BNL4E/8H7XhsVijPILUBHOy8rQUYdTHSPIKQgvelTIwlEIhDwYOO4O7CHc2VrBcbg53YAQ2+wXwV
/WvIrby04Aqpykb0AfV9DGR2VfOQIyCECCabFi8CIAvNZt4f6SwYfOKE655O7BBUgKNpGQJuKSoQ
tw2ChLc6dSKWoijXipP8lTM/dA9qW4zQiTXhPcLWGpKpvUZohXJP4Sxux11IrAHQ2+6uVA+slRtn
MLQ6jBj7VmgQuxdMHxjfuMXWQ0KC5f58HcllnsxYQclbrWK4ZBT6XXAr48fUv+6Uwd5Tj3dx27Xx
8Yr1itsXZeed307FyN3b5YG/Yn58ihH9elnFTjBSWtrzuadqMo5wyVvF52aS3p+vz42THbP0rO52
sCC2eVrYUkJiFQu2TzPfrPMxnX9AWUsi+S2J/w/KL3HqKF8d+JPbWPm63aiojRiiJ6GXU4aqwcT4
MpBJfh6nSn0SenkE2hgFYJe0kLtzqfeWBAuRxHtiVF4y9Xw9A+RWrm2gmix1sbenQJjFj4uK/VVo
m7bghNfCDE9d72dgmFL13zrNBpquAkM74g4d7xGY3TiaIqecj95D8dniHTdd5V4IyBLI7rNe32+e
uR1EXsufgb9uAKXUcURcLUGbw7nUGHx1Kw0KQIMqdEfTSw7wz9ZSB8zK464HmbJx5Ffiwi7Wj4r0
tQM9MFVajUvXFXxbFvvjB2qXnwj8iJOEXdIul0W/FMZZ4JJ0yrc/hTiC9Jagyp63lZKsKIH7N6BX
U30+QdQt1OD1JlFj7/8ZF2QigXkHRl25ZJm+3upkrQ0hO+4573qWJ3XnEzsgbCDyoOgxYXXijlqI
wbafmcnQff0nbYv/B27yY5eCK4qkLK/o05ZOxzTHMvYxeLmo8oINxsOQw1sWc6JjBS8JRp8nynAp
AHzZFDut03RVLfRt4VN0iJBa0C7JF/CGxccAxqumUOB3EaqBJnmbi9ucQxGl3u7RGSfmtq8qNNyH
GY4dmxGEeBtUU12NA/qs1Qt+lv3EjNk3gJk6DSVRL1mtSwsfgOboGqpOjaipC//Iryp1UDIeM9EQ
ZRlWb4i3W4dhEQFDvaeON/GPa2Zp/fN7MYytEzhOCjhoCtY8fMoYhsOQMq4q4zDyZ/osSUCAl876
sdM2sjqiY8jDnbDxu9gDMqMuPda42xGvRWGTAJlBm5IZFCPvHKXbZP+fnR/Jpv/gL8rB28nkvkiN
32nkkiA77kgYsbNEcWJfIbXw3YCDqtECP7yB+TcyAbZwav5n7MF3O37rbLnmkLPmeS1S94+Xo/+y
wz94hDAgOMpjXg4dDJG6OzS7Fux+my+YzojsSCoQgSYa216nWQHCbEGMFkH7/wrEwR6aHX81vea8
IFa8Ij6+3vDKvEBDBQ9jh8vgDX8TgQOOK64jBjXl9FD9RSCUdkmHVxIoKuMH6eN3+3PaycWDZLsI
7cwz9dZWWn/5ndmeGaUqAtT2EQWXEAkSSZGPzuil+MRBZosJeIpwZXCj+J+gZ59siquf4MpZ3cxM
zYfRNI1UF5mFW7pxJJpWZCaunY/HQJskHckXCWcDi2TGyojEjjFGN2MidUvxVw1OJLgwNSteuZeS
UR38fjJAM7I2WOuR1GPx1bqq6P5c+cmiQsWVS5JmbsDgTWY5RTANwEFwd2qZ8S7d//aV+WkvpPEY
Z9hyh3Vt0IsRFpG+wZLuS6IYYORZwMo6sPCHtpUGOfOzDZNtlr3MhoaQpGolqb0ux9qLRQWbvvMR
+lz/MWDhn4x0kbhNGNvR8yMS2yaJkugBBDXxPciYDmkNLjupme6mHHvq8Hgv3rMUXoCZXFQ18XCz
GXRh7WeSTYIR45Q5RMDGQOebrMebpl3Ff/mo4M0BVcYsaGW8Pg8pumJoBCNr+jtnqYXONwpW19ER
C8A3OtMA83GcqcM1XQuXWmX4s1QmX9LnpLtqz8MQkpDydlIsVj+4ragFxm3dH0eMhZqp46NI9J7C
CFvQthhJ1zGxjoei3eTxdFaoVret6SdCUKgrPJ+8SbQ5yhxMUQBP7ys5kk+IUtjgWjwvsFpEn6AH
u/Ddp4ZcNH9T95inr3HoH1PvuDmypBFX+Dsj/J5Oai472pN11IdYAk8ji3qhRVag/R/P67WCgJ5w
0YeoqBGTZUUn56Cblvx5+MOpVUtQf/SeVr8E5VGAJuK8hY6x2N/ROr3+g5FwGC50V5mHiH+zrn1l
n1mEE0iv5wv3yrZCewaD7mhdWKIkQB8OA1kWt9MBoZ6Vfg7UBh0Rwr4zMUq7Jd+SV5CvmfNLaHN+
3lrJHmv5Yud+Bi8TkGOebavQDTaVMxaCOZg8oUSk0BGhSqRnr8sLxIi2vtp5HQSvE3fDw3MqDz0e
8Zn/NlkMgFLTuDvgimtw65VGxxzgpb9MZwiRbEqKe5/g96x190HZlgzGRe6O76GGyd/4kLcQTOWA
MD4pjq7WciqFlTlEU8frVK0cc4oZwp2TlA/QR7eU3vDBRTDAMZabuk98v8aCV5ffKNDy68WK/zyq
inSGEyQkE9M3UUFsff3mLGYOqvxy5kcrrws+RqBnxdb9WTCfgcQ0M53BJFZCjri01rkKdE0SS9Xd
SjO0GovZ8bWhag+nRzStNYzAydyavbV71MRuGIuDtnxledq5rvK/1TUfiBZo18HIP4UxP1BHmCdd
YE9GNXiImNvIDqlkQSDr1Qzw2k+23DMzsDcrwz7SClWkBu4tnB4Dv/02THLGB+saBSvUssxjeIF6
9nQxtdtU4UcWorv5VjRFOsDPArTKW44u5Gc7gBD9A7kbzTS1g5TfbHKZwqFVHzJe4Zw+VLNbuism
mlXTn6YLO6LTJ7SGrzn/SU0dPT5nPIb+ygI10govG8/rFskRQg0DXz+rPbHXhEoLIPUq7PGzAvzD
wyiX3n5ElC2DSc4ZhRQt3PliKeEVSlDxZf0v7dlL1u0rwqPUbY/gVEZwmqyyxZDHbgWj7PFn1L79
V3iNOTPuAiHfjyaUaCKlQCNFnTLOFj8+eF6LeYIom6K98xi+0R6XGmQegdeq2b4SDKcaWFwi/5ca
9K/VNasnlXIwmGAQKTv9SfDT498MjcY6Adwf5pSuAMmCnwH1lukKl0L57co2M+DOS4bBh8aGAiq2
8LNchfm0p/KTbLk7wEtRlED1Y+SJNhUUFhnKm+9DyOvEUisfKVpp+WLYcx+lPDpCRcZtCqdughnk
6jfd+ORVGzWU1I9Rx4Vdya+YFKHT+/Iy/yhA1hlpG1ZwUQKD8mIWULhMI68OrqGFc5lyxEamlxoU
Hu1xEQ/HhlktF643IGUbFtS+5vq2bN/eY44oBt5TawE8c1bYrtullnm+iQ/ytopaqwOj3NoX6Y3a
8W82+HNE7Xfv/ud7h7uPaxPg+lYl1RXyjxvpiVE2TZXmfGFZ1IaJotxTr3r5QUKpwikLH0eqLfKC
BgKcCQLbIKGn8joRE6DbTaGbAFr09PEPWX2SuIHKlEjgIZIEArEx3xSUcQ7kWUOYqK8tKSFQGDEg
vglPOVLNUyiHi23tF8G5+8C9IvKafAr7weZbbF8x2zuYkp9CE7uYeMiA7Tf7NRtUuNwoflZw/Plj
WkcoGpDMCYb+yVWYc5WKGsS3cwhbzI8cCkAB+P0zzuDltwqzKUat42xX7LYnfVcIFV2/NRmJDpfW
tPT5R/Uq7hDVEL/X0cxzvcd6XLZKI5P8Qp25yNgMwZZu1DT83XNNR+L7sfmq2ZheS9X0gU/Txeph
P23C7ONp2CqXBvlxugBN2zl7KPBw6QLWT28qvdUJro7chxRlHx8NxoJpVyE5xVRj7Bt4tY8mj8uj
Frka7GQIzZJFXm8YqmY7Lrp0arcZwAVoaV/WhW6kpO/EQ1jyjMOEd7lwS3gEWiklrUjyKPj7mV+Y
DYQaLHkAvJQKGUQaT9gbnM0Il+E6vCdzHhHfdBPFpvhj31HyTfEiRoAb8V/5MIGey+O6n2Vi7gO6
5Z0LE/3ko02Sqadf+jp7idLLZt/v2fgLYfsKOAcwo13247ExoiyOSMral2zNkZWJHOtuKz568SFJ
9LhPbOoiZs8UlKK6YftdQqMcYT+hbh42bH5g/RDY14cJf3Il6R0BUfmG6N6clbWtOkKvPshcC5Ea
gUu2sVA2FBzv3ObEWM7qV+XzdVQKDf9w2lcJMP25EK7w4wYnUnZkDBk8b/7DED4W44q4FeuGvPqN
72jyhHMK5JrGRl/W2LEjLQMdrCIZB+4hP9oz+n7G37DLBXgvuUNFLCbA1itj7sQUZ63QEFAlg217
JRT58wK7p34ZmVZm6Uw1chCBY9H+8dWpTa4qv4nHO20PpIlELvWLZ+hPaanbp7UoIOWeaBExeAiJ
47WObZ1HQru6h+jHbjgAvJj8/9BvM1/q4iiGDCnFs3cd+hPSRSoDZYruhrme3OSE501r/Xd9GwAC
yI6jhGWGUS4iPKlP2Blm3t1aQuIc6RBb9AN6TqrYHnPKxI1JY8dR1+wRRd9Fe7KMas+e3Ybc0v7/
40pzFjjMUSduM4r+SVnfd41eB/hIwuMxlbSBAKOfxGdko3DUm3Cw3uCFa653ag0HOi+E597fqj8R
Qn1Z0Is7+hgZP6aLT8JgdzEsF+LkXbjKKClr3kloXwmQ9PEj5/Hn4xtoFZ6heGy33Zwychn1R8hG
9lnI4GLMKMM7udNwSShyc8YAyqn5tEFn7K0zZFPr3ZbNW5fuD9z+z/DuF4cBe+QpbPf6cpRTQz2g
SKrrO+OU31giT+P61hFz3z2VytQP5AK2RwodNzHayKzlOgF3vokYYLlh9QqxGifCfC2ilBQ951MX
7VeOaDu+hHTcZGyPgzNj27gbtt6InnFvz65y+s+QVHp5o3XAS83ZXhCa97zV1vo8MT6iHJDcl2le
XmdKSDtFCK/xoe5+nIdGd2HoL3qtigvl/h2djr0OeFwcFWT4hRpQREwKuMnqRHmDP7aZtDbVlx3w
VSlPhAbOJZpa8aR4XyhVPDGm9CwGs9IDPynlAd0HIlj3es6nsG4vvp8E4eGnvkxfz6dKUk7v8mRb
8nbxo6F0Y1XHoxDxEeOqCDe/ABpUnOVPGooaVUdV0frz1a2zhPid4FCXbYu6i7i+ykr+JmIj76l4
QWOinxDWYR/zl40UutjpxI1cvkyieMtNCtrYVZYOKOJDzrKqELQx0D8/aKy8PNw6SITbT5HqVCRE
R3/o27jX4Yg+hl4jTp90UPzoRjhtPeSF7zybgZqusKTRUrC/lmrjffFPOOfSgM3YFAMi5YGF2K4F
s2HTTA+xTyJPGjXHJbKAbSrZhf5JN2vKrBApTSUo8D/7NIZctPvM15mFmCG8M9zO6rTdhqamB/rL
T7+M4SsrWEt+Apy7/ENdeBWOa45OkSoFt7N6VURtW+g6eVTAOweHX9xgRgbJ2NfD98/MlZhAiWWv
/MyoovCm7V22pUX3krlXxOd5HWcdpudrGX7UeszUtV1TVxjSz2Q9AIXjURBLsj34E548L0OkbGBO
Z0Eth2bjSPdFpNd1/LyqSqQ6oCEe1nUP68pvR9+BalD3lbmma0rsVCqjpCFBjPOcnOEORrY6Ynyw
ONYS+SSrHa1gK7fSNrobhNp/5FjBYCTHcT7nD7BbRZ+EV9ntW2hda5BmUlAP5lpQ6ssrpSBUrHyz
Ik16b5qh3NPCos6wRacd9N+F47XTgebdmhZyhz56pemMKxeRLQm7PPb5kBhNtxk36Vc2cboDVvW0
hOwV/g+8OmHxdXBtrPPv35F/2mN/ICIvwcNHvqS1wcoa266F5T49mJoQTHIUYu2Eluv98uWBIWvE
MbeniHyaq1KNo4q7XQIhG2hqZJMzQm2WZfJPOr5mwqbi/9nAqZXiVMt1Yi3m/M2BQw9z5w0bnjrg
9jQuM+wZDoK+ruLIXeazpGDgpcDxxPxuYbYhyp6wk1QojBJ5qB9FZE1iYTTyeuUK2DKkkF1bUof9
X/B5upkBmPCY00cu/O3+iQl5J7RBZ6E54lW8c7Le5VT3XJGRV26Neqmctdh6v/YUbYv1eP20BISh
XyLkAZ0BekWURHz9R2UPm3eASx1+LQZZgXjeyFmLzsvH+tFe//UgJPFfqwfySt6HmqGxAybNjTte
+K5haYuXxvgiJwfLgBqAIyNVNvwjXZwvfVW6pig7nbc96xIFcZh75s9UPB5tT/4TtlNkQQyZz4KM
eN1L7fXe6l+a6hcAySn62GpapIDM2IcJAOw0vOBwR0HzvYLFwIMEuwtLY7Xq4QzCWWiZHd89jjHj
++QUCcp1KR8wx0QFErJV1tINWzMzc87wIa6Lt2BDQGo6p+7ZFQzPBmfmfS8x9po79O8WkHTAuqfG
9O0rokyfHYxDePei5MHbPYHKF3+QHO7CatrrJPMfKoJtK+HwB3ITlGr4ql7bo8e1fQOD71gYKYsb
cD0J9MNLz7YfxH+ASX4TILBSc5DDhgwljic2BL7o/HVXzUbKKfOl1HfyJZ1e6VJxbMLneTExZyXP
tp+RbncyUNlOckH/BLNXuem3bVL01qyPhPyjhMCIiDSpVURPjxWmlcMBdwUPerTMDo4XuCHZFAub
ecDZT1cG3Wkdk6TzzCjkrzmwW453vwQ04jagU4N/+pi74bQ9+X07kei1aWdomRzb1vNOmCGmhQUk
/DNYSED2hcUzfvkA5nsxYem3X3vOFUE5jTXSF/EEhS6hfGc3YF67RuoqbqijjHVmDEjED6BeF9X5
H1an7oj5EqT8G8BGTlgfH/wF2Y3I3FZiYxEXpbV62YvDRT+BUNy1nv7j8FuWVMZZNalUE6Y8ZIte
8MaE3FFQpXKtKLMXILbIV2E6gNxUFgnssYW3xZyYbLhDP+m1hLGhQlrnSq9lnPTaMBTsRuZcQKDA
iXbWwPz2AF/A07p43+mOYgR7bjkJzq3XmMKvgi/K7tiUeStqJ34DNlTAqk6xfe5kozwln/ZBldHt
Id0izK2MjS9Vsp9zsCLQuYlDB1A19rRov4ysT84/gm0Hu36QkgTh8FyTAHkWUBiqDpYk7swykAnQ
Vz8OMgx0mbEWo9YGyLHq0iNTb5UefuebYu84m758MMuIRo2c941nsDbvvm6kLoonFRvXPq7SGCHB
dooIPv8/TnZkj/ZhE6BYR6ZsKugt3eYH+KDaOqoKYecIH9lQGwQCQ8p3fz/pk6QVpVyvc3wuvPgj
MnssawAiAMcQfoEIi3/ZF3w/px54DHPAvhcKwZngjd6Ib9n/nzES+yjn0pgcIvWw+obE6kVyi+RR
icG7uMJQFWyXO9aVAVwrdr1Bu+0nXUTxICfJGLHR3Ms9vOkDDIu107VJoTJMuDlMxZpvkTLW6aAb
oiC4yJ2sMbLPXc/xKC4PJkkcs3FoT0M2Xtkn765Me3TRW42iKFnVayG6R35yjHkUc1NtRlnTMSzV
YCjf+C1UJTDbnNG0bw7uB2D+kjYeU4SUia/JB0IYaHzszvWkPsWjVJsqBjZTUXlwANiqcRCbdAOT
yrvRlaSFKndnc1n2Laand396czyRXX/doFgZqp1akGZoKKFuN4HLe9nfgyIajNu6sIE7Y/VdHwMH
pEDniI8mVX0p+y+Ffg8sr+vVKaJuTOp3S8kPCcIEPKiHI5ktFup8/fjrs1bv+7Wh96FW/JtmvC3f
+B0k9Apt9sV0fYHGF6QbpHwp+9AaODaw7GeFFRSqbYGTt8sJ6cW6j35JTCnzw73dllLn5vwrqsef
DqLDfokpivhBOnSuQHkSSpQXILInvirTzes5UJr1WtauT3Xi0kQsqkCxlDQy3RZduVQNuzO+zS95
ZZ9XGa8Z2bgsW/qdzDqkMKjGhfLHMR5aB1VfKNApFnZvoFavLkdNJVOpN/x9WVcVFZ717bQWcVJm
FuPfLAziA4SepFGA7E7mPhs8HMCGj4TqD6RqvyK68ShG9tM3OegcqlFPtNjzVHTOmPhAG3GgyVYz
iBLgdmk+ZuahQRgYqXfBEDaudY8FthXAfrnlHmAVyxP1rJhSbBjlG2fFPJjCsTY1g+ydv5OQCWqx
5LYw1Xhi980T17erqGq6403gE2aACHhWbiQj2BJpDx2og7eyD5NmK8hmsX/8tO6rFe0GPWpmCg31
31N5matI148bWREcv0eUcRrZpIlYqZuZM78d1hVaZ5rurvEAG09+RJwVo1sXe65nEi37ffk2X+G5
9LE2GZozMCcgjVcq5QLhSKG74Tm6K13/+mEvmwDwC8ZFTn4NRyfo+eILnmXMMayaDe/GSp8SIbRp
w1tk1gOhVe2uIgPmt8sC8DvpUfW8I7wuX7eTmxo12Xe2Ib9eBpdashhZFmOLbhpldoasTHHrZX1H
LThGNazoywHCjA38evPC+LwGszNEBqb+7EKMNMWs+pJYnMOEmKlHBb2tEEfuDOvBfH5319fg3bYn
+pOmAn6xQM1in+zx9D3TCKNv0aXsf+aL2Ye2fNstZG7AdIkUse7Q82vFc9DHHG9V5l3JR+rM8iFT
9iWF8Y54Aub5fhtWLJbmEM+VCxucXdlISWK2vSF1u7ewdwQ32QsUikbWqvbeuKg2zPEmkosGmBpa
U6876Nx/P8CSr55bQHI06wyeO5XXG9i2Sdc4joH60M7Fje+hQc5kmVBnAV+1eyq744m37qSLUcG7
A7UFj33rHuj7YaiFN1LzKBB5VkWmflRz+XiVQHFqyrySWKCg4GRK48DyfzpD3t15IGHvsxhPOOPx
eH677erQsXt2sNQNsgrrUXv/3ZeW657TRshD0SuNBhazzhA8yr9raJbErBgD173FxbJrYXKEGZTs
/hwxciM1qIfDc0BnR5PHGY2NBEIF568Gts4OzottJ8jCUEYV9LeMyKxFy+OwOi4uoDWWpBxefVzG
9MG4lb/nCMEqm2hiXgNGKhyG2zO/ypuUFAKWEAhgZzAAHjgNatl+t7f0t7VnjIxReR5Rg7PAm8T8
FCw1GMFNMiDEsAG8edWzAIXd4vwT+75blGOdk1I1v7UgrYSxsDuzylFVJiQrf5ZHaXnxNGsW1MBJ
WMLyb+gJkTyvPM0tmqzlA3wiBt26B+VM/hXRRQOkRSMxuF7I0tp3TnAEDwFOCL7ohZvppMpPUzHY
I8TAC75m/FP8vL5CGVaD9CpBJ9ehyK/cnFy+T3ig/D9ZEeD2oJyQIgjRmdiM68Jt5EffxTYU8aRX
nZOCmJk3epX7XRVjz+vVB9+rKZPo1yCFgQOWHOHlJgWD5xczFBKXNPS0+lTo0Xk5jc6CoGH+NCHh
XzYtN3ovGV8b8KoC8vFO0ad8nHzsReCsKuU/iqGN60O6BPedOwkWYfKsR5VSnwIHL1PICXu8468V
dvFfzobJIZLgTJzskJ5JeIQ61t4J3uy1+BD1RkX4OYTZDYv97rihTMHr6YaMM9SYopoQmZ+xUaaj
0wXP9LkCse+sFiVtRZVBFZB87dPDfEqhhKfvcSs5vw1K0P+AM9VIFkFyH5dA/QH+V48hXUtH61eO
cKtNap+7t6yUHY5tqhhho2EHYSFImoWW/xWhaj2TX4kaeglyqxkOAgv+ZYPh0Y/X0yqsaEzTGHzM
e1zLVGldssPgQ3wpm4gzlCZE0EkQ5QtRJ21VafSrE9rpkDgQLUYhg01RMoib5m2icxMT7Ctq1EFy
gcguAk+Z3F0g1/n+KDUsaaCD+yw8G0TswcGCOeNXjgXjNKGe0IE1Q5Owq5z4wSlChi+gC4YjjDTS
yYWUFij6l/XT9xnWuGiVtFzI7CXMAdnzF1hEZ4X424mdHe/uRb71aH0OaaZpbAkaUVJJQXxCi3rX
7DcCqNwoLRmg/2YCdhEJNiz6tudm1UYM2tN0DTXK4bejv7Ud4kGPV7vNKqx9ub0Yn1jiXpysarFb
02/Ju1It0yMpzKx8vPIaQjJgEQyF/jq53Dssyoi3Mf7OhQ6/weerpUIr6jOFKGXBRFG46wSMuPCp
xCFM0B97gmF9pag2kztmA6LTAHR/eXwMGtWLUW0B2LsR9VdPa5MgtBRBHQ3MpMuQMHkVznfXrEj1
HMjvx+JuhqifVMN0V5Q5tC4uezasbk4z7+l5LkgtCzQSPAV7278SZmkFya1LhIAGfTcOEUUaDSfM
+kaFVomeIzAXXd+AWNXqrLQ4ANbjeYAXIjs29nK8q8ezKDK5u4TqT1qP5913nw2r+uz8a6AudgM2
NZy3YfHfj9UBFPZpu0Qa07kTDGSHSbzaQLLLx4O0Uy0DrFDmjF8n2QkG9Lr1bklkWXLL8RBueKAn
8BkopTRE5S6F1yCjZDUizJ3UL08rWibNPg1zDNTDqXYnuBwIwrN7JgW1rnqcuBgSC6W6/FCduvv6
6bFrVJxqtFvnRWqukPHnTAX5u/90+gk37vcySQ+I7TpfRv/i6n+uE8lLoSTk9g+xAsBeV4hNr9WQ
bVZinWF2JVtVftKikZ3mFCR+lhtO6AUTJSwFOgn+/CTntoHOq2PUG3QFfnMGxUP/vbA3h93r47bn
rCZhmbKYt370yRYiPzHmqduKzd3gC4nLQeos07OtiInLNhebR512iBpd8tVK+qCCtE64YYkEOSe3
HRxDqLbtn5V5oK3YgZHArzwElLPz/0NbqIxIHj63KJcBCglDWVvpjvixHUgYGAYqBE1K4tLsOsND
G8cvFpB8hNKH/2cDMNSXKZsSDwUqmy6Eo5WQxbhs6IQB6kruM1OqbBSLxI4++W4hYLhhVW0l1FAj
zkePY4DdmdJ4oArgNuelp0DqnLqltdyaJxYmRlLpmgR2Dy6LwS731qmOHjflKB8ElNaIOC4em4at
cLxtV9w6mrib+o6tZM59dQBnb2S491o+PSGTsD/RttBqcZdz26EFUr4uIC903/FDuQuD8sQfzHjS
1pH+O74xcAQwAieOwMRKCLRn04wd4r+pzf/fyJjhBXkY1zsEnlvUFP78q1GSpMrnFv1D8eEOpcka
FiX2jVWxeSMZ9SO5i/ANlMYIN5yj6wiLNLEqhExxtkWMFQrG6ZfTh9E3iS1BXzLtfzih+jdYDnYB
dPrLiw/UwMUYrO/xLD/j60Zr9GYT5vBxlH0X2chqdjKCaxtKz5Hi7dzGcCDXIKKoFJxLDhwh+nig
7RYDuf3K3NkUULW+OB6Isdnb2Fyg93Tfjv5deVfWNXR4582X0O/j+adJXmJA8Ks9fO6t9TRWqXAj
DCu9q9DRCpEkdNpK1Ar9CvQhqFJZYKuI8azCdMfttjRj8kJNfGKtMZdV6Rcu88m5vyb8SwgMHZPc
8f/r3rvYnFSYZGepd5ysZRKsbk8QMUnGv50wl+m3eX7ef/z7HkaS3q+jPTp0hRnFYWYjRAIs5go6
/rH/LDoBXZFYHpCj/89KMd/aIjvyTr1rt+9lFUwZBZLnjDlAzrNzm2M2yzR9dxoHZo0J6H6+xCw2
z3Wt72jlF7EQlVmj+FOUkgNl9iZORXp0x4rFduN+7OAZg1VbnxTRH885UUEPot8ts55D1yuTddyU
3BiBXcG8R1zEEvU2RFxu/Eznx+ijgqqmWCJ9JdG40at424HzhAQtdVbSlQFuHdHiQk+4jAL7pidt
VL1UIbsl4FsDcd/rgRhgdFR3J0bZ2INujOCOQfVM/iqqe3HM6OWVQVwIz8P4mPTAaYB9lUy9x4D1
bey3vXClhgd/BzLT/za4Dbr7NnF1mDjsK6ha7kTbZokbhz3kA3tWXiIVbfQ+E52GGL5kiPdgi9nE
04+csn4CKtpZWvGsy/enOYF9mhevCj3ViATnocBnL/zRfM+bHAhPRsXO9RZWJPJaenpBlOcPvnkr
Bt9s/DAkvcS5Kq2ilTPHEPfw7jYEA3mbM6Kwahyk3fLPMqEPHoLT3sfwPD6iQvvMnEkcrbjXM5Hm
r3gQi/eWx3VzMr3mpLy6qAcdz+gsAfSX2fKqaRnYmAaPYxrKc6yEEwv4ZqJbXzHf4SjCcJk3CZhZ
AiZ7liuwWnR2kQh/S2jPrryMFiRBtKBYHX9nb/D7gL8CYRDfJwj7ph+KTaTmuMIcY1MeoRo4FVhr
FcApQuE7VPN3p3z2rNagg+pcpfvAREpiTWcC4+SlYiiWTfeOpXkuCwMIWS41BESBoN5EhY4SitUn
Aiw9W3/ED6aaX2JK+1JXJetKqv1NbuS/qI6lyXdjExFN3FLFzZS9Vqlut+j9wxTs+K8ZJZsEs6AX
d1oaz8ShqTC1kmmtf1BsLpT8BdsTIbws0f9Xwa2CxWIDpaLLMFfopWo4w79Iz0FrB9jlRv2101Ur
ebAhFf5oZAygQS3Ridy2GIcKAwJNtBDcdaSqLOJph1mBF7o9f65cuB8F1yaFxBOytrMxHtrSlMy0
6G71cNiwr62bN981lMR54n8ajFU2Z5eyIXuIy2P7mxxaaHZiKhLiEGnBYCuGaMO9LVIIajUn+ZeM
fEAemBnWAwrnuHzrtTbZ12sXcBM6zQSubESpXALlhPIA9fhNatwBInuzX0AxnjVoR6rrQklWjPyT
ghSwog7NQeALcN0y/yMyHiU220zIcSossOcpGMYsY3VcSCA2hrLAfp6spQ/7nb/uIcBB3gh2UXDU
1IvPx7yJpRl/w9dcI1XoyFc+PcvAzUuNekOoyZKJ4YSrYK5vrwCD7jxeE8Os3SHiVy81CkukHq/I
usVQt+DSpMXQ8G2c2PgIMuu10pxzZYM97t9Ic/gTABD5nWNoehQJPz7JayCvRpqlbvjXGSOEk0KW
Dvgmft6prTAnud/AoH7tMpXPUIMcIxSUPU+d6nK5UhAfjHvcThtJd5t8mIfmkLvTTGjf7QroKaIS
MGe+lZ4uj4zbQeLgvWZ5Euez6KqBjpkYQo2hOuFha4XPsT86+r4KvP4a04E7ppy7r5qpNa548/Ml
T6sd9KTlH7bK1YEjMw/5a+0bvhN6juasEQGlfTGwGKdBNg9io1FZjs+DrERULLX4HPv3bxQ/x60H
M16EBQllHjoUJJmaSo5qOrJLGQsRQn05+0c04bTYgQJzBo/C8EMdQneyoXF2m1O6ED/4necdLm8x
cKRuPrXDsJMKAvzZc82eU3KFLed545w7TFiH4l/hHzdOBz6+5NGmBOnm/VS8ZBFTH6jhrtM4tMB5
gOES5+lkj285x06jjwoj90X56Ibp0LxKSeuuGtEi4f/ZM6paNkDIwnz7s6IfpIIUFHqObp6TDtvb
s1zho3N5RhksWWfxHMNHD3e9mTj3pjUpcsp9Jmm8Fx9T63609I9X1/EjFg/3rCElr3sZ9bCoW+sP
tHCIcS5t2BmVhoWPT/GQ8RY6Iq2q/W0LoUjxgyGAqqEAkBCXSABTEFkJFMJScmGp/StIiruKUceH
8SIKIQ6RhJQIZr5qMzPuLMo16NPUQn2Te4HVXFpuQTPOf8VpwZpHR4qRtIbBsDVRuhiqrDA9mj93
44fdRj0Fxq1AkLfsytg5bZdtVcJuFk1xFO4ZXZxbhpmNynuX9dTRu9bdJysNhc750I2ib5hWAIVB
cI8TmY77jy45+OqBrKC++4gqTHro2JSCX2KZQ4JWW/BN0JA4rIy0GZC7bW7qbTYA6F6yrGRD26uY
jXltXKb0IHK8PIZPQOimolCpHYk4W3zDqcCI5hZwrvGWYjes1lBulEn002kSkXswgiabfEMT3cYz
igMROl6oZiv54Z4IaDcgZ/SBpWo6N4EvTU3llZC50OO7USnxsWwh8Vc1Av/9XSYJK/6CoemT/TcL
MActGvXkzrU55I5vzSgWQ6SNBftbrIIvxMnubeAZ5XdhI2xLUnzP28dw7MjmuJGDYX9bflwXHTfN
WgfoVFaTYYbT+zdQtYCh21e64RqSFzUkpeirSChEx0JWgZhDz1Ty6FudYnW1ZFGWQ7TYhJYfkOiz
dEA5pMVsY1X1Vbmxwer8KXMEtr2cj/rVbZfBz5fJ5fV+ySOEzfQi9XvWSzojHGMbtec6eW8f6lm+
iZm/Yk+MHLzRiAhBNnDa7zyjGpmVOc3DgB9qGMXrbtOIDWUkoholxVawqSQTJAIOw1Fx47zC3Xek
DI00twdN5CQCfqTC4lc7g3CvCIH0KBWjYHOxWO7UiYrfjt1UbyT5E5h9lspGlXFk6jBn6LOfx2Nn
X6133xQhwRWe+hKwAgMPXWk/t8oSqz5pr/xXlRfaa89++3Ff1jzD+2I+xzwTJBw+J7YCo6nxKKkg
XuQmz4HgzXSahGoUZpthbGQe4HtY6hxppq/O/gOQZ0DlFTdIvuALZD27Tu7iyjvpWjb269yOWjJq
sUF+ogZDRDU6FfdtNn8QlQVO9HJDlDYqLuW9rgSLvapzoz3QuLAr+khaYwnoRUJIqF4DJsa3URG1
ZM6wcGqb+EjdS0mGP0TZSHcU5NAdS5Yo/q5VCJKwFW/KeoRYr0c6UVF+r3NNScopkSR0lWAv+kVu
olvb42D910+fs2kY4oSR+dtpUCORb3yhTRIoDyg4W+chCrRLzt7nYNkPHigooZcQ9eoyMmwVG2QQ
lS6mkM62yVmhEDXHFLoyvoVlyh8YiOslU5Y/Xp2eiH4biVaRw94dwfw1eLJ+IeTmUOzevyqjOCQ6
ACXQzPE5xNJYa6sYzpcBTQqVDceZPnVEqJFE6vStGhJQI8oND4Bgta1S+0TvDgdZ6KlQSXTV1tR6
CAHY5Dsy4vpsy3YNF6jPKgIS9Rv+GRSlW30wKqccExxepYT2WtTLkSrkosAXDuNuO9hijGlvDbRp
thUf2jCMEk3AFQ505hHOa77JEaJyPuQU+uR+/NDMB3lZtD5zR8/x+2K3uGo1hbR58q/VlUl3HjnL
+C+1Zsr30+0TQD78VGoLco0wGpTyVDa9BWjvWo9DAEEfDypX0U9y2ugQB9nSpD6v9aSA+ne7giiV
N84zm1qS5uRzGAZs1XEd2XwPEqxqyzAO0zY4o/j3LQ+IdtdgFUHEnnj+lZFLoRRnTiPSZfGkPy34
Lgvup1m9D8elUo1qDcoXE2izIXxv8eSwnY/qYqib0i4b71vSBVPrc9dqoQpVKDYz9oyDegluXio6
BGInzO45nxnbt8GshrqKDRdjfLvcgFhV/1uRgmkgn+RKszqhmVIND8EhkRCrhAYm1RvKq9W9GlKc
wC2JUwI0JFn70q+dlDvXasXcgLJZ0y/12HaOwnKE9IfcFAMFrr/ZBCXXGfIaMT5IKYRp3jZ7DFLm
P3lGyJoRYsOY/j1JB5xGjn2sKaMOcBDJH1QRyWVIStmfvgLQGYCfpFl+iwNHqrJ5TD6mSVZOzWR+
1zKut8pfhs9qiZ1TKFgOtjJmQA7yAV84FfRtjw5eQaJqe/AudQju3OKpSHgXkX5+Mh8mj+V8RuL1
KVH1iWDe657AQaJnKu6mWWR/vaaQQm3I0i6LiCTICT1qiWoocxC8HSpNF9v++0eCIXvAwurHuQ8v
z5AWRenN/wc4KYzBFscVD7Mn3l7pybFr3fNk9gjM0a1f5L8I7v2JMNGn68BGFn5ujv76TBRGfQ/S
AjFjgCBeuS8WiujKkccK0spHVbm2bfXrMQReWi2CUDRmaI7umcffHLHUsW0k2i5TXyobKb+yQHSD
WBsQKSYQouhnwhRUuWgvZM3FZ1Uwl/q4Q99ZF8B6uUR6uBDPuGtJqKQpXrZZH97As0Nj+EUlUDif
0OmQinaZkYpcZIjetC0c7dnFwYVuGJEZoo4qbk/lAioWMTadB+LSf50+mjL+bReL1B5y7EpWiIrZ
5hMTthjt6FW0Bdy4U0iO+iWm/10q9ych3CMRZD151/UjJKdZIrxNirKskHfZWY4T2MbkNZ1KcCMA
DU8I6y3FzR+O+JiV7tgQ6tl06bvmpJAFFlQl22y340a6K0FcesmQz5RiqSJxi8uG/H7lPu9vEYkO
zJ7cK6cmhPTwP+wJ8GR5TBe9sig3IR4hrIQwvlkFTnso+Ez6f17uLdO0wki2Tb5x8lJj3zeTqDD/
XrM5xbh4C8nmhJIEDkObRFL5mlnKvrkJb8a41yDGLEWEgL/miANX/riW7Lw5mHognQCcyMC94jXU
vy1dZHokv+lcZ8i/s2Pr+6sEmq2KBAMLS0eaWGxDVb6wu37BgBrkKPOY+HqtSTfXte2+Ihysdyiz
2mbiz7ugBqE2jnnNIlUtrYZEP29813KQqg/FvcAZOn4LcC764pnCRIpfBOGjjTJ+uDHqM3Pw0ov8
UffvB3KS2YFOHGF3Qi6CewS7lWI0OgUtz2jRTNibZB1PQO+zaFJhoSH/bqqOSHkkKBB5UTJMvTq4
tFhJaDgRnwAxFXTnB4EiolPid6WHMw0szcQUFJwnqrUYFSjz4Jruze7bb7Q9e9fG02SfPoaDX29v
fhPat46ajk4qpVvExnSLqTD6vtawJad+XjmrF4lTMNV1NYjvWKjZ8fy4+p9bqOCAdwjfuPqvpfcs
wmNzw/7N+FgVV6UiUl8G27XnFRuyW1Qo3kyLrRF303MIXo3lyJOo9ffr0JLMU4K23UTkC26U4Lyy
/ItJ2r5rSjwCxfHf212qWhpznE91Hrd4ce97DyTsJV2JgJf0Fubzg1Ni+8tY6EAFuq9ixAk/jhvc
LT3AFhJIgzMfY9zh4mCOaQVIVfSPp4K4QHy1QPNpLWPtdKVGL+Upz5/AtiNZYdu/mxeuJncQ3riR
V+MzR4xkn8ZshUBDJhJsnKvz5iVVon9iYsMbMIaLkACzVqGE6mKgQr6J98iyBtGCYeLeQnNg4kLN
ZfnouQd/Oly/uEC68p9F1Tp5Gx5DNDPy51I1JmT9/usWlEGOeso+2XPpzheqKA0mTGKK/qGlS0Qu
CEP2WZC0lB/4YzcTPph8daSikSYeFfTl2KT6iM72B6sjfDRHp7/PnaIUJYzI7onf05SUqE9hxbjS
O6UWrBBv+E8Mmu589Yu8BiDtaRvcbQcHzMdwBWyLjvRxDp04JDeglzQpgRTt6E+i7hjCGBEvyKnP
rKA5cqXakArB2CTf50OYvFCBrjr2Wsi3ByqqDBrwQG1J3oNsPwlZoJcy4WwfCE9TO331EtWch5ze
w6mYsHnSeAsujar42J2dElAk7u/q74soLYzqZuiBitELPXI1m6h1byIKSHLgJCJ9lhdp/FifIw81
TasNT41CWCkFZJegVG2pCTXijxONGK1YMSJl51xX2ka0zKfwA/QfSWmKh1E8bYkr2lOrJxj+BO1P
rLPIzLsPENPJ1vhmYlK493MZTbgMQN1RA0xMwl4l27N6qAqDobo0dUh3tL5KYkaxfJHefzcyboY8
tpDj9FLr5GKFGUpqYCe5cdFPpH6/3IxqyrbX1VNYJ0QCKlHN7EicRmxJzt9obQBubjbgOgX7Morf
6kRCGz6X/hRs9LDe8pIqHwtoP3Yh5/4If29e2MBSEXleiZ5Bh1e7BCWer0UQ9hwEuwF6G0eLY5/3
CvBtP6UeP0eBR/yoilINA4xmw/cakRnhIujzkJ8SticSiRUtfJXFuFU2tt4MB8z3ZrPSjuPbpgCB
bTDCFBltvjNL/CYzQs5RleQlrTHlzowI7z45uSc29Noa/5LSDwNio0RodDFMSwa9EN1FR5VkWO5m
kSrtsdCNO5AqxH5AwWzWx5zsjrejMgrluDNKI8XgmKDVc6bLfzO1GKdJ1DSYIGvFTKXJt5MpBKqF
1NYCQJOSbIMOSAAy/0LDhgWbrBrguUJZZHMnQ0UzYWSCqiYckvRlD7gpgmXg1PrAEUGPZDPHY6PU
bKL0xjGePrjJLPd3A6nrdweFgP+KPo/Er68zNoKDUhivCf08DGbEKVC9jj8yFq7tiDjLh1ABX85y
eNLjinVlVhlaqQEusHvGoMdWYGdxnvT8QRvKEASkbx+n5DXY/aagtaBigCYcpDBFhOuCBdKa/LBl
Gt6tLIT1xiSGkN6WgCcKWwA4QdjZZkNr/hY6TwxnrerOAN6Dfj3ny0mWG8BA+/8mtKsrtDQeg14P
hYtC+7DnvyfV3YOP91fiekHelJHtl/JnVmzdvukDLJHhr7ZWsmkBmVU3KxZlf4VNhw1dQQ/8PHmN
WyOqZCs9HcRkdqNxPZgzBvPv+P3FXngG93PvFpm9BYzJrK0B3ibx+igL6Q/STZ3EBaxJ1PSzOfzF
CQcgD0P+u85NfTQgXXWzknFjYXSDWrE+v4bh+GAERxuQsdfNchGVksmnS/auyWMiREwweHvMRUSr
k42wDTD3uXRka0PuXFziQwndF7CyRmQutgKaENfyhIRoXxBzw0yBWmCyYhlR6/1CfjjBXUSrxit9
o/eAoxiJNY4FDlEuwPdjnOsc25VyQdqsoeXi8IupPNPmv3uPFrTJt5EVbFN75cExFgxm4//eWDlX
cwY1S1DkWf8xQ5vce2GEwfKsYPviFYooQBKSxvO19Al3jY8WWApuQ5fdr+oIV0knWKNnxUh1GRsh
MEUFZP6Ru61RflUL/5AjlidjGKFUcZATEdGsdmIAmAskeZUIOqdPR8QV1JLl0scJV2jZZ5hCGC41
86UzmBGXQ2aPqKBeht1/ZWKJHX+aKeAzGiYQKiO6lCxzXQjP4eYCGM9tbF+dR1pJD39IF8lKFs/3
/NSAGnYABq/l39JCfXpVMrVJPGFMeKr8xw9KMOOhoeCMXljSOpWqmDi1LnSzI9sLvX/w+5OK7s9g
wqcc9NPUR7pMTKCjOtN6ipc7hBbNRQWQwMCWQrP8ADNxHZnD8DfalPZHwOwx8jCGn/IyCaqekadf
+rlKI6KOdvcScrUMEZFomKjQHo4iP+LKWedu/99p80lb+vxMFPOsvLe/lmWvaOuVLgNxV+TFbFAG
QAaZhy8eRJFlBlbVIhVSQfiOcZ3UtfTctIqsrRXr3b6lSEqHsEDU6XN5SXB6MeZb9Gzfib+vmmjC
dBrfneCTZvuQHzzMh94+FJwl2ATrzu25M93qWEmLzVQmpZEsI1ul8jfaJXypNcsqClm+dJJiVeCa
ludkdX0aPywo5WsXisV9W3Vfvla/VKhqOHYlFV+7Q1wVSR2/sVKmS6S/PYPcYq+au4dbrrWSbHQ+
Z9ClFtXwmDyMhxDN7Tcv7ScwKVl7FASdL900BhtQiVRHM3ubEIgC2eSGjLvADQDPR9yFU+Homgo8
H5qGtEgNhfMEbT70BcLrzpgT4DcxBxA+GofQ2FewEuOHdacHzy23ahDMF+qo35Nu8vGCF2uIg0m2
RdIFZpepf791YmVKOc08jeqbO4qq5YYZ2sb1B5PdGDraK80676yiS31zqppj8qpoPyBB9/aktmKH
DfsLHXCveW6ua6zj4MCkNSUij1pVWxQlVfXUzfnnnj031wTl3/KX1NUBDjTAhUsF5xav47A639yn
TJX7UeVLhPsjNgbByczOBn5ZPLfmiqQkT3qAdswNZWp4GzLEnRQukWvzaRHvba2BSRXaBpktxSfw
2sEohIpYEWXmW3Q9rnRwXVibyeMQGD85ltzHz3HyuXRE682H5cLMEP5GY53hI9xudXLGplSj9uXo
Hm34j5OzkbnqqYaxiSdwHCeFM2w15lJHoNScxYR0RIkMhXPg5iqObgZOD81WeuNJr0HmxfOuiUpa
8XInn4C092wD/ylA+Wt9U1BIDSKq5fI1QM0CzufHwuHkTEuuURwxLBXZ7H3CqfMS3f98UiGhEPjf
z2E6BgoRhb1LjzS8riKH5urnahKtkGB2hskCqUseYWMtuhZ9350rjwscSrD8jKrQMjFFfWDRYgtS
Id1LCUW/HzaBdkd6DB3sEmJWYDhEsR4RrWRQmcV/gCCOcSJdHqHMg4yFDI+BJ+GS1itcMjH4/ifP
MbceqQ6BZF+Hk4ya3xTzbvG7qO86Nhr4TJnQAej/+ZzdMzfwvVP+axb1qEaLFWN4/i4Wp7kSefGK
6Cqu1A5xFbMtfO1NGuary2G9zjMph5ndoa4ze5Y/u206veic+QBFzjHNNn3u/+HE2PTdT6pBXWZO
/NqfA2WqOeMoTyYTByVnNqg7YHgvBFwqvKL5sv246fVapjEZDJYXODetelN30HK9qUG0C0/HkOwH
mGxgU4mIAYqNPV3B0pTcx7Ky2xLQbpcuQdHDQr/N22fxMgVjdG5AH00lwehbYAJ94SHMKAXV+xna
Fix+g4x2bcWXJ4v4nrfhyFfpYhjdQXaBHpbVD7Al9hmtRLR0iargkGnNOAYV/IvuFLkVn4ve8omR
FQT2n7i+oeDVBAjbFZlP38xe0LlhCvjqA9J8/d78bI3MBKlhNFjP+2o+178D9JTDrEcwEDVKFcm7
dU+1jgcwij3jkO8C9r04pLVBskVYqIQ+y9bhjkOYcrs4GFJrvoq/34F09o/hgotpuY0HwRw/gI5E
uSWImNJyVUZo2SS+eIedQF0NQMY/NJRNdlk5MG/5MeN4G+ihTo2oPDMsp1HboCxrkjnyF0w9EOWF
IKBAkllHVBu0B4mcrxiyu2/whvvtHosD3zGyCkgzkpRVlB6AkiVxOkbvzVCkJnGVFBIr3vA6amyB
IdDnsN9bvLLZJdPP+4+sR5TM6sRckUUimg25mUjLncEf/KdBO0/387cePesNSn+oXLxFVIrCcT+0
zZRi2AWJQG8Nw/8Si5CRgqHM6merLLvCB2feS/rpXHFcsltRpSytLlCzcfk1fqfStBv5kOainOQa
cRA/l5wssAe0stV39NM5syyQaqa5QjcJOuXekitRmz2lRAjw1wg8Olg+HyO8kagAadCTXFSEeQJ2
7FttDKbgZfNWY6e9Ry/LSfEuPXEFJMX2vVFOUZAivq0QGvhS9LWv5RCk4ziRqUXsQOn6krHY6smP
o5wLK1iYTNCDrVxek+BXpEpT2rIypZLD35cAdlTbczoTibD5k8EH1sIzEjEcdSkt3iR/MdTK2DlZ
J806jppq/mNspCac/xs7DykhtPhIMmS0GixE+rGbV1A2DoVOObPEpX8sBZ6mR8NPNmfj9OKco6s6
soabsRSt3DezRbss6qYINyJS/9aRLhRQ6t392pUUIx8uqISjufU/hAyJnjNM6Ja9tXLCA80LPAmY
uPStVM4n7WkaecCTl+hj/c/59l6nmpXRRrdk5FMYsiyEY7+UP7+YSTztghk3wWyF4uK8tmTCbyWT
l3orZSg0N0nWwKOyuP3o/mdE1twE4uyaHMscMjFDqw1WqiDIRGBE16Kl5rugFW3yFiAhx1CgNZ4W
lMCZ4+gmYQyALmzsCg3LTQ19KwrOasMshX9KxgiEK6keAvo2KQTmzRO9FGLsLhQIFMQ1msVMApXL
b/eHYnOzQrQ6KinaZEoPhFD67ccHHnliss2jdcNEAKP69x1Mr1zLpzrYr7sedcKR3BPsgmGpG2sZ
+BID6FrdBUA9vyJIhwBvd+WkPMvUrC3Oj2rjv8uc/Fu44ewJeWIIMOlp2Js+7lUBcjJFkQi5RM+V
fv9BX6FcESKYeDieo6e1JgM4qWtNvLsz6QUmRfJO1T+vLW8ODKC093372pmrDIFwnpoh51NQS1D0
kkjGJwtcLwqqu+MXIK4eD2KnOpLv9kNoJzUMFBytAp9Am3aMlESLHccxGGg1g7NQkv6hiG1tGMId
Uz+P5SOOXlAAleMbfoI5OPNZ4zjMZGTeBBL0jZCl9OBFT5SrKmoMD2PAEczXlUutDfeatLum+j2B
iHlRqIouiHk9cuEVM9ImKqJvbzYniZRDLN9QOUSMKEELnN1sVGe0RbHw5ho6qYKjdDr3zFIMyQ6K
enXQzo91gTpXeBS7CSZRi1Dqo0PDnRhaQWJoEhm4hYBZyZdnGVljoDx/YgXgvEEFk9iSiZkuUpoH
fARxCMiZ78ghUGi7T4yi8R+P+QfdTwKRd6a8XeqM+Cc7jacbVeygo3/CRucXIqyeLmSoHgxRyc1K
41k2heAPbIo/VbQ888LpFUa4n3br/7PqGLyfTWXM/lrcXdK+pqgGcC90bCNgDe01Ko25pB2C/2ZF
HR7CtmHK0TvhaDhyRcN6Ng3yVpUyjKH5hvjuOFtjK++xfVoY9KG/KSwmsB0fpMZzyOwnu1bq+8wB
efxmtUgh2dTb1npBXZdJPtdK/CH6N/7Yafsjl81T9V8ILrt0p0/p7k7q4OE6zzY9wnr1FPBdVuEo
Xwn92eB1GMqCMzNfnGkYRFGAix6+gooO/WSX3AdvNTUscW/Qf69Y1y1a+fCd89N0scfsAc1Ck5rJ
dXSX8onbD/yRrGf1dnQiFhSyEc2VlCmbJL1rb24eSpxhoGZ89TudPeA3mIdUcAUbr4fiZtTA6ZL9
kWKSaUcrdEhpfv7XrDs/GP7gmCul3UxBc4leAfoTFck6qOwhu9cRGcXgdrIPqSx80VSAtD5GTi7J
INhiJ+k/L3WNamiQtbu+BGUSLrzmcarM1S/UQcs7VrD4sQwwKTnrhBM7MvmNC24JCk6BJnQ659Ph
lz+NmDT49zhYs7fvePjv5mlV/BSdAI51PW4Evu1hcrNmrl70X1DnUEnz3Ax33YBN3VjFzXykOVSb
VwhL4KDxSzu15Ze5OTfLiMZtko+ptt0ToEevRw6OPgsGSKG9crb9mTvFOaxyjlcf8f0JQAOR+CCJ
2NnWXaJU+M1mn+pmv61Gm/CIbnxxqzYAwgCeQ3OfzMNPUPTBW5go/ENYxImQs7OI3ItwX/9b83+B
WXXj1r0p9g75S54My0IbvmqXYB8LJifT5x9DSbgvFNGKBSeF/XtDjyxj0qenlTvFS9Rj87ZOzgwt
k1DRd7n7u6W/citnIhLInbJiIX+lZgPy2XbNC2sKijBJM6M6bV8eDBIilnLXtqydrlEoy14upSw2
CnKEJo34RaqFsu2laYh2FKD9asLD2furDtyxI6gdFQ8Tffy8DB+U12cvpbfbdcK+ucCtEO+s/GEv
jWWZ2Tcy+0miP/wyiiGNkHn15T1rZ4hHjcqw73K2We9TnqEqZy44ddBuPslh8+nPbUcNYL7Q1CfR
oSOZitVGylP3q2OrCYp9o7iDObVAd5c/P8wDSBI/E1Uc4hYIwlTRhuHUXr2oaQrq5SPlQJvfGFV1
LtWcWGbZSLeNFK8hsk8q+w57/08ImOQ9aD8c/gO+nFQKoHfQBnxY3ocf5/x/49lCWnHINbhAfstg
pqsSmebPhWh02aLppDMUL+F+TqKjeOJgUa4jUHMgx9jshY9sfvVmQGnZ/yOFODxcpQwbn0/VKtuH
I3dwwzNc+lNBmUyVa6nW3ypFzwT0UfrkfmiVEIqTx30+V4UmRd54iWJPeE5bohu4YvA6znW96kjJ
hPBubfDCfsfGcVoxkllnDDcG4Abgu7Wxmii6/lcsYG9+9330OV/8ILCWzaVJ9+6EwPbUP4bQ9lXt
4kENlVTZAfWxRDFbYBRwUzgqncxlwxIz4cRiUppYzVv75ZQkfpjNmh08tennXeDETqVJz5rF0H/W
al7nR7Y7n7sWrMWtYl6nWNTG1QUJVPMbabOZSk8dHTPzstdbEY9ngz1OkRlsdIKcojF1GYXix8Y9
N73NWeFF7Jt1OZjtBtldq5Ge7Wsb9c4PrqESHEaeJjTfHCSI6LpB34vdE67+wD7Yiz5ZzpW4Nj4k
V8JEPYyIKvVWu7KjxL5rtlZ+F+ZPy92949dP9BvxlPPDHHXOpYkg/nFmVf+CYYteMfq6jK8C8VBJ
6hs+caaGsC85fGl78dLKoVs1WQyGvy8RQmSnLrWO1HWg+azu8VQZ3Hs0rELs3fFFtLwA8VaoWoM5
vH3ERDRcewI5cNf/AhcbrW4SRHe0m1XSerYx07PPyejNO18W4tjvbghoSfqJYP8WyTNjDzb/+7Zo
dwQzgqAX7W3YbiLJjnMTUg8WUxJV5qsGgjYDmVKW6XzWBllPKU3opy0L7A8yLEkDKZ/OBZJQp7PJ
ckJADF5dnYhl/CkP3eyZcjqFVK/8Dhh9lGoCyeq/1LvEHknAiGSLZDNdVlz5jPPKo9fRIub8pAcA
mwSijOqVn3284+prrCXrs+f+8ro9mIGM3xL9+14RB9wccLL/kQ81Gge9BWedkg8UNZfSHp8GaZCy
31UkWT6fBpvPDgcNcGYa/E47qDjO3BxpxBUWt7ti2R6CoeKG+s8n5YetNVLBNALO5y1A8w8Yx89J
+ULTwY/+D9h5VoAeFEz0aobJli60zwAghvuE3GFzDa0N3CHHB9kdfnqXDENQzstdMuIflNCdGEZj
Q3khFQHmsj5hWKVrymqDaBfr4WkvH8Oy16NrUsOQr/Qj7fsNpZyL2c0Rj7Zr40dbg5+gJjBQapua
Zup4Q+R1760zez//A/bEF1wDO/FFVRZefBayftmsFjo0gmkTW/W/SgqBYEBYT1Rvl0q5iGY6r2fu
HJTJZBe43Btv4FQUADCU4gJPpTqfbGtFsSCPBbhE+/B7+nrnmb8P7k8zgbHrCcu4iGA/9ezsbXTm
FR42/jRVf1NrinfMk/7jebChREVIG8jEW0yXwHkj1Dtx77aBPyNmUTfIRokgA3uG8yAx43V+VBmr
eoxsvBTSZfgWw4KMaL5nLWYiwmAqU6A47+dYnSiIef9PsK1pfMtI/olFAlIN+Qu0kpFWHM7L4Epc
9Z7PNMRD8RZ/8PlMgEb7bWLdPlqH0UjRVEhc6vBnySeWLw9lShhHbH7NgAx4i41s9F7sL1b3PMG1
AHvdC6JSY9iV6UR4acyZ5UXG5Bi//sS0vaEqZd0HuK4HQ3MYMOrd7TXLhAxIlEOIXfANafNC8b3H
l+R5wC92znmDVMTDj2eCM3W+B1Qx3oUQ5w5yDeSs+hZdMYFkhLeARctVv84npPP+YA5GDz6OIxVO
PkFFlhVaju6YkrfiYAt+CrbfB4h50GmN7qDho6j8VCpaN/5nV+hicSoEST8s1WFhBFY8RMhywjI5
Jwx2HKbXt6e/Q4u4DaY4/kml0QgYYHKJLsYY4BCiOiOytQRx/8rK4144ntisF7IRFETgDEFrfCK8
Z/T3hSirgxs6cCVwaClDq5hT2ttXxW7LERvky5p3bs4Z03LW/N+cQYgLtdd3DWu7W6uLLKTlPqhK
2cxtrtAboaW7ai+8cOt56k6ttt+upTYw6DgBb2H3WvLKDSznu6Zm8rZ1/pnOQSfJC6xryR7hbDqs
hnPhRmd7Rdaov5Bi7sH1cS4TYrmAVLkg1kzatw2jwZ3zg//wu81DzNsqU9QjJxg/qAU7wscFQejh
w/PUBVPX79gbZ5pOsFl6rUz6q5kd2NiSntzweeRykfWGQZUPQR03COVQJ4wY9szbirKhvNLQiHTp
+FdaM7I0raMnoDU0+pj3of+PZf4kWI8Cb1qtQ0kKa4TiV3F17AQRWFGsdSSt2DbzjKJb3dDp8EJh
PK6Fw1A3LgH5f4r3q7MMjXI3jFFNlkR3euiHOMW1w/PJvhK8eR0/d7pCe37F9fW8ijityucq33UE
s1bBG4cH1tqjsbjFh9r4LP9+xdAKn4xql5rodfg0ypJWZoAGjh9l9gtgtUtUKqZVUGvn5SkeBy83
OsrYDwzIURInkogsWbQrqO408Dk+3gR8PNOuUbrz5l8F42iY5Gfi2WScVc6+xf/uS2w2Nbszr+rD
cnA/8FfwCJDaVnb8SrBobmmMhZMNETcVgKL3rBt6elepSQnsAcEDC40Y5onmxAdglXCx5pP7t55f
VUECoef1eOHkcDBn/qYfkQxXkJiEdgJqkTDSDcktK5gybPlKO9teO/mjRxNpA22w5Rt//0J3c0Pr
1MxevkLe/o1V4eSLlrExcXcHlZuYGLjAHyVM6iJf1jrRlD1uxwS0HTu9bgNqbSddGz/RaEjERMfg
tXhgtzrOiR6awmfUuE3GBqoL3hDyFyKqraJCyGR7dyU1qPGsieaqev3vcribN3Tesm+murwRi8ag
b2/oV3/7PpBpsJn7E18S44cTzwnqxmPRLG/taXkUEVxgJCxub1SrSUrbaQrItVcDlxwUviEU59C4
1o1JBLDMiQ4iNVm44Xgy+z0y0uuaPRC+UJ4EgAD/G2bGTsJwyqZ/JdnfGty+QBQSmXNZQzpgclYh
vXHvZ/Kruu5O42OdsfLXRdLE1TsJ2CFArAsBDQhmM6X6iZCEqDxFpF6wEemCWl0P4Zj9Z+XpzvoQ
cSrwtFDhWBdd/V26wLXEt38adKXcAIFnzFO2IUlYboXGqJpJfULFHYARvYy9QDJ5ZIgpY4/5e1Ah
H08AZSXNkWCzyfIpEMtY1Odsv+YiFNKMwho00c5IPQ/MFQa6Y40UFPCmOs+mOLN78psYYlpZGLiO
dsdrkh+MA6Iah4cWrYFCuHBD3yBYzDb6Py2AKLckWnnVbUf97Hq44LzLQD1X09y2VJETKqGDkiQS
ibhihuR90gZaYPTo8doDarZiIDIykqgHDzQtgVMhFMu6AYnfCEkdJE4r2RYef6dezp4fq/1Uzhg4
khA708hX4ujKW06dlh08o+HfJy7N+uDfMQv8yFf/BoyuB75n4ZFoK44do8Lou3K1PPhCZ1T6wyOe
hhZHmDDrnz45ss1YDuDZPgEy6zugfEUWtVd99jqhe6aCXNDkBiXIKFXjgRjpmbREevPvaOu3lfDs
/DZrQFxWHRPj48BWBzu0I3jRa2kgBnSTZx/baqiKUxHcwoZUVVRfx9T/cCxNegbTKlEDOkKJ4u8l
2cXQ4ZWSoNQjgL91X3mDR7NUDXmQ76Aj3f4yt5vr+ENZ9GEFMlXLIcWRJIaBWrZn+tQy+tXAhvuo
wh6RMUQqv/g7mXu2BRNKERRHIbjyD4AZDtZawXrJfsGycfPFKW4V8DeSkKJRFwUN1Xq7Jy7GlANj
Vrbdexr8JVdL1fEzuXnfIxLRPirJqQ9frzb/IieAMcN4GAuMzKWDACKyUhmzrd7SOQAZmyR4ED0V
NUV2W0b9kFD1nRhdiT8r+HFgzJr46GcHSSD81Da+Y55hTMfws0cMqQFWjrgrv8GLXgd2bP8hqu+l
gaqEYWfhbaKT/vdmywKjrvMA/Kv0IcGPWaj8G//3QpYv3hy1sVHDDbtYAlCxSRQsArE9pBzpGpsE
Cv/+RwPxifIQDjj/1Qu1DksZMvd9Vt1SMIUCxibwy3Pt/PGvSfeu6D3YjUGpX2grVV7/XTTL4veG
/chRlLMzPiqnwMQqy+ecjX9yk/RmgNC6xpW7wRzzAU1HbDjzC1QyTPba1I5q9iW81ra1KMgJpwfe
SozXuLezJ/aWT4Bhs8gIgYUCGmzmqfq2VVkueyBiYkHwY5c9ASP6/8VdYLGej0Au64lw8k/FC3Pa
oaPKEqFQcQ8Fd61W+uVyX7NFr/JzjODsHv7COvH2+gWI2N19s1+bFY3W137EbPZV23erHR/b6k2v
07Yq2H0MVJsuKWsaWd+7mo0acno2PbC6KCR9NRIgeeW3zZdK8XMm7rCRStOVgz62jlDNhth6caMu
CYYwl9DGMaopsVQdv33oSe1ChItvcqRKOQrpgItqPwaWc5BBunhISPoJAeVY3Xow4PEtRnUqU/kl
hMumxpdzcyxfK7bx9tzo5bTwfosazyubNrPM7/r+/plSQ4bzpMqsb4ytFpJP1//QHWiy4q0kFCr3
e59hJWyf93C3mp48NhD9W8ZzzhUQccc6D1FruHteOxhNJl2q19Bf3D4n9v8oOKFVVHVooJAgnmu8
efkjjyGe16PxEthHVxXFtaXwWi2oSofLFuKVh2ftjjOKM4gcOzWOl25FYBoW5eHnYYb6pgx+ibp6
2RQGdiyJLhE6QwJbDuaTbaJa7xpT/mL13OIfLSAeEwmCOcXnq7Axg7O3KeRIGW56rkY1HUUlDMYw
7u0b13nye5exyFfwM70JJLuj289lAGukAXSGaDJYWeI/nMVtgP3IdeMaVy4nBPvnP7rmi27wicIK
WdkE+BgEyge990lEUKVUm4NbtcY4jwDMcPE0GaooWcNn5VaxupUcM6FTtpB3DljD9UPjAErGKOEk
ncdclXc+x0RatHHfKE4D7LAuVgpO1S5IB7WQJ4Iq8G9hingfm1a+5p/qYaXn6N+Cz7+dV1XRss3x
XbTfQyBzFYqhuqKq0rl/F0yg1d3J/RSjfzqopwqwgv4w4Gvt5wd0IxzuJ6DlJ+Pyt28nPBYvr1vP
9h58xyJGPM0JuXl215P/fuVaZ31NvZm1rJkkBKEZcmrgUlpyYDzcscQFFE9C2fxy6BQguA60mXDi
W5Xz04/cC/9zhysDSx2vzEu4lL8lKTjBdGrXUHZYF8UlaatwAYWA9QKne+ywyo3HuPZlCmmTBiwW
YO6yI6OksIt7/55/KREYsT3lBTFdbkXeRtkOVDIqOsSzsqqguNn+wtBAPqlUwz9XoKowy+4+t1D0
3/DT8kz/Ntj8zhEYcyeJQNbGi1cefT6yHnt1KdJHRSfOBljONwA45le+KKeQ6udpXVwCXuORTfh+
hTYNXwMl7Nkdu1tU3X1LrFSIXVXvfN6FkLhABUywPNcg+Alq4otdupLcvYkHcOlTxS6+8+3yqDiX
UjiTrX9eDx1GyBvdCwcgEcLhapd8FhXwgALzEVszv8wMClNaUVAS/zLJXCn7JGSu7KcGI3iDRJa/
iBrbUpuMK0szd1vknr1SPxcvaXAaGxNTRTx+6t5bJ3/YNqGMjQe/53VOJovV1Q2gPCpXEG1A/XUD
JmNkPXjSNADMUaT98mhKXo3Oh4weOqNDvVgV5irAtP/bQU9uGBq0NOkj+BQWmTbFeboW2K10QnKB
l3qbuSL5JvuReepyq56Ed7r8YGChS3fJW1J0cfV5PEkwTSJW2fg5fr+cnlfI9ic5zZ3ZsqTaDqGn
3MkhzpX4kZUFMH8neZNNyM/1jsDVEQZX0xXaH8EguaJzN6kvavfQE31nd9JKfcxCdctIXE33njJL
plIynXfvvEQzho+3h1YG237Kgelv4/ScDm5z0f2eRGAaSogJISDlMzv8gdl3w25gePfF60zmNmTz
kkLcW+Kh5O1CV5u6OgcfdLV5ITgpucsIhrmNOr9tcyi+TljL+IzHr/wVuqiDF4kD/mgioPD3IXin
6qX7MWmSt8YuavKB1zaF3Xt89T2f2Ghzhij2XsKxbu4us7HGYfaImT/MyuD+YQZL8aOl4/QKkYlM
8UfFLhWN+lNc51T4AFjJrhe0Z8CkGtqRLzfqhQjOt8sqjScT2urf0T+Cql87j5+LtT5t84GGjnGd
AyaOzpvuMOt0jh2eMndZFvGaRk/2vQt9B0q1XTn0VTEJAzY/WIecsu8KXJbtOJWWkP8srZkQdQ7Z
QDpnuEfGm00h6iyExeJdBZg9U8QgUHshxwuuR9i4dhXHlhivnGytlnJzJJdrCHp8J03A7TLau2Xh
y2zaQxdQLTYtTFIK3KKwqhTNktDMWGVE4aINTkhkacNRrk4+WS6BVYmRsBG5BySX25nIilWwrGRy
D6519+0DVtbNX/aQTIkXfiIjUrk532vNTT0tQlI6Oq99SaWi1V+bQcOfaiiczIPp7qwEvip03/xJ
Z5J13IrG3Viqv64HmXAmsTDbqSQz/8WxPhlu6GJ/JvN6634x4e5bu05yxzA1+paf0onWuMsq3euj
Aq5t3nG1GoFmJvPkCLHsTTi9EXPNxEBKuJuEkpg+2ebNoeg0obyGxvnZh4fT4zW5Kh1xI2w6+gNt
Lq4UylhCWWOtsnhX1fMVaiTVdxe4zpdoXHhAvmSlytK+pqrwZdEu4/LVe6NbZwdBBf3lMQQ4/BtG
6Hn6wQlmSLWoQRZTxLAhsjzEkNymOgXRY6YnZNgAz67u7fmdPzpVz3qSKrZlWkEuZzoE1G9xNPSw
nF/FGEY2C382bi8s4hGL+rBMqpPCw1ZM9sAI12/tgdPUbhXqMWJCo+qiaJX3lHhI5YBwVKl47NwL
Gb7dGKnAobgP6znyxe9F4Xh2g7kCxCep7vsp31LGf7lAMXS2ybfb786Wfr+lACycu0gc9eVSfLaB
9UKGRLXt2gU3JXhGL70B67d3lGYWmM247ruz/07QPgiymfg1ZHX1doEMGQsGraLjU5aMnSy+v3Bt
hyARg7B0xZlHkJ+6Xz8jB1hecLsbsnhuSgbZt/b9dpvSR7961YcaQWoXW+pKLitWxTnF6XdJfkWJ
83uUyGfzsAeRxC1Pv86k4sypFRi9TAdzzNiryiSwe+4BqDHGf6MSx8dbQ51W5E02+tAO6IMsbHz0
jB7/Fy94b0bvUgHpVbID/5TwUAYsBRyj97NKqen1UzFIbAwZ3e8N1wBF+9nPUC9jAHXDS4sBP+eR
UT4jiVPfYP9fFlZHSV/0YuG5hJB6Bj962itAKZJN/G8rgVnfSLzB693LBWeGsx9xZl6o9qxaE3Su
nSFcRooUi5OcPFb2urmsNv/fl+t6vUjuwGC6dgQbz3xPqxuTQ2sJpwEo+XnWtz5hdX9Eq4BeRQby
A4GdAalh7BOqNypA1gWurUVBs6RsWB36q6Y5mN0GWK48Fy45sES9Z4Rv7LvniY+TmH59rlqBQJAv
VWw90uPv7muKFqmxRwZC/P1HDyl4bXV7xFUo8u1Ojc8zYqdkfvxUu/sqPLG2M6HLRpHWUPGRwKZz
vocOS5hxPCRUJ2SXoUSc1zr5c9CLTF4ohvpkRH8+ji76AlOstBvKAE4eu6qb1Ra8ED5n4edAS+vw
89jUp9NtiVyWAUqdfGvtHTdivYbd8GReIhW2dbtJGr9ECeenlt/lXa/SLejM5o85jwK95jHFUPze
nPcBPjNPNBSXsl7AcCb/YKJjf/M+wf5BWVQHm/l+l/J30IraekXgS5alZlcZu5SMQu8vt3n4ncTk
7cFTYi3sL7OYFbPfGkZm46A9VNEA36yru5Y3uLcH5wf/gO8TmM6oDZBq+6Rzb7VL2a6pH2MDx6zW
5jLLCd6pe1ssAi0TE1KcHwwGcRVHQj8St/NiR844FEHNLh7pC1AVAJPwjS8YHLhJe6HzZlURVn2b
ye71Ti6CyETRg3jFc0Fw+A0Apw1gdtj5i5zCVkeRMpin+ef4ULPyCullziIALJwYFB9w9w6cJCI/
BkG84d0U23gh+ksIbg/UPgNGQ2J2RnVqsa72Nj9aa/iz0duVL5Yu2PrZkO2UTkBNpj/xqMDEz3Kp
aRfgSxZqnNlaVsNnVwbMDXvT61PRnl/3sF5JSo+aaC0Vavm8ybHOkP2P+rB4RcoM5VcX9laPKIQ3
7b4LL+szjeZaJ7kpBbpnu813Vc9e3S9+/Kvcd4Ff7NcBdC1p0HcpIMHGNIY3dYnTa0pvzVFw+uCo
Vei7ZrIvpvZvcJ4TXurr9TjFunwTXcoAHFiPTdsXsalqw/g9Djjnt5/cVYKUIbjNmaLNOlfQxzsN
OS0I8iaKb+daEsbbdMEan4peX/BcJ5wm0ZWj1Y6dU2e42HlF6jbOwmTuArnru0+cMkGCkYNgxULl
8t+RlIvBbdfFAbs7yN6HoYNA2XTBrVOF3VJrkMbPVpOwvp7/uIGvWIADRF+c7KGefsYwZu+GWANH
jWiEbwiIn3zQ8MPuVKN2GQ6IAv51loG9SmL5qAebo0cnhC7ceqreZ2X79M8nkFLZUZErkmbeDG+n
4MeW8OrOKLeGmS1LUjqhQz1Us0pK8HaGa7iCBT9n9G0Cs+MnM+TivE4gtRWHUIr52GOl8enFs2np
8GTq91v/erkZZPJjTX+9ilcKHjPcmt99wdTsK4FiFu6gezS/3x7T1GxxjtMw4/w9I9oZ2qGKElm5
U14Mcj5t54ELAxzy8Nk3hpeUgVxtiYYsiRoQ6DWjA52HcED4BK7NOB0JglZY6ClioAQI5hjX03AV
R00QxOX4stNqJpTUAL2ukHigiWjcFoihKv6hG8eqiDwCoBWTTZlj5CBJJo7VrRjzlktupJTdBQjp
rHBGJmS2OpIP2xsq3WvBRGB+EsqfGhAE07vPf0qHN664mZOXgMr0YE64Ee8J5KymftHVDNJfF6I6
dB6AUDLprdJywe8+10Ev+V9C7GP7iQFSjpIonYHP/PAoSC1aL21O/Z95uoR9+kd3ZKkpgpzxEiIT
e5gxDVVE32GnxKtNRKmz8wLmv881NYpyOPpMXJ2IdAZmvfClaYrh3sJ/L7Q0Xzs4z7x8KMp43ZuE
yWclKkPVB0mrYXm8jYxERkb6HngRbxbhnrKGrRfG8u/A2gOjNRjixTPlrrCQt/5U2OmR6hL2hVo3
DWxUE1l7zeUV93tz2PGkqYy1fJKTRhnRV192JO3IWD9AX1TOBhIY1ALIbYrtRQooVvqNgtLByILD
GM3f+T25z25/3jns9C6NfUWjoF9TA8/U0syQmz0oB/HnCdbL9FC07sFsk/CA394y6cyuReCK/dYf
yungeD6k3rhsp0CC+i50A8f66SjSQSCtijrklEcIXFCdHwPq7wsVwmFK8/qZDOFeMgl7r8dJhMdE
VfUcdWfe5RqcdKij0MFmkPWbjZO1bYZIZS6uwZFgR4S6ByNUKSo/M3gUcb3NYgDKQOUmMfq++mLp
s6vgcDltBScZnqWZwzLXCdpB0ynDp7eJ0TaoCRP0jyTUZpuXxH8M4Kdi+50udWHHUzr3rOvhQuzh
Paywa9iZ3IWzhrfB67aT6NU5+gphjk0QVmZDoOqxp+5TwlBcQyWzvfrKUmYh6NwH0/Muuv5m2MyW
/ptdDlLlnxPIXVftYxijtG28s3lpaNydRayqgpUbendsdP2zs0TSKZSaYv6aAyjl6tRnf6CCgGCB
DH/Xhu99xoruby3EP3R9SN9HqsHxOfod+z3b6M9X1CS9gLK/DKeA1PbXy6HjXtWhVM5D8ii9TFe4
jUm5PWnzYwOko9ACgnPwH2oU2Y1ogWVMvpinBxlxNTsvivWuIloiTCDT/68Ruq8fkFAFSGwx6EAz
j/Bvem7PzZPBiBHAYG8A7LZZ0ZT76ipEL2WLBHMUZr+Rr3eJQUn8f9z1HyS3jz1ME0NC8LhJSquO
NUqqWopESb4rvTiYYsLNB9CMI291BP3oxt74zFp/RnHBI3yNVzZBIo3LpFem/9g7XXrPgqn1tpFm
xxoRPAGO6b+UmEF+a8v624LRumW9579UnYT/k3mjTJHbfzSNra/2itA+l+bduvrOJhMKKgmULW2q
BHuAlLctjQYa/tGepXYMH6RUa+AuQgrYYTAKU0Xouipmgkze17XtoT916diaM74W9iVxeXvzum/V
UexbxNxhplekh7n2pQUlTiF+B3p+qzimREH3TMQsQlHh52YvNQoiF1EktchkNNSZvFASsF+Yb62z
RobP/klVT1sXtQ/tRD31KXvMa3e275fgsVUmc2FF84M3zRTKuQqJOOrXAeUkDQwibjnpy6BfMmN6
n2i1sfi6Gq4yu+inrZFPYh4ur4gFCgX56pSNYXN3syRlj+8t+MNHChye0tMlqBfjAB2gc10G3fLd
4oUdP4iTEmdnlac+TzNY7elas30RYpJJSpjNd7/Jc7W9ytJt8VLwRamjpvdUcrqcKNDlV2dMmUYB
4L7yofH17s8SfwIHZ+9RUXN2D3TTzHKu9mJgvfIo12j3F/Zk5UohCuXj5dHGfzjZ+ZPHkxJCY4AL
sYNhU9Ygn9myYiBfqd23aQvntlOUw/Ts5EZBKvetJ4zNuCEvrWoVSbfQu8oDjOExm3hmDxs+YKUo
tpLjNOnIxtD336aUu2hm1X47l99ROL4gwrqqYI67OUFBBvOEIciTQLTEGUMfXRSbmhblFcCEiGUc
f9GrhyrDr7WvkfgzyF97JmPVbDpdUkCiz7r/2kCZv8YBoAHUU0mc2W5tXXGdhb+KxULMteaB0K5Q
RWJUlq8tL1qIhBcfak/b36eJ4kcmxCX5yk0TslsBvygJje+Yqpdmav91Dn7mUP/FdFQwqlZD+nuq
hYUsLjBHr4r3keY0M5+8N8ezeAL00j9v9s0B5AZp8bnXtYhzf2NQcPkTwVX0rcw7jjbDlFQxOD7R
u2e/IMge9FNcyeJ/PeXcHhnis0b+U47GlvzxG6vyvJv4QkAFM/UdIFjNGVEvbpRc2gmIyD3G7iQl
v/nGgeGqVZyoBGKAoPGpNvAhPhnrysi+TSIji/VltzHTMhgIHK7m1eOTbtXolQk0j0rFY/+jkAcJ
UEVy680nox8L2vMLU4IiyMGhBAmASyZoaG0qET27RBO3Ei1B/bub7FFLeTi0a7ozugp8jfGOJTtk
LkqrspA3PLFg5jzn2jLF5ZKxDJ+ytWUBW8GIhB7FFjwMcNUxrBuS/PsTjn1llfkgLN1S240WGBhY
ERpscyg6j8pouf6zGt4LczMYnmiLnHq1ZqaiMJS86nyElXWxoN12vhfjkjH4fapeVO27zgPT3O9L
Cute3ay4H4/rQanTE5Kv7A2DjDyY+e5Zm7mWFE+3UrScOu/Oha4Rz9RHSfgwCrV9TpvQ3jDvGFah
4sw/IHDRW35/D8WhmSj9rh9G+DXx5ir+bJ8dZY3Y96Ph5rktKHtR7JrEcYuxVcJS+JVNiKpNsY3V
N7OpPzFFpWBs0KwJm8459lztSodqaB9Q6afJrVKuAWFnWKB4Awy4RM7ybVjEe8KZwAJLcIBxoZZ/
HU1J+W9TyLPOH/0VCKK4sHrSIP6YVcaMZLEmAelrds+Um2fOEB+Cap4/xwuYEx6fn42Rs3/mRth9
C7GO/8vfh4MAmC/vD6A0Fxy3CoNPugWgLidr4F7GkvMp5uCVIwrflMI7jjomJuzb9c7g8fyFO2Pr
HLB5m7nbHU+YAMgvjG+JVAXFZgcT89/71p/XdL81Siq0fUGcIQHx4FD2lGUIkbEKp0CkDrde2CsQ
JxMjNUpGTGqMuQ23lLca+nZuDVSfRTA0mZKbxL+ubiT0NdyfKudvpPh2xHli1ypU6SPpwLLwqQoX
L6m8nZfUApGLU2EW+Wmjq5EpCWMpuZNPQFAi4Z6J7kJ6c7k1MIbzPCZKT1s3NcaedpHFMROQb6mD
oia4uNj09A5Pf9l7k9YR/1a72+KwSIy0NNw59+OR+RvcSZZSVx64grKBTbL8clhSmWZmyhEBksOg
Ah69f2SsW3HloLUNIxqpnO9acxHY1/Q9DXwGsI2huqfmqadigwHN5J1aFK/deDejxfSlYoQYL4RH
FChUnahYMFfZrKZj8ygrClDoC8g5o8aeD78fP3bidhqG4aAbKXEuP0kup8NSaYf24bcIDARW5WV5
0oqQHArBE5n5ijpinIvu9L/gBFp3LRA0a8WerlMtD3p9Rz1VM2VKILmaXLcezWP7RmuhCm93LnRW
NqMoFDhfmtWQt3l/oajm3SPGvgOzzvYuJ+N8GCVoaIc2/zctmXFdhQJR+UflHXP9aSkGTrTcHK3w
VszEGGr/gZfer3zqT9pfAcie62Wq7OCgXup4dRyEAwn9RExYaCr4Z04d40CWkT/Eq6zoPgVU7sbu
oa6K4wNl0Y+ye+tSXEQP3keRxN2RQnHv679pzadQJFo0nEytbBCAg8nYsPm6UXTI+88DaNKTXwgV
5So9c1YLHtFJo8oSJOvhTo7LyohZgsSv7baE1QhDz2v0XTA4P0cEoQ5cqTFKjwRqrxMukvfEI/6S
EJK8O8TY2LGvQVq2KZEPOZfGX62fakp112qz4Xq8193bgzVOK5pwvJzx15m3lbzweFXuElCoPoM3
mY7akCUr2CkfRaT5c4TVVWar/3Cd13TojlZekwVrujJlkWPtCM4GputSjYUiemrQqIZjtbKn6MpM
ZkITO3P7HkbI7Df52XQ9X88BjmLnGs7Uj7QCpYPhgdSgS2a0MT+jVZzML4AiJgx6S8IsLnCmH21G
5PdyMPkKC16iZEdCraXJpgSlvo6nZsK7pBeBKyBUL2M+/NWhLByuCZgAMPlMP1WzqhtLYpag6Oua
8AEaB2Buvmx2NFfgOk9V5g10fDLsnw+qDT75WBlXLHgEfBDJLiZ9sv+SPFExnLUySbMj9lW0Zj1I
0m63Wvcy1O/dX2rDaDffvUl3AK/Qd4h4Zgjp/7OTtEGh7MU369vk1kdpZXXHQDrMQqfpZAckyFGQ
Kenk5VSIIszZLTdxVA/V1Fp/2ghJj6gQ9g0/8+U5Tnbvz8Virh7AeXNJrQiYnVtLOtTdyGs4Ksn9
nJEU96366XvpH43w1XyFMbo3QNO3z0MQthdsEiZHIoP3b4grseklgEgrrQO6eRDog7AHVa5zHVwZ
uZsXnu/dTlflklGzyK/QojSAHBzWtjuhq8JVga8USxvTPirDXqfMD+EJ6vjbJVdAYubIBQ6yOM4F
Jiyvaod5vT7Bjt+azR4RoyIxttmyILAz+M5N9z6WN7Dbih/PNbt37nHqYNZyuwXzHJNOxAyvAqJy
35k4y8/TpizJUOdLKI+YSm2GAqDrWYzYK4ez4qGhJeH8pVZi7lyuKKi2paMyciED9LO+Ix2aEqUi
cNThEXO7snfBztkacK4e0GcL232IfxtUqJUHovMqT4f3YRMLtPSxj7k0Yt0lDDqZZoGxTHuZHHEH
G6VyoT0ApHWLI4jDXJZ9YAFgT5NM1Z6ibZM1jJM85FzqS4WTK3dLiKe8TPA1iPUDJEmo4enoEFBN
ElaD9Bsdz+gCXR6gUhraK02UWdmtvUpKJcRhnxQWlz0rvWMhy1PYOY1jLraQa33YExonsTydxUU2
8Sov4IeR6+NtIgzEDeIHj0RdLO7z70UtsqtBf4/OkA9tCAOqOA0TO3kHUsrdtRC+3n0rdf5b8g6Y
zPxu0U+p733qHlSPlXgpP17wH37PW9aWFhhAxVk3QIDMY85Ww5nosTaQIXj8QVDF0CzqzrbzQffa
TJaNq4At3Ir3AQecSOD0BlH9JuI4apH9AmvMXAavjiKt5aIRx/5FYz4T9NTBHseeX0LQzP4AnsK/
N7dlk2Ug34L/p1mmd1f4jnBZnm9YXe0xiGZVVWE8i6knANqR8sN4sbIzOX1BS8Rl/fOYw6hFWJ38
Yvl94cujM8tNC8RHEB7HZppp/hf1FQFjysNGhqOwlCelp8bKV9IzEVOzZA91ogC/8IByPq5LQqZR
EzI3ihQcmM9jA9sFtXgHzCmskAPA/ud/Q1aCEZbOWCLuxoR1otKMs+li3sj7hkey7pvdPuZHw0d5
yk4voNQQHW+70KsX2609/cjlgZGKhrIYnJGQ8B3B303l1BIER8R/vmBTgkAP1Zc9YEuVYcswzRqY
lsRoYXc0sxSBZTYoVJQtyslup67Rl/EJthhG/AnnMZEEF3Aj2mgjI3vCI3lbp9zIcstVzfSZtAsw
qQonDTioyqN09E1ddDjSCgm5Env6i8bIQzEkCLypsqBZNtUAcUMIh61Un/pHQdV9XBc+odes/FjA
Yt77yhvW7jAZ97VXFyhFyOKu6QL7IEHqm3YaSnyQI/8R0+rIjkzUfig9DDWygecS1WSKrXSE5W7E
MAhZjY6rUbeNJQ+DTy1oIlmiXHIN4fnHNLlbyoPz/ysD6+qTyfI3f4PbX/MTsBVeZ7z0gyizoi99
wu51wA6wKeNCto0JoXr3h6KFLz4qiNAZWjFD6YMGNXAnvMcQRnPyofioZ/XYiyC2xdh3Agwmx8wM
hFHljJ4x0VWw3QDa2BYZmhBpcsW43aBgBYa1Xe4gY0MeDJ4mJvHyb1th8fZHOi8roIzY63R1Qi+N
2hRCJYALZlVOK7YSGXoDfUX24GjOcB52Xrn+f7w7/HFP5UfJYYF+4BXktKZEzsVvo9KTFh4zLQIi
eRZlwoC8Sfm/Xk/7YJ6Dk56vjDxhaZbnr3EMcQ53V7Diqyhnic+OS1gZ/6QowyRuloWoazXSqe5i
G6lerAQI0W0UrzD/LLOT5Ped18PjOoxkCgTEMLeXYcaxL4o49Zl+NeqFUMIBXyN8YonVR9ocxFSE
NALQFsW5VGfu+r2MWHx43drqthaNknX9HaCz8oL4ShHLgYmRskZHBf+jzAG8UQ2K4Ci03Vb5C8+T
tD5pMw90Y0Oh/6JdTUx+OQFel71OSSyNuRh78vEhObzLySFJzr+/9cLyfDrxVV+YxR5d4mv5utpy
V2JMPBorfWDYK9N+l4D4RHFr4rlmLwdsti+34LhwgmK+lQEkGSvJZBe9kDPgA6mJrMwQw51Zl91q
eqm0J6S+D4ax91hK8XgRiudODN2BKkfwwFnwVV3P/WWPkKQrLDz5x2xijXlFc1Pj6i5chzz7447a
UOlvMwHbnZ9ilsAIo8D2mlZFKK32VX8LkwWQ8Wvk0jhcWcTtG8BAGNF0iLML0rs18GgjkyCgSDTq
dK/sNeRRPbLydMXcTw7DZINLYfoF0Xb5FdKF9oPZvL+OWwMLUiuV1RzcyI6cr+YuGb6CYJ8eeIEM
p779CJ+fgNouqrvlUlQhozPtKUms8d0s8R0jqqhb10iyQSLA9bTDD2NyRPmjrFTufGK5asP4KqQS
LWncKQnuzfHRmhgTnt0EqGqIFQuoiRKNcvhvoA+XR8ECO941VLa45/yWChHHVmUzVPnvuXYiqEhf
NdUvRUyG3BgyuyRXaaKfG15cjK2DeXDIObh0ntyn5Hccx9mRrTXGYOUZePQjOvQEq66jcWz8pX3P
KwzvUVvSwcQsxlU8h9b9LgSrmTKzFbSe7EFovVq6YKJop8Cn7RDYSAtl4fglSWk6TUFUOCOocyfk
2ikAP996tKAsawV9pcQ5YyyQ/YRF3x+yaNvZ49ytAVeUejvsHRHiSQR+bJsgTjXFW8ovNNJbNfca
i+19Ij171fd20bO47l2uDI0zFE+K75ZgJIFWcJBSuem1Yn9TyhRszdxysRArh/4ZxoQPCJwYDuKW
DmJ6Py7cR2B2BPw9QVmlcrIZBiYP+9SBeJIEJb6kPdD9aHOVCD9tlk0xz8FAqYdf0lNo59CkDJgs
2zmxNOWE7lh4Tb4cyR0FJX4qiAYEJ7x75/6Gc64SMiQ14e1EUUsNbH5utQMwYnE68/RLqooIwKWX
9TUL/TyZt6Mkbr/wd2R8/0nLbq57NEzWxm4qQRGvpAYP3GGK8nROgcMuyBI9VKx2/nQu6vYZDnvw
Ou3/ZZ04iqxwGeDsCHlpmWmJuEGsNOqoE5IiLPKwVsjh0MknjtLnci1LWKfZFUmAClRqBdsc9MeZ
cProc4LePBMAnO2n1+5SYwSGPNdvwPOtQNAsMNiN2ZIEHGsdAr8kHhOMT3fD2EWWPm6qcZC4ATCG
HwPQa4fGlHfc9lBwLsSNzdTuJ8AUzoHS+uM9bAiiBETqtpttnLD30O0uBW1DHOjlB+BNvuFe52kS
VuR3oN4q9QnT5T7ZilVSO5kmhoKlLZxln729pQGcBZVDVpFt/8e0ntDB5WI6V5sJRGyIaEVFJZHG
MWIaNzjYDYVvm4hVyVJIUXXK+yND4a4rtXmcaAlMz/dBdCQjz7oFRrODENvrWuVDxnVBZQN94jaQ
neO3kowi6MWx1iuONtbGqbuB7p+F70HWC3711qqRGeut1v++sJ2iN61oEPmBmaYzw2N3WUZairx0
lJbpejSd9/GiMfTG3lA/jXj615qlWHP7nPypStxZg5/d0epAsYRMNqZvkc5sqC9bxChx10U7+yYF
ahMSVpZsFgXeEOOIXDLKBaRBDzB1uNecfvHydU05MVIwCnW9Dve9F3UPDQ0Wo4yaz8IR56CwmXI7
4EMQxeC0ahB+osvfSc9BFSgtY4quskuUM2FegUAVnxxAfJxB7qAyeIsk5Y4ltvKsZjfHy2CE3GxJ
VmCgSCnDkZiORZy8BynTWS2BP3VZ4zT5yocl6xAjfbx46gWs5Pf9o466YY0ZmOom2UWiCCklpBzB
fnmorQD/oGEGVem/xGk9yMH9JU+YJ93wtrWRqkL58JUt0xVSktKqx4EeHr2FmM81EOi+M+Tl/2d+
jl5ge0IuPaai5hulF3RfSRH2QeiibB0vnQ8sIQEc5qEwf39L3ab9B+KSlYVfR9aeA4LvrWXS5fAf
yHf69aqhppRoZZpdzbzq9ple4XeJEAXHG2czl/ciSnAKM8KH5QaJ7mETItebHXWJjKn2uD5ceEfh
xD/i8i+IEwVZs/xJULnwv60NzFJgqNDGh50HjCcLUp2PQw4t68s2Am5NMwhe0mi/8BMSQCns9Ooq
6Fkfjs4Nh9a966hUW36T3Ame+LD3hFliPmsyqSgmAMxd367oc3TKfSlXujLYLx7qy29CkcITvvU9
F5cPPAmSDDCGDoUCvWtSmY9NDdf2vLF83FYhP0RbtHSdAGwsEy7fYb/1IUZK9O3dHVV64GOv4lEC
BLsFtJCb99kQ3WEKAWenZNk4jURTXzZ3ImgYriOtVP/zwHOyXh4TFaoO5LhEDxkaG6zLnhxFt9DQ
287rc0TCrpdITkeMSoOrmNWtrUHwmGRqaAaU+/OWGjNfU3ZD8CZpldXxHwlEGB6AMpSRfJKdihtn
ONs3KvcHieFFkDXVLPRdevxZ6e4YpcotBN4ox3YF0HxLh/9w6ivxJB0c9w1mKphfef7GN7f8icTp
nIfTrbc7yg8ifgKFS1qdj17Vi/ykIEm/RndO/AWVsScnFOcNDZvAuGLnY4u8BS7lEIo63yxY4Hww
k3kHVdHcx6EODD48+eK0tEYmaoD70fEVGInCCe82bMHG+NXg3HoWc1e0IQM2MvjF3GuBlzPX7dM8
sxg1KaEj1vCGuHrk0XibQBOABfNplQPwJy1wmgtEQe7E5Oprj1NLP0dCpwrYezAbCsKSMl/mxcLN
+PN5+4rEy068j1Xb699ppavo6X5IuXviLENZ9nyXXfjy78LG894cWsG7RMQRD5bCfPL6LMjzRuFp
PD/fjD/2QpcGhrRtnCdorMQUuIgV6jVP32TCg6r1OEi1IpIgQOsQH4DsGh+2FdtwbMUDrSOnUQpk
WrZw2WB8E1L+3Lixm889NBVgPiV55uC0nBS20PyE+eHmTa7WKxZZVNSI7VraWOtTh2OCj61PmtFO
xMZ9I28ZLTUbJrKmHWTIKnKBFarqoJNauugW/6vS6WmXYobRBpUQlWyzZHAs+CrH7HQAAMJ1wKK7
trqt/y1dj/qPGLdvh56iZ7eNZ34hrPaC8wr8AYbPHucrq0MQYIWJDM3z60/6YMuXlRyQnyaOZbTD
rKMxbdAWrp1BYO3r051VjyhryfDzSge7jPtTCLrkhpetsfuAJHndt6qv9O147ebB5esSgRteNYiZ
4Ur9HgvNGeb6dFmzQh+W6bJCoxfcfir9GytBrnbmMuJAyMmd0xxRxwTEDa//mgjWk6xhcMbf2svz
6Wtdwnx/mDR2cHZYxdMlvg0C+VcxQUoRhqElbCYdSJzuv7CO+HTh1n5B7RoVHj0UYHHZ68D6Tayr
UiLh6PagTK+BabMv3hdwkYHh3yV89jnRFIkp6dHhxtXpdhu9BzwpK/D6SKzcrnsOi0syVzf/0Iva
YtVPWoVpoOcDtFdtAAmb5dNMtI1X6D4OaOCoZIwMMfbRCdZj4HNZxwI9ONPDiSk9i61OpwmmQ9Oh
rh0yQJbYTxKKsBFLaYOd2MIDa9XpoWB9Wf3LfiQ/zI1YFhgXYpwpCyN/75w7z7kBOSpWOJm6Lsa8
nNLdPVZ3y+s323pYgkYdJsUH2S9xoQJbYKRDzM/DYynSbN1hYhHkqfwtRNHPQ7Bjdb4m25Xk6tPB
dNHWbuwwsyN25mEIjA2nleZZm7Vz7f9hNqZf7yQyRxhaSKNcdst0yC+AhELm4ROBpYKGD+FSOxWf
ym7n9dl305UjV2aYB1Qjpp9OZsP4GAIqGYeG1sTAeaQfWOFh6YE5ifdiRnVgG7qzVq8HbYhV5qm1
yLXQH92MALlDhh95fksBxvwH/ksG2ENaQQFdFJ1seb8WvxJNB9yoiRDC7NmPfc8U/u938IXlm7FT
vaTo4po5iVcAmb24I5BbuuaFk8LZ7rX8Tfw8M8mfl8foBr+XRQHnnDtkDyuCJwp/+UxlrxSVNSOZ
tzqbIM2MTYSLo58kJ8M/eiuii1fydhfFKZTjMCTGOKeTj9eJ2c7+0azU0ryU8QvFkF/vIVe4wHR/
npvFLJNHC94/7znrG2Xj4/vtIvg10gZbqh60wV5fWSdkNxaM1uW28IXIXjzQfa1Osz+qz9PQY37b
hQOXlNjG7XrZPqLkVnWlK4xFJvXv0zLmPrsIkA6XWcg96Y1xWdvuDjto3M5Ws0zQsfdKqa+FqGzl
7IcIPCCD/HT9wu0h02CKa0ClBTnoDha82lD2TBSaWncoK928H6/5uhh56pa2QkTEU0yciRxXEivO
Vmw0DprSLjprHH4gyBKRUDS9Mjf3wihK0fS7icUs4HYUaTktjVs+ZZHF3GfXZ0f6tX8mKdbAERyv
d0fw0w0BT7h2jRvKNhLYysvI17puG5HGdZORZT7wgJS2vpA+OiCSyhIOrqIRu5hWCtzh98MOF8/p
3o53MV+We1Q5KcPC/rbSrkKBSmjBM0ROQEhSI6C1D7qQOziGe5PrfgkhBz614dT5KUO5zM4/LB4Y
2oKQBaiYjRXk2hCdSmsfvQiM+4sVtREpHD7Z3aFz66L+2HuKdEtiIzoYk5Z6+KBScWzrc2J6/bVR
KZwRDKy8mlnWUW1H+UpK7CHrzRvEtSgVpchhJFVRlprhpXp391FJlXXvoHiD1BjjDLxHThDSsZbK
8MTu9I0O4+mjLnVHbqRG0LfmUP9CpdxAuiT20RaSsqtmkKrxI2PTSMYCYYlc+9675YF/1rT3R3zt
ovuRR0VH1x46XZYI1FC1wkDnuXdZnjITdphHh7+GEGBbbVQnnxz+wrZFslsnCb2jKaFC0+iIqMhv
psWfQrVq13ZfrEH6yBYMpqWvcmyu8ztMMSKtzsiwN+hqizTujoJLUkCUEY8j6vjxxXm7YUgDLxUg
+HPx6O8QrtujDh2t2MtOE13q4swj+YfkJsEvB/9XvX1s/d1Q0DjQOuiqUFPH3pEgKofS8nX+bzRp
euIzTuaJ/goPf7cqKtd+jmrJFGwj7MjzEE7iIckVu4hKOnS1TGl/4+yrTACPgANuHn4DEbvSVYD5
w8nRPnyxVjXkvsJxN292SCOfujWhJxa/tEc9fLXQqOek7jKqu8GgRe4zO1YC2tOtl2mGZty4AW6E
YlELAf2NvPm/k+Le7XKBpvB2ytySk9AGSm0E/hKggFxtgZfLwl+4mNFHmGgM03rC5jZ2a4cU5VcA
FHfNnXnVv+mL2AJbHCwF8vMUZPBBlVfXfNcgXp8JKYyYhgN29vEIBWITbpQtOv9B/GWPjafxQmGn
3VsC2A7DTx/cw9sZJdHVeON45WCyOj9X1N3O2TZYJdWA+xyZNJ9wzbRFJKjOjYC7Sc/WMQ1dMcHx
n2BxBN2R9hgF8rHDmUdi15W+kGB79s1iTewhcaT+roQyHKIGGmoLn1TkGETfGGLixoyW+A53usBB
CzvBBGeTh2VmD9cfLSXnJxUemKvZZ/L0hk/x0J1TnZT+FEGpjbx27AYNWBNyLy0EWfpC8tcnefKr
14FrMTsSCREasOtjx9Y8/s7SBAqmFOUOTuK5FyV5uiLD8v9f8cnQEiFsHaT6JQkcBKC0AkMfbv9c
TMma93GDxxX85YLulvYurj3aDAqII2j08PUpwnGHrkZsxKdYwmgH26TLzVSE4iKADEeXsgeX2uvW
GqrDZTTkHnceSF65NKhP//ebIZgCgMNafQQZJZnVZZJdb1jphBYJHaXLoe9Sc1GVRuR4hR2OlhCD
uswNlsyjRnNauILyshgDgk0rQj3BlPFremfhniYL8adaRGWMWjS5DbYJIdwZpW/5PCrSlc4foAOy
MKbJT85aZapf/fWEODSC/a1cyIHEf6v8JQU+fonGZLg9DgLIEuHLefQQyfRFlRYfKE4Qol7mwELh
4VKBDXntVPL58lg85wadBOmQ47n7ScYbKlBHxF2mMsBIH97zV4oFo0i09AuYh9xHB3Vk42ZUtj20
53gyipDZr7lKjJ5X2BNFhDseaxfDMy4lG0dhSahDMnWUet7E0+UjZwDDNWkhxqAOQWwBax5QO7Hq
4DJEbRty665u90pKxAH9FkMw4RS3+t4I9It6/w0Ql0KS9qk9DFBaiHgmTCPD4oD8wYzNeO0/FvGM
CAA/sp0z9GmPUrj510EZ4aAVvqr/VblA1nZVET48sKTWL2l2KOCl7ch0VKzhRkqF3kqQUzPKEmZf
RIYx7igzwobzhnZsh5nJDp6My0sb4sugpzg3pSns7CW3zqsiKI+QF+OzpMVcYP6E0zArNjYXFoJW
Mhw3aS9aefhoTxXaOQ5rQfcD+NdFIgCfLyesblrTio69bkewQ9Lk9gzNvKxrb6QeaknRd7i7Z9js
OigueFTGnyv+VBLCaqha+L6TnT8pgCq6Zj3wy4LlxbHm2JVOii7puMvCFbd4i6KlObzh98n36OMX
PmKqgF0gGeBiJHgZY+UEJbL/ZPmF7+XcoM4dhqHPK7pm2zGdgqDu/wzFnK13dAUD9CKujOmZylS9
Q1O9/u4+RlZ7vTJ8zaq69TZG/pRVCme0qMs5CGopPA53tb7rwcoDFDDALg/098pk2qAP21tVKAXf
tBuCmhWTQFiVC8rcmCwMSVbsAfO1hgB0dr/YVkgsdSmz4lEvOUuH2/uYTwXoJHnzCTRy7/xzI3Hf
h/KZ5S1jvYszq/FLP0YAjDEhjdvFRDfbIPvxq1npFIs/0yPhQ6+1Gn0G+JwI4RDWpJiWT8Sfg4CC
SXl2VK/9o+bDIMu1AHFa5Nxab/PHAfrb+cNbTXHKPq0GFN2rXCokd3+/QCHvNpx9QVwzDRXIATUi
rou3SM9Mxdf/vCMz28RNanaCyGq4ZEKVV+El2BXaRfCT5McSKY4yFMKH8vgYuGNn6ypvRwHBJVZh
lzwhOM41h4CN0Pel7SEB50PBldyC+qtLzz4lDFZoMZhePY1gLFTn9lm7fKjFSKfseKCPwYvEhDY7
Z9tlV36JhnrLCW+I9+x6WUzPsPzR/aW57BqQ5Iw5eqgz72KvfGtwe9TbWf5vsX3jnMZ+9If3Big2
GlJv+0qh0YrJdBfIy1YCPJIqzwHITyHKVe8MFgdKKSVkVpVACVt+5VZpNVJ5WW+i6E1BEAR6MWEw
9yAobeXf6Y08khA0AIPkEitQGZ0DQhJg68amP8nXPj25aXW7anuG98aCV2lZvf+IkoIxvZZ6vVEJ
NEPNNwBQ5lqO7+jM/DoH1znl8/zRdApwGHfoe3uXxkte6rnZGcYUkBboD8GSQTOYs/4h+zOho9H6
ZP2WHnVaBGwQh7vY0k1IN6pF1xMZPkeIoWLfqt58yi3XokVkzOiTkz95n3n+39YNDm2mNcCzc+2A
kV/gEWyAiP225/7VDKUZnABgg65LW0tXcT6bWxO7D10gD887/v1YjRropTWevjLvviURFlGJuZPv
rqX0laPytOh3TJhEB9JeikUNcXyf/NPwj72W4LD6TWg5iD1q2ru63LQVHr67QGpbwCidnvE0wSIo
cCJFeWKGi1fovTxGfECrpniJGQK+SJocK2riFza4Ra0a+Hfb1zQ6kTWAk0lVtMna9zmlTO9oYLXc
cxYXeLPIMUzwcPcKVOvZS2COTpoR8LvFLqG+Oq+0Mku50dPP0B4WX5CxjSdlug2EJLrg6sNysz/7
XCQ5Z88xBLn6k5ybHt4UmY50Jd8NH8kOug4/lc187H5qYwoiiHirwUJ3wbGOYIixvqm7qb84ld5k
pcs0sVBCw4JdgxkNg4QMfH589qmtHu8Pk4SyuxBNW7fxBF+YQ7D/EoMfZF+/iPzDmy+fIiVvX5SF
KBhS4XMHS1IPA2vsNT35JI72KWJcuqyi5W78WyXgYYnuzP1OrlPh9FMADN7bLDqzjHB+/O5EKr3a
uC/0YT0tv5i+zzAYOeflL4MMko2BNKKyOpuwrcWUIVdi1WGyu8dIt/B/ggEY2jG4YWuDpm9lfLhS
zIPuNBALuww6Bihjnnztqouj+9aBkbuD8f5PoQQI4jVWWM73/IDzFtaBuu6nxN029RHFN+MQY+nl
4zarcE5nh4RwFrO+J00SlmWxiwYihMMB0YSdRHdSiQirF4ST4Vp0c2adgq7tz/mh8oZdAgk/X0yx
ypWIeQuL/QD3ZNiBb1mV7iUowvsAO57Ej7AHq1PN1xB63knRAqPqOkEwoZWWMrlKTNzsEGFOngwe
132jSkFAOjAZQKIDdq5DhJNzsidglfDYBVoyA43Fui6XHezSHIFvJcmBdEbHJcmmOTz8gHtLe2GC
dBLKkAMaVBmrgKo2SOMOYrCpP3YrGoxhMJyUb+opyqCryyCDreEV+b3f21Vruv1I2CVbCmTxupVQ
YCIq+HbnntD3efc9HA8EKPDIBj42T5ePjIug9uvW2XfLwjBQQaLnQOWLQat5bqcjRKvoovT63Cmx
7YmFiPU8BlknshJhmzN8D+PhAtlkFUqSFBfu3p5aajDEdMpYlg7Y8xcI0JkUooYN3HZJDcmFqn4x
5RCfY1b7l9EE8KkxibKFlTg/IDUCfs3QU9xgxSjpq2va3qWxpuBuj1yLxOKjXhQqWvV732g0/WU2
vlHqeF2snc7mngt0DmJwQiVg1WEio8VFYpvDOLXDcZp/A9vE4h2e2qx32aI/9Rid4YfFNBPDI247
FJL+2cCJi8hj/DEOklA7cY7aNjF6pRwFqzAE2TqlPEL0HqEix/IH7hCmXgkkFUBF9YXuQ6nTwu7q
nR6pFryPI6oojS5hH+vEwzOOv70OCL0YCuhCeEF8iy0SlfsEQ/cAv6DqV27nMERXdSbCM31XM5AZ
gRESzm7CzAg+Uznkz5DISbEFg0DaLLlUFv4oa8WMaGw7hYOUEQNmVaSJloE/M8przejy7M5iMlBS
6dLIsn2DyBNadO0Fu82iPAw6DYHC4yDrolSEgUH4AOPL78GEhJL1+0vOjSt+OQiBG3eSigJm/jjZ
SBmvVNKa4CHOmxe1Zez46eq/7Fx/QQtdUFYKNHO/j3W9thDV/qXVM8gPJvx/VXis4iG9AuQqRZva
EO8TcQYFvnTzG1wIlroZefuhxTFnGhtg+PmTH2TxXJ58iyC4T3dqSBKRJQBwnpZupNmheAOof/hN
lc+fslJAp5hdoIbRgJvekEg9eGBrExnv2hq/KsDPrEnAl4Wx8P4xOm+KZdRqp6VkwW8UD8HSx2w0
UZKPFFh+7VKJB+RUguc1fsa0fD0iTCvTa3EGXH7aj45gmgCLiXtmbaCD5YmpFCeMlnnWDtFpOho9
JATZ4CofIlJdHYNrz+1whan7aUnQc3yFAUWKp9i37nvMZS/iarlRHaGZtcx/xFxoxR//zKkxFTaW
WwXAkHPIKFThsjBODJLkZigg3A4g5WPGSS0J4CNphDZj4gwqmsVlNAFByTmwbH2i9G2A3eOT0jFj
fO9WXZ9gqgORWu5vqjyvEOnaRG6QYvLPkhFBPAZDoafeGfPHWguLzL72jkscB8EUcMPdrJcjk790
cxPwhCYbN/1GhAc03ji9G+tPGhPz7neuWLoNMcCTCmbLl4WfZ1+QCAwwR1qMjpYug5aEVBWlDYtX
qtEmvE0c3Td1byz6YzBxuXdrsfSUf+hsWt0305cu4KptQa/aB+kHnwNFWPDye0tkUSEsNokaGln4
FhT03odsi2mZH6gU/04XcyIFXIVcrWdqvHqASv4FCBOrJ51NuiqPwxY1cEwCTnyItm+if+m8EzYr
D0+HUhQNBXxmcG0YVk3tJaaQ4o1roxU5UfyhZ4eYXpwwdrb+ai/76Lb1rOaoHSpBjKVXdOUM2T5W
B2wvar963B646eHajavX6xUZCmU7C5EZq9lxK/i1gcrRnJuRMJVb4aQ7Y3A2cTJyBZmPMatLV9wT
5oDo2iV+zt8A/wAui8HHkCwJDynI2hQu0K5RchokUPZ8ACPuUWXbubHbUBhEcS0x+KG3kmYmdCe/
ANZZDY3jylUjapytSBskZx+HzRJh0Wi+zVZ3U4feL084kywQR7mInnRcN57TjSMS/Z7+pIaa+zJL
zulQAWbaFL0KBWgb2WkiPBGjhF9WLyJZDX6Br9Mt7jUQzXAr+uF4PGj+T9aho9tPYsai47k8Tr5B
H7H1JLzg1P2awARfG7gUOBgcJhX8qy//xmm3IDqImXLpId9z02hGV2Svvre4oCiov3frJG9uSBsi
pTemmt0i0fGOQZVEqkWBCm6h8a5TYwkKyZWBBUm9vMPOuHmv7qCA8uzVORmBoCA7qniEh0ZRnkEo
B5sS56cEel0N/L4aChJa38JUDGWM6Cdva1Vioqcx93Eo1RfRayQqTJFC+ZGohJAiqzCgLFAdHC8l
rENr5A6EmNWb0JChgB/zTPzTAqpSrW4Q7L2Lh3VRdpk6yu/AVIih+tACFAkW1SMINXOftn4Hs1S2
qwm7T8k1oMelQ/Xf3qPQm3Bubyx5JuQhhgLnIII3K8vc66NADFDMmVPoOpoyLzzLmOb5NZdxxR9y
VTGlvFxS29u6fgCjiqVtQKsWxwgd18k/liad5SCk2oT++vwLw2SaY1dfOQYSNZgN0sS8CZVmj2qr
PHow0Ga0e2LTNTitnqvwoROWAN93vyY4CJG6icKWh1b3YFmtNm4b2GzPqEuUIbdnjKJJLeBGOklv
WSuRPuV5dsX3W4sdioTFqirt4ox/AkQdD0w4uZivacXbp/54MYfr90EGV68KXkEiZrqsiZow3D7K
uBYaFtAdb3VyVrDj1Y1UEgjQiLaGC3Pudx5QAe3uLwh6avFUSyuZ3Ek4uJWG3NpvPuT0KjAY57c4
xpLhjMH1Sdcr+mVnEzyaLclBaIH1vLZh1Fp97WlJeh/bUuN2aDVT8yo6nyHspwIJ26WEUmdNenU1
zrYFKFpZVD9iKsKi4eIGI3EF3+Tb4sKO3CNdGRp5LNWX95Z+5xbaDNAQfNdrkYUQWEjHmBmR/VwF
ou6/IWsT++OwvOQ66M/NAFeCFOG7Rwa0WtKWgO/QYyVlKSho1rl8Vv0u+rN/W6zO+tERBF7BXnaz
7ckd/vOc2lf8PFJnmb7+5HxVrwZFlUCNlF7Roo+zq8skPtbn093I8Q/TUINoL3mHryx4bKB7du38
3G6hGJmfIRHatkSWuzmahjRkTc9dVbp/uFhg0J5DztpOLj0OSMRoDmJQ7Znc0YND4i/eCk6TMgKn
Nw0SRgQRvtLg0NMRd1jALjYZQQIy89SDV7Z1zN+m8cyYFmdRzep6EVzpb9PALs7j7rRnabaobAvx
C8vsQbfeu9rAMYZIFdPSEukgwlaTtLdjNWotb1Hbgl4sCwSCxfulbcBx/8pOgBUBCzXJKX7J/D6e
i9/DRUIVFWZtlpIqL1ffvQuRVdId5zNVRZLp82ItDTetQgyTl27klvRnvHGJpZIidxoUxlmIb0h0
G0JWH6EJzIKBuuf/k4nZjdf0JlrzS04YBq/cnjdlVDi+iuW5kjv60IDhO/BdA0cZHthRGprmvG4M
1e/sr58g6KRwF1ynXcYIX//8IDsvbg6tjK5Fw92nH+tk0rQq8l3dKE0lE2ID4hMKKOXQBgDBmEL3
KAhe8pDQpFoGY8FUheF/cUo8utc8HlKm3L06TKGCbH68bde38dyP78VBkmlHzowheXIYOwVUO8pd
6lNa78Cw541ykD90ND0dVX2XxL7aKwQxMCfk8zCTI8/bsk6lx3kpNFJ7XtA0tsc1vG9kEMH19mgR
JLS6n1lW3rLaV4Ox9Bbd7qQgClkUalnBUhQgGTTjm5wMNrvYyACcOtQwQQdmwFqbZZNuMF6pq7+R
NOfnogQAmwZcJ+G2TnzwEXlCq4yIGW8bgnAqRT25dwI3WNzQaIt3uMj32dK/PaEH5FN1ZfSNPv8S
J+zCcXdw9MKf47mLMtZ0U3/lccVajnaFYOXQ9tTgLdjnMJj48nOlj5G/EhpMl1LKX4aqvaNQ45uN
KF5PHoPcAa255z2BH+WZ96rMNj4MqAUn1JkVDIqw/wfpkVLiAJlALGNAJds6C4C1Qz/QNpNhSigX
wXA/wPu7fB2KuxIXHcCo39LcPYobDDpATJPw/917Oq5XtWofZovnj2f7NCduj2EUdmap2cJZpnuu
Ab7hGDyBFjobtik393ClPLanc9YosVjjA1x06G1E9438NghofawrOUWqk1ZHPX3WzYCv/Z5ofZpC
U67QAFuBH6drUKYuzE8JKpkzJp3iKQWN246aDqQ8wFPhdn7zV/AkYOREq4OSGlhnghXUX930QU/c
AW1qXoEC4cDgQD3RatgjeRkhBTrX/GR5vQWVgPwXLn0bPL86C/EWHNOFUw4UU4kHBX3dESuGHQRq
xlWAQaw51Nq6Pi3B0saAVyzWEw6g3SwlW1EjMJZvwxOMjLGbzLuoDXQaeeJox6tYKgpzfimHGekW
qxgr+BKg0A+5y6LkE6HanQqauXtLxehzszHPtg7H3cFb+jiNpzOZuvbFgt7vClhTt8T4z6gqeEGM
Y75tWk+KprI9gse3rHz39E2zvp6/OPbg0Pb+acEsVrl6YBXTNMAH4x3Xm3ZaEl44VMSiKx5UUCDB
eq1UKm/4KUm4pdShz42doWqUmdTgjObuijomyxIeThA3X8bNuOk5uWEdzCcM9HufDyDv7Md4/YoH
OaZXYCVPxHzAK/Xw5BsaLqtostSEG+QVSZhvQGInHLSTzd2z68TUS8Ib9NJlLHAd6zZ3H6VHrTn2
f+e8nmNGsoCB+s/hDvWUCrkoZgDS48R9OTZTqlTTVvA1H6vrixXZyTaPLUjgBg3mGZjIFoLS7pNb
WyKhHpiZX3ZGCZcnVhf+lmTrmwVcgCVHkRR82UWg1tEornsPILFkF7ZPC1lgfF8kZgE3u9arIcji
QiPCIuBhY2Ul6GxmXJAAG6kc6Qz7aDO4EmlhMXn/po62w55J+hfFj2jWKeRjaodviABBOZ6Zmhgu
KhZ2MAqiCzmJRr7v/TTTwClAHfhchh/HT3CRWuL8luS5LS6NozcG7yhVU0nDg7SHmAt/0a6/FyQY
KmBPlaGo0vFTMuK8uGWUbOoyowWsGPDAzQCLuouZ8GSbI2ZmlCA2zbenJVXwQVQPyAFWukIGv+bh
jfPLIase3YhOJWXA9yt7H9nmIDMt4Kgolzk0XxXEmCH/oy8182UnogBnyt568bN5F+j2VmuaMU+w
Q0n93QPJQOfpYbWIYwF5NPOXZGGpqm14N3mwRTfmMxlVVRxlE2vd461S4jf7O+XvkiiipnMjwW8P
hrhPOL/wK+5EuxpkLPKnqpbGAz0HRkuCYqWRPLRPi68NMRFfLQd9KVRktgeGuoZ8IMSc+9D1iAG8
eev0ng58m5Q43yypisvB2HXkW4Zc51pyNgMv5JDSSFGoGwTxkJ32y+66ZJyaVxyXx/Kj2s5aUnkd
qiCdroUBwXGANr4KAB2WoooGAc+FC2VGmtwHNMxgEP0hI6QsKAVHXHvuqWH8d0leGa0yTQY1gdWK
wmn1774lFmG8Se7e3IUaDxZgzNDra34CpmDrixPIRssVAQxvjBOSRP5TmWkCcBoexgtKpnmOMrtP
sD6hdVGJR6BELjNZ4OL5NZiRMhUt7SwufnEymRvYr4IbT1P/Yc6NGdU/2TdBE6sg7wmKpsfIQJV1
RjnkmRPOsyUcHfzGtxPBciDRvhIRosp3U5cNw6gAiuvjgOPEGuV2kUK83aXbPSz4w7pQrTkeJqbd
qpNDT59N3Alg2OkPyekfYiDLNEXIlNIPW8TDLmGgm5BapWuBhiUzuyfZus3t1HINUcdJnMAWf/97
mbmZAO/C/y26N3e9u7pbVly+RmurKrGMd12cWKmusOhKnuL7dKxDgETNOucJfdWKdSKU0B0UkwzQ
shGaUCbChle0u9Ebz4hzTkacIIVdFZ43c7rKLZYCD+AzSWDDNZW/6kX73b/g5XdyPjF1s2y/DZBB
GsC1Cxx80G8TxC3bBTfeStb8Zy1pWLdK1pzxcDLz1bzV0ju1ErOdL+i5kC9ymOwBvAilj0/VxaqP
GhY81Mueoj9xMW2SXA1ECM5v+LU3dKTeccrP3DUjCaAPkPfiYKoSyJ4WeE+KOM1bSNql06w+Wd+e
V3gbd7MjPemiOamhX/YWm7uRDq8x0HWJ5UsS3BPMSSGsnWdRoEPeWz2phoi/3d1lHRGM3gBdk90b
igLgDiaRJGxncLon+421QQKImcIBa/4c6oyP1fmLZS9He58ktmi7cb1hcV6rzCKsLd4nFksP+TKQ
iN+gxZxiygxPLbfpmrM2viSSrBYDPrnXb45lL0nBRA1dOZiBcSMXJ7Mx7OyakJ+uh84nMmvOXxNC
jAoPVo6gsF0SuZGGj2kpyb4Qy5Y9MYvUlBZLVoXqBdWdNKLz2gnNSqTgG6lKC1gZMBVNnCqool+w
7OHz4q9KObWhDDpPDb+KGeeppBztuju6ZFqWYxddV+8ZdMszyj3EM9kFAESQSD1PpPVmV2AmWERS
gbTBs+QTyqoY1HiNWA6i0ZIJJtHrguRm/+AQ76TQeg9xWohtLNenYKSHyNm9cq0de3o0Eu8yDGEy
+cp78VH1ttFjhclAjLhmHOJFj/5kv0Vo10u6jl6pVJGNyEpTuE4/xoFSPgLmT6aS2WlYVpsVSI6k
oJlfEIhDDyXWylLitOeCVkgWM0duCzXW2TF67K37WIVsIx9apKiFCDIw26BJhPbPusaFr0vZnWZs
/txZVcD6vNBJuyPSuHNpaCeBvukOY5Z1Z1Sf5UY7alOmOJ+fUWcZRttLp1JJthN+lxca7WtYZv8a
yOD2Me2gazIfjQWUXZ4HnzcGOlNd/8oBmDex7hZ9q0sq64v/iQRlmwkUlts/KGkadtKPYBLa6NrZ
2eAz1Tvt0LZ12TIycEO6YZ7ymdyccgvNIK085pN10otzNgSOX/M7EM/1OuuOicZ1J4CpRis7OjU7
jV9v/ZK/1QemoyQCdU+B7w8BNdyY/mh7twISB+zjerewnQOdgJuFT2b5BV+jstMvvZUrbxl8bHTZ
BVYEVw0ERBUPo/4oNp1FJ+gQz/aIxTgM2Lbj9MWmkUgeN+oJRNqDk8torwboaVWPNIPij2Ua0+Dg
2Z22tIWeKntJc77Yq770qNZLZQa7mo8Ahd5SATpWpyR/JNYDjp9z13S8vWu8TjrASqsye4dF4ZQD
I+elJw+0mLwHg9BZiRQ+QI+lN6uN4FJpfZJC3SxBiYr1wEeeikEv9QWY2FLrRMoru2OmDyZoZe2W
Ua4lSFhievE8U00f4zD3JdZUJrDsMB6T7EtrKmm92kE0NaSLiXPAd8xSK1rmbtLsl9w6JVZQGFuK
BRZFyM9vxff6EJ9nNuXv3j0IcWOS1f/izZkb96NPImwkBe9LUURaLMtlmGUf3MFoDi5Zv5ihJFnm
Ztdtyim//OSn1o4zegcdPucVby2GXRrYfiJyHaSqXVe9Bc2XyeF09GOKGYbivcdBLNfjlMutZc8Z
EAEKS3Ln3/7ScqgNPhv114z/N3O175JaXVnM5Cpnyyo5XxS03E6bgg4YEvdXq7McOz8qHeIRKO37
GVNn6VP0YQzGexTGhZkgM7j8pDkjLy/00RE2K5wMNHbwHzwY3Jd3vjfb06CFoh8a+BA58T+gMo2x
cULUe7tQ+Z/29c1ivbQmeIBhlc9AaUzsv1qg2befyVSIR91QDHmOm9wC0A0S4cPPoyK8h5j3Gxj2
bSlqd2UBTxpKgvlaafDThSRk6zvf5iVsYZgRYiAk4yKP4ajSb15UdAo8eqrfg3Z/MS1FgvYK3DdV
gs6s1FgXWqTomcE2OX2uK+O4aawuHt5SZaM7ckr8SCqicSVXU0RlZPNaAuLmNZ5k6wLo65tvMmsY
pc0KO67AdeLge7K3Paz++FbA9EhLSJj48NTfy7sxyoaGvqEFMYG0yM5mWMp6152Y+OmX9+0IY+0K
pIO/Wse7D6hgIYbN//Jx1rPfhs25VYvgXXPxI88Bk4SEZXsWotB0pDUFRG+BHxRIcJQ8SVAL4yH9
7ZU8RZAQFsA0onc5xwrnOB/xWopSIMhEhqoBIg9iq4K3BVQqeqKHQiaauhckqnFH1+jXlZr4oVYt
UX1ULAQACdzIYL9T1kHA7Oa5W9b6FX5/ELWZICiVq2SSj+Ue1Gmgo0XhwXaw0vVaYf1KvJdPaztc
oyGyrthE2Xto4ZaknFkoo/YO8Ol4EO1n7Nh7rOhwFS4M3Uo98FSbImF734PtyiPBhN0849VNA51q
dvSW29yNg2yoogNPa81DeCSX8PBsEP4T0rBhtICTKV7nhjqO26nx5P/j8elywolqCTvRQgy9fH5y
Mekp3FkK1V9eHErm21ZTbnPdXoeCAWU7UR5j6Y1zoPFwNXbfh8UtrOckzrGZ5SRttUOtqGOm+eFZ
8VLLrWVkB8ah7urFnyTGmajazXi6aVpdg7Wr88Mo1CMG2je7+S//LjrzVbidlSbCKxq5KdC5jLiB
a4qGCvHd0OL7aPcqSTWprFIUOCTjQLBJDH3mzQf20Z9jlT7VhSYAW3OYSHBerntUMk4OkFo6b8Hh
7yeIgr7hgkJLF59DvL3sFHyDaJQcZyYWObhN6x5SMsifm+Q6ZAgVtQuh5NT6+D3mhxRWO683XDA0
45DyMALxUKcsHJtt0ZgvkyOrKIiokHWNnbb13/0dexlKxsRLMnNgZH75Nu6VAdX0kG2D+FGljCJZ
LY6/TgXZL2v9wE9+NHjp7C8BLZgx6yjAU5rRvv3LfR/h8LIqIm88LsALIsQAp6wIjJ5s7xGXRJpx
i6r57VPJw2didA4tUMlWvr214IQ68aVo24MlzNg0qoIy+VeM5mBCfPBUAY4HVaH9/EhKkJmzscLe
5E2+C77WPnLJjoddgScekBw7HJPo7M++LhcKT9bkkriUN5Xt9FDUQWl/P/cvljW1bNjPoF64f7o3
QjL17Va6n1w13mU2yFlqdW7b0LoPXMMgnncEr9gwKdvP4436cqR4/6YguKo0502Vq+OwF2CEAuXA
FpBO2TsVMiwlGNoQXdqpYYn81sPeOJvIk3MNpgaTcouH3LE8NapGwhxnRTLBMZPzwKL1A8qCGvk2
FwQj/QFP7Ri4boxBTpW5CkkMI+XL9V8sGPOTZlx0OESCoo0GvVNTlyvBIrsn+b3zLP+Qij7qXiqf
z+8JFqTAhec6XLFATr2HRSrSsy42d+xcI8zTI7J8qEdq/QBOq1de0qtZCuEho8xeC+gDB3H03kpx
BZzraVUR5nxOaNQPGWT4tK4fqMdpe3wcvOBqxOKJigDeZuBL+rYxhgiwwwA8DNpphvWji2a4KTNL
4uFOztswJDZhQWLpY3OeHaahEwxus4m0ICZumdxSKQgHEVi5cKd0nnMOpRpXOqtTMfI12Wgw77IN
2P9Y/9rgj0pR7Y43czKsZw8+B07tL7oPU1O2zJBBS7531O9XuuiQlY0DOanw6dmpWSn7grnw/p3b
YnJ1XZQ9IUqNDTmdy+XsEDjodNXgp0q/SKkykeMSPLZdKkrNtwZaUqeZ8N7p1o9Qouq1ot8RgcUO
ygMKtbFSmPFtpoOUGHnLQ9j6wYLFzp4pyZCtbue5oEQk4Mu0Jj/uaPvl+tHl+xZvjiH5MAcE3zaN
/dZxghCdPztbl0OnHSJcz3FS+5M+IN5erXZnvKUZQWdzsMRgLiBzP1Eko79vhueW5O6DNC/42rzc
jXX89ecFNDjo+hjBDLFkY/Z7yrtyclFPyLlKKsmyv8wEZoCfDOalrDSCOLBtH53ZA8C8pTytpc3f
ow1OzToJifhKYEgYdg04fN6R3VYWnHpW3l//erVrflO8StIhqjlGhpbEkNbp7SwVnvf+tS1S6Ygn
/tmQ7ZJE9VW6Rg7wHAQEqfELIOLKJg4dbmOvQTsyERJ7RnajBBF2b3UgwdocYqdPZ5zquFDRHD0L
CX1MrjVWx8g7TCaYAZax38n0DbZAx9QvPgq5HZhlvwJRnJ922MbVTZ4hBzuiZmvhppbGTpOKE84C
on3fpIXcK5+ZumwVQmavNiF3GdXDXUBxMqoY+/hIU2/FDRp16tmE5EZ8boZqNkbmA0d55GHBW0JF
xQBvgPy3fY6q07LvHrNG1HbxJlYoHrHxejY/3YEnCH3m7PdM3BWVBPZzXxKiniplj5Ruo4g3NYLo
/ew5ipxvrVSeDR5Wh/STUXSnTlKHasy5zrFKuQ5DAcd+fcOQC4+kbZaAt69H9kvO2u9iUwvbgCXN
ECM7Z449weUFUvOPohqlkeoN0Nnz6NgZLpcPCEjBa0D9MCscF+6UE3JMSXoI8a7P4BvFP6ynJJXu
99UPb7A3XIvCtOWs3RHH9/JvDAmHcVn1nbtTh9NGROswvfVHcDI5Ev5MSnnoQITtpef00XclDMp4
K3yJti/APIJw1Ox5nSYnJnUPt1YcN3YfGsRbPw2GJjKcIvv2Lnk+FUSoJK7yH04GxQZWW03yEsCB
lyDtVDSWSFB9r8T7G7PuLOD63hq4iVskYdT/cHOfKnaqk35Ke3qtWBoXNEYcL3G3vJGPStPoN6I/
0bsgrsjGjIF3FSq6BhnPjFgyoCTT3ACRwxYtWbtQP79JkMIw+4NlUryaVf7/wu0EMJItOd27HD9p
vWVrSMCYSQ8w3+1bI/Tyn2kkmK+cIh44QNIRH2XwU1agcMIWelK1L+fMwf+gFgLBI/NfKx/nkbag
WC9Zs2NNZFeG6PRrTTPAxmZvNTRYzOklnbdj31oLWRW+atRhJOr2kp55isP7tRaZkZWViAwvTAa8
n5Wy95OU3vDgpnAFYabkToOh3UMkd8udVs96PDxgigTCn2xNAktNlq17PPRpIvv2HNQ/kHu3shzQ
hG8Zk74Fc1Sre78ETp4SST2hpRno8Ih8Y6XAbogJfG/BWz2TmOsuuP0hdrz9199cKeFpprbEx+oZ
dF5EvtlSn2YRNoTs/VuOcc+byWgi5lXCkVpSXNBnfg/E5gMYM9/LVgJ2qfddIe2mx0UysxiDsTQU
Q/pp6mXKlRb20oyIiYZCfRWfjetzAuAVMk1JuBuEe0HHS7kmB3G7/Jk/SNCyQDcLsJ6RzllWR4iO
Z76S5359hzChk73RocMrvTWw8/iSLSoBn1B4znhLPw4vE/Im1LzvhkoPJ/VQekYQXcLYcmdmx2Gu
HMSJN4M9ZI/eCYE1bpPmdcVrATOXwDMN/D3W06FnDZXsXBZPNmyfljGQRL4DP1LCmLBTSkuH8bhV
PTOF8j1DqqVZSCvzOd7xnpyE4mbylfMZh1Q6SNAe2CJwBaKNEjaPmr4M7mY9mWEs33CNhAuQUuga
mUSk2BzNWdcorzgUl2q4o/fd4ZUgVrck9ybn9oLHBXvN/guCSXDmnYW+8z3VQ8bJogSRmVbPVwPO
i4w01EhoVzCbNZndsNGb/kuOi5G853NcWTrmPvp57JxbQKr/0WFINPDBAvkL2Gqb9xII/rQG7HmH
VkYN06MdeASeyKrI1BGBJSr3CUPFWE/ps7LpCo0h900Ytgd0FQFEOsJcU51h64GZ7ocKJWmUqA5h
wnEKkNnNy9Mm6HihCxgcP2S5w0JW4ZPotAFHOrW1NWme+Ks/FKo+UfmDzdFqrIFLH7p/+8x11utz
LdH9qjuez1Gp5lrrOIkJsGz+u6LJ1xi00kwenM6lfq5S26QVpK8BLMTDFxUJzsHVcvmuqNd0TO4D
X9aySg4EBa9QdRhkZVMAK64bYwFRsBmfUvGEEA2oAVL82/bcSHwVinK+CF7rTXOmbZmQoiiZFl79
77dxH5tcwoevYwRKqx3DOGgpm2mfzJyMSK90KWaQf/e8K/gXw0wrOoHOJehmOKUmh47YAid6woih
xsV96vSHdgNxzJ8xQnjOuqOk4kAcOJVcCWUzLwzcAWH8w7BeAmDXYONSWXah4wao7bH0x7caZh0B
jqmIp+OBF6Mqu55ISwuBfQyVJ20nM9ZOkyM/loiSutDJ+AV40+XK+oEx32bUyoiq47Rubehe45Dr
JLnNw6QX5OHA8/jxFFJJPw70Y2UzDHYx4JegAQEGdqlZc0CdfngTlf/ehZVgj49/WcekqoYTIHd9
sCymG2RCnHa4wCyWfZwZMBywYeWwjvOOYMwULopR8fJCKtPn9dlumm9EAdJcwIodnqYp9Gx9dcfL
oqxUS2+IVdv9/0PH9XJFbLv9oDc1vXeorV8ljvM5vYtJbP1WQdXPvVcRbUuS/Kh9AKHW6xNdhO2M
b8VzA/adOAORaqXkOH0G2tUbrQwHRWxvCcpVS6iUdMxmvL6J9hKQHF6LUFKM13UwRsjlqP+VKf2D
JidKjzpwD5kGjxr2/b3JNDTHwSiV04h+RyIf9ARVihM8J3IuLOpcrKh+ix2wO38yt33COF0tjTjw
LVcAlCB/NTmbXIWRWS6tU8u+0qUzdHT1rnwTXGbZH18GU2twFXewAaxj35y+hk0jimaO6AAdS2v7
Leo98fVlrBakrt1+qATceB5lUpZ7sS2x9x1tPZVovONySUDQgE1ESDkztyp1Xcw2nigwwBPZFhOi
1YkBxG4yanbrPQJDo65Yiic+834ORSKJsN5NCszytJmX8domKfYxwsVdSdxHNACYhfDdYIOka6dz
0n1UPVUo823BCFl0h5W0C+yeV7t0nB30fMVYQvrqwtFM4zYe5M2m+1HZGxC29sYQAmG8lToUKo8J
+LuJ7c0JFTTk+q0aqZKuvv1Td1QEM2tPAg17HNhYqXrFuG9jUoYaMCYLrPWwEc4eGrYlQuURauOS
VdqoDuCgW03ISlJFujyNsDqqo2qtPpgDLI9ykjNpiiMYDaem0ikRBI2C8yC2+MTvEG0jj0x1GJPt
tu/t+sSVzn+4Yo0FwS7wqE5I1V+PT9hGJcHlNc72i3Io89GNhSOee8R9fwGiwk+JrnWSbXs2GSi9
P487JN5QDThaEr/MWlBIXdrJJTdahKWKLBkMmsBABZhnEu77+cexbKXl8I6s5k3YN6WqN5WvTJJy
XVC5wJBAXsqJWPV9FcSSMCyns/uorlEVNDh/V8UkXxG8dAgVjIl3QEBTuF9v8K/NRXBaOjEc0O1q
MJPCLxzSkz/w0XCyUCE4F3VCc7I7RzRzDsuhvGvqUrqZdZ+lruqMx95H+YJYjAB2xKWVIiNZasYR
b7YydQYcVz6rIJUsUanuXGdyB2ohnat9gIzGBqW38uCZnAZccoVN+aGnAiYgsoW4mok5MmBwZpuo
C6/dExzGOLkWrf4doKU24wlRKXMklLQQ/guES0NwvxV1UUNw5gVDavJJiK0bgbZ40c/vz4YhMEol
leKt7AlTjm7GVvRHehlQMfkvQ/omqdtfgNKObtf8CF2MRxiyxZ+aiCkjn6KuU4pLsHnyuxgUGn2/
6OBx863/2M7qBQPPh+r7XL/2x99Ks/c/lZ96qkTwG/7IKlLF2QtV7jcNjP7lGx1USzAT6CtOWwz5
ST8EKzt3+rRLhH1Ee7Pv1NwmPAIdenWCp7MVPwFlPJHcKdQ89bmf19N8gs2pitm/fDPuI0rc561H
ZuW6OHa5pELZf145iC64eMYQSLX9Vi1kbLLgn9wNg+9JRDz/8+tWTwgf0mKEAY1WfCMxIJDrwy+h
PRn7Zn31hp5q2Qrof7L6hv++3+CfZGoSQ2+cvY6KMIKqDuhb807ByjwIZGYI33KsYQruy8KsDG8s
irRvpgtyA0pg4yk06m9H2abLKba2uGDXGYNxJlMo/1Th05ZfD6e1fzKLLoiTncJaM882gY9CcrNb
XrWRDjAhyt6mAL+y24lonVkhLsK0fNhupvkIY8bdWsucQuCC9T6XgU4Zed+iE2vuIIFNUAGhZNeB
f8b8Yf2i5E/sZ7l2B+INk6J7+0PmUQVWgH9Vm06WqkbdtYv2+m7K6ER/tfqSAKypGSeHTik3l/lZ
FCwEHla/z6jCxgHwYqbZrbSh2H+FfFnjbjX5HqBIyDlRN/Q48giAn7i1ymcwry8G0HsrVYS16PtO
03ZhAyddCV5Y/ZwnLyH/KK556KF+g8K/9eNNvxaX7ujwmeUP7xV+iFyAHzsQRrn749b/SuP7nrIZ
jg8rR9g9MtLh6F7NbFsy8yQ9/hoJ6RSQS51ynE+6gIOFzAiYEmvY4sRbqHK9KUhQXsS2TpjpqfvP
8p4MLmoi6pT4WTZxD8SQumdSC5fXhZ4zwqq8LMtR9VBaDEPCNbmXXOlG2bJ+J5HN7sUG25M3R8Lz
ilHv3tyw03JxlzyLM+lAYfqEz58H+NCJlV6JwLYDTk7afMSX8lPDB4cVtRkbSUEWv927g+iuofXN
MMIUUC49IyMreYV8AhgFubJEe3VivOGfcgQYBRprGr/OngevSWDKJ6Yzl/MIrxW3L2RM3y/emBp3
UImnzCk15wpXr3eIoPBEyUgFv7rfgEyZrUCUGR6M4NAkNNfCKAwIXbh+r9I5Hw+CJbwhFpbR/4w9
R5JllnHpdjszZW3H92sRovUB/nzZ7FXWm/HvMOeAeV6eWuLkPyXq/iOYjqSUpVnzNTowjbFru1k9
RnnsH5lA9+ujDOqfYFSBOmyzINnPklUHx1cpM3LO6yV/fSInvaytaeQMLnvM56uNPGEvwKeCmm/a
M4lC1uGV1JT8TKDX2/b3wEokTNXGm9cG82OI551+b4hVP31j8HZZZP5TiC6gstn1HkDzBtFFr1nG
3kGXFR4tkhZ2yJl+0sxdggs8W1dH5wObW0osQRbuyQFmrLtG5IRJ+dZaNThV1zpbtCeKuvkNdyht
/YhK3adBQ9Jhd+hIXJ+K8YpZTfSPEOU0p//IlPkczv2naE8MBTxzbC1P7Cu3LjVsrEAeUia3p+vT
qp1DB/gn21TmrDdKhHkjjwWVGa8sUL1vhD+5VJyPR/P/pkCIQw9Am4N+OoL18wZoLykB8iw0/EvZ
FjvCZ22yzs0HiPckKs6PyXr/6hfrE4gusQYj4kNn/YrPcWnwCSTS288s3s2O0z0A5ElHwIutOyOL
3ckmgrtI38b5Man5cbVBBT/4AtaM2m8tsszo2UxlKxOH838kAr06G11M/q3DVMdFk/eJw798ia/V
eIJduTMwxxZX2ct58VwWbHLyg7gLSbzQ4enkqgCSWLWluFJGdUwnikkP+ZumOr/larOYCLfAmc+V
S0Y8awnQOQrZn6YMpgxOcgYMDVk1BhrN/TFcaCbCypcfUXNVcv3QHSMyKbFSAdXRdND9IoaXHG/E
X+1o3PfJ3MfNt+GMaGyLSRYq/wAKbg3xhHrbPm+GtppLh1kzxY7JsX0ik6E12FtOPY4tRlqccBiA
aOtkDGOBAwm+OiZnQ2HYnVIj98dW9ssgNcRFOM/t275vQsmueTdVWQZgVlqWivkg7eqelnlTCoA4
zXwvizfTxzKVI9n0BXTQIdbbdVfHcNAwVRwoXEOx3M3O7O3T2yL72sb/CVwwhXYV3m2eGMIvSWaE
lzGWB8ee/LP+Boix7b6X88npsbJmHphkTwGUhyMsgd8neEvIfUj1KZyZdFLSgnOKFTELq0RXxMiv
iHO89KUbvB5XhEESf8+86WeGGC3HCIB+MzOOQpJgR5PyzFC8G0gmBS7qaIYy/3UBVKqzZSYYS1PV
dzMTek7W4w/Egoy9Lw17YjCDX6URkXrrmcvqJ3G1x8wIWmgA/cBdyRfOrqhSn6A5kkvMkyg7T//N
14tykCLELlLIK+Z6rQHM/3ZOTTtCj/XV8oGYJQNVxtwtggzcvOITRQ0UXFS6NmU409OJ3jg70g+g
s47A6PV0fnTh2INTI3vFQF09Ps9wvmh11W9rb64Gx2VzS9OdWP56NWXuhigJbX3lRwDzh/iBukEr
yG8jrw7XaqMk/rdT13ybZF8yJokTGItan33UKmnsdrpBaa5GUnxIkzl+JxNTOgDV2KegoGjanftH
miGYE5hgjsj7mHFGhiY55qMo5OdrCsNyr23TRDQJIyYpB2q20BZ4c9tZddTzkh/TQM1Dg3bHrZGO
KGlkDYc7GSK1yTm8n4AKT3PKUBOXauAyk9bv5QW/1iHjRpexe5YdZo5cuJWd0c9aQ6pTlP14sou1
rhQvBEEnH4fKcKPHzto52oKPCJs1dDMvdBrJ2xEleL+ZY/HWnPB9PZ0gqcFRKQqNfm6MEgXlskKj
Lk2a32nU0KKUNL3Cg0il7qW+oJvHCHUw8W18XlM472bAvCnAXUfXHXZI6BbB4FQ7ukPwC2J5kP3M
yF9g8wtQbtRtW9JkGjfMuHew7RuDS3gS6NloERn75/PGCwIKeDuQgPmT+fNDcBSGHrFT+yH9HDqB
Z4tVF5JpZKckOzrNbQNRssSOlg96IHwNIN0Ng/LcKlnznbNpCiEoqNQlY2jvmmiUcixg3lQZDN33
3ICnmW1IgagW+gjklLn+TEDANXSBBEih6L6lBiCSHaHFDkq7qBVIqgSKEZBJmyQ4xyvUnA4obrI1
ZN1CP5ZGeiTGfX4HRSXdgll2S43dMRGRCLfEPvp+y82y4NpHpD6qHCwcde7EFrAA8CKcxh2+L6dg
XueO/E4K8lL+SilGXijtgTG7Etmywxqn11ZJGTacUUZE1pvl1WJ1b5htIbEU7wQkf+Shyqb5WWys
3/k9MYaFBm5SEaSbWsUp0auCj5Yy1nxyM11r1UUcUFLcRA/6KrFKVXKibZL1pHI+VUcf4ch9dzNe
dVavr9lUHLRs0QH2AvJJXvj75qkQa6GUNRTHGlGO7OmXSY5yHpuy2eun/P/kQ0nT7EtFMMDG1tSn
2/HGkWGZ34delUXz7rAeevwSQm/6K+iKhgoVEx7svSA4h54uEIlYNOO0tP604WmkOL32Kol/E2iF
u+GdKHi7W+S3JKyBdYiro0kEEgQXpD//ZdCtOAwBV1OozCa7cX/anIetRqZ2vxokn3gLlZ1DRdoC
hf9a0elfKDuaF92H2juPbXRKWERSvciZi7ixJ3bhl0Qea/Da3qKSlvT4vXjQ3Ay/GCAzStzXU6+6
CiqKLIozs1OetBWymvCHVFZeSgRYBkLaIKKbYcmoO8fXXvHXqL2YHa5kXgCZOLd8754a8h7WuQvw
JuPDuwQaBnQ+SZhoi3SydoGobkdjJZSV7I44rxotANeQHd6ZxAKT78NH4EoPEbc7GxYbM+yw0uaO
mWQr8B2u2vtdnLt/KsK6n/ygRzAPGEhu8jhF1I0bxNk+EXpkH7XZ2tirOP+rZKEkYvCMvt8zpua8
G1ozFHDwvBYiKfEH+bs/EoNSUVkguZlZ8JRHT29rlaEWwoh5tg3paLwllcRYXTa0lhn9gOYyZXva
v/yRyS2DYnu2lRd/0ZBBP2gnVqvkV4Eq/TmvvlvM6dbcrSw+LsBcdxhxh2Pn8c0lBgxxtMSe5MoQ
pJDxNvj4QI60y7uT4fj8/+hTnDKteLTqItUiCPHHcsR+93HuiRwJBt5vpZP6zxTXqzy2Uk0HtJg4
begxwedqneblLCrqR5KKj54m5s+7QoPAYmZ1uQiXrx3TvJt0grJdOi7wcp9+528tpJRQeXos20Yt
UEuSUYv1Wmh1GFpTRnido2ZhjrPRGgmEBr/C6GQDFeDD81h1GYINrkqPaj+Bkfq3s3WDKFd8viGm
HFOfmVGv/brhJC0g4CqovfeuZNWyjs0eZpoc5kkrN7zCPrX0M8mO/k0iXxTD8/25qgn7mZum9r3C
Wnp9D+b6QdZ2O3ZuS5+Ytk/JBXb0WyU7qHSQwej2ilWzewjfnS8xoCiTPqZ4YCa9/PK0UY3gw4Br
J/CPNX3Vw3HLC5wIx0edMH0+yHAYTtzmarDnpsztpd3r+lUY058+dak1WT06cfXhWBBzrC3g1omH
GwDPtH8yGwJnU4grVG4qjfD4NolsuwWa3wBPVfoXTnMs+IdrK7sc3re1PJqQuruBWeH/w6M6bMmc
mplI+EZR+sGqxQqhmXcgD79MAuA2lQ1lo+r/qhaHn4kzIMMMzDE29O7bCBKMz+cBewEt+qjNVscm
HZP8Uh5+hi0ztOj/QQBBh/Ea2tG+3rDuKvxtPT4ItIEBj9DKeVIDLHYx4snVPbx1Ra+2TCkhDD0c
suaMR2vvIHAR6tKoj1dnofjWO3byJNuFtjzAywTHT9JlWBs6sqSforg5Eu4oKJPW74xPtZCAHkwZ
fP4QUzgsfbApby4U0np4TM5KffBfVIttSeYZW4lB/8xcR2pZd2M4VdM9o2B37ApFxPRIaI6NrbMM
uJaB84VMXAHpgwiGiPEhMCTH8GSrI682ciTtrgPyhUiadhcqol/+62DCIba/RpzXx7RoFVe93Us6
IU9cIstHIwPWoOHFdyrinpWL0OeN2cHB72+Zqc+Pwsq67O7usyRbDSZDQbQqClkahQtxlagDC1o8
5EPBFMQU3i2UtZETVnnCEgmWiwONqtlABfcNlLkEn+Gr91c5b7xDWiv11ZjR7Of97L7YV3Wp1rDy
pPNCq9qtGygrmRPo+vib4PmPEaNB4MGi4DTsvzsqNBquR6Q0T1MK5FQRro6v6KCEKdxE3ri3yEZK
OByegvNeWWiFczRqTpvtAfsvtmj5j3yYYDLNbMp2BSoc0pUnHHJR8ixn6ZOQuviDkyCD+wQ5QvSK
pG/ySbRk65fiRTCIQ+MVR0a9zGN3+rrJZHMkg/fS2VwqDthGH+kf1qofdrvbBno02x0FwkKTNg0h
32eqiDHHV/G8y4yPZILZMvBw63P5YRK6+40qhPIUNykM/7KcgU9owaJRTEeI3qKV9C1EwsfxYfSk
jVGSFThGc0zbiG90IskBgNiVtEwlJuy9+3Jaca7k7CoT7D6bK13w+rG5N0+wEY+VAMHP7+VyTp/H
bijJmPnjMqhwvk4Qs1WROjCJtW7FhHkuOBggmW+aF3F1/63WJ/KbVuBYzrApYEwS9Dhsl05oLlHL
7oPU+VH1v9mkDJvZqnDz3d5li/vA+XvWUyqjaZuvX28Xb58R+KMpBZDJhJak0X3NG1mucx7tJWeH
oa0ASgvPIGo/IOk74jVoPvhHIhQHAYIzfPk0iSV19aEExaWS44RFTUrYTou01nWz+BJ0Bj3+7ruG
+SLjOaw2EuaFDBbWYYCt36/Liv5J3//0x8PBAY5vz1/vbdKbn59FN0CsYsOYfZEdP6Kc8Oxe09ic
rf5zgo2KNR3BtwblPU9GEefsktNvWUBELokNEVp5v5UTWo3+brwppCx8GwNV0LMTdd7DQVUZymTy
hvzxDeSDOJBLz+vbVJHw0sga/Mh53SSlTFLw850V6h3xWFa8MolD2OSK74k6AgWxd4ipcrW+tAZs
AWPZsA243EHG7zxIldbF++PGfFd5xkX6iz+AKDAxTM0pj+ehYpvnp6Lmx5hdqTxa4165te6Bcs+F
RasfJKZGsY4x2vwCK2C9veO6gayi2fY5+A9El880rYfF1PTnz4UZZJB3hlacTHUkCCJskAXqLvJB
feNKagB4r8YSC2STBjVlTlzJENcfvapMu23/T7VtTPxYKj/OVtVYvUOr9/u+xGiO/X3DrS9//FfV
LarBjpgNWuKGDE+GBl9KTE52Kif5fAqgyVlst98VKO1e/Yuyvmc1aM1VcXm4afZcoaNN4eaZtypB
gbs0kuNcMCdjpiRofjOzzvC2Kx+G9OWv4q6aNwwepnMxQpEBngQWZyvuNAgqCJ1I29bKaVkxMunz
tXzg0j7+IQRZCFLDTS8LmWvcA+aObvYmtb+8FhtcuPbuX5ejqOYrOA4SXduavzy+B3bcdY/g2CFm
U6AtTP+5+fe0xfjw19fkl2VorT23GN2zTslOVff1iQ8xfWKgwuhQRH2PP9VOas8SBffZH0NlWZRS
9PDI8Ph24Fh7TEimaCp78MdwQF3+KblCGUBRYngsx6UXs+7JEs59AO6DgCdVScmwN2qAOy8Y1rUb
+b+8kWxRXpIUXlsyAL5FYHVzVwLhv35qkgpUxiVNrOXI/yrZEER9SQZkObdBjpEHlfW9w+T6JbNc
0DVCua8C/bX+2Pi4n2FcjG8Y05u/03BPBwKTQADpbpBGlU8n6G0ZyWcaa/aBLWOo/G4eb7MRtuKU
RDlHSOOyQoOHKBUuvHoFCVXmfASkAee2TvJcOCS7yHm4Vh8Uj2UeaJb0aGHGKJzV69M2mCe90pgy
qRstpwdAo1PdWsar39bGF7BXtVHUoWv0gMaiclVWcXj1R6yKjv5+IqtQgRm2B9nGdEaJklhe3e2z
KOvMzWr3MCE22kf+POy6+SdDg+snT90DTv48EAi2ipjGuMPw/r5ndhX8Q3JTJUMUQONNaHPPm/Cj
eCBH0IzOFvIgFyejGaPDEJ8P4hzmiNwWhYqv+9pPtwClna4Z0fCk3rTLmP5SDTmyB/6eozUPwoVp
GTw5awMu/WkxKpXZ3dnP4gXWIrZPPeX874BtkrZ9RabQbeNSSLthuwfZdpLzM/QfW9FkPMTfoYxT
P5Llk2tgdS9CUZhQwy8mwlib+07T4Dei0mmzs1tkIzs5Dlkew+QMDsKe7uDLRJTXP/M706XJJ9fI
8PbM6UHBvHIVrfMbmyD4Y0OLgieBrjmLQSOlKy2PDfCH03Cdr8xNK8pGmCAlT1ZLs95cRGWG9+/R
PlEP8jGnhXMm95ULJWt/G1S6JE9bMT6Fqvgq3b4kVn7kfQWwy8L1wgRtGBSXisodsajMOO0FkbRV
g+s7tIC43IgW7TBdOb94G1EKEE2vJNamW1ksqkCXwPfozy3cOoUHIIypUD+auACmt8KTirPHwYmy
x/AJOcWBSMcY1sd3jYkK8Urx9H2c6mp8jkb1BrxcK+8KOf+92BJY1qrUHL2g+zPVe2VaB0IGlRh5
4dHmRSyARZAqrsYfpDJfK6pTifmlzP2brhQl4zkD+xF6kuOGaPU0yInTGeSi5OFttc2llEB2oqUM
W9e8Rv2MfnST0hTJrQFAAqXEFYTQY8MmhsXB0EHxicMAWKaiQ5EAd86OFXXM1CIoQgxS0/Q20StG
N13KI9V7pEMzXG4DY0dc5YP+DHhn4CMrKpv6mk/otuon1vRhbGtLLatnmDk0jluw4G4oAW7PyIWY
kwoEKoZkmNU6AAQteAMdjr/GruXyPQQmvr4vikf0AHRWKj30rvasM8U8w9ErGlPpGkThjff1H5e8
joR9Qq4bsvdSyStNXXEHuT85MZVYazc6rcKHgx+tdR4h13lbwctOB3lz77jP+wGky/cOH9kN1c5W
7Z/YcwKBijY/4QclgtKZZC9rYj2m5Hej/1PxJ/vAldhj0oeiUcP2M8iZXKYOPqQlF3cgF8Dg7vqn
emWwvzjbiHUMFCyc9G8IXEscn2mM6J49ERYFLL9Qnlywy/vMG2H3v/ad2usTYY8nAgulLaOSnPrJ
eYyEVbT2IG4k0cXFwdqlv2S2Z14K/xgMVO094bg8lQxYpydy4itso3koCRRCKXBZ1q15Aw59l2OR
m0+eFrYUuYnb3pFW5LogETm0UxkSzcuSWze/xytqVh9LktfXq80+Ig/aihYLyhwznBNqvWT1SArw
61pkxld7uqsWFKcT7cDK9QeX711JF4C/3rjc53MkTkGbZ9X4jaWd3U/Axhge3zKH9YZlbE5ZZ3tC
4RNpoeOUpX/Io7aWbs1RWlw7Fx+Hl3jYmqXVnGsbKWviSwDmPQfbpu/BbCtMTKehC9xxh5a9bUtb
Ua29IX1ZJoX3H3VqWloQEOUzSd7fEGFJJ8zXWkxBSTh7D2uMrEkiur4T3OXlDOjXA3u0IoAFF9Q7
fWcMJ2GYqehNuHZsIN7a3MWUqAQbGJgkS2iSi3mu7RyIUKUBDLO09uO8BtJJzlEusD1VENdc+xui
Tpf0AMmVaixPIUJ9T+UuB1qfTtmjCclvaIan9RW7oVDjAhr1NHcL5P52+GtCNlZcZYjR4wYtnjp/
3wd7W9I3L/OvCC833XH778FWHgGeEAKomUbcME4w8x6Vbb85L7R6GQ6gFmxbkeMCcG1WSNUPApFA
W5oyB9jt5NfJJIyCA52b36Y/L4VvHnoESOsNvdIK4QSdY9SOVbeunMx3UrVqivwbYPzb9fki1ygp
eCcYGNzk2S4wFJxYQwODVs54frRHAF8GxPmfMwLV33zxp+gkUGaoE6hE8VK3unA5jFAtErUcarH0
RlI3odXU0W/lnql6nKSrHuZ/Ba9kGPFYpOpO5ljwf6fBUgz1HXtEneajiNYa8XbWTI+GR8tQBnnF
nKsd3maIQmPATO/S7NzkPiT/h0Jc5TMkjcRuFrRwvk5ukRacVgjFBZ7MSnQOB/QBc80tYb6GEpKQ
IwPE2KOGbbuxTlf5i7IqeDbJAKwq3AjnpkobQd8XDuAhqhAr4UbPJdqbPnKUHjjtAriySddrUUMr
jD/J7STg0aqf6MwPPH+fGOatRAHsLWa+NhG8TuC0cyQB0tN76BIzdZZa+AvA8cQjA1HJCep0CyHO
2Jyk8ZBtIozKsCAGTdhUyOOnVpje8kdtYhUDW248R3KoZmBKvLcJrHSxlzuHupeD9yDUkR4hFm3G
PzrErfJjNIn7v6GW3GiB5Anp6nbkYxWhwAoaGmnXe3kNMT45nOdal4PSA5vc2MLQmS+pbpRJpDsR
ikKjuHipEXdGznJb5KudcT7Ywaxl+sBIEvpRFtB1hN8E4y4TDX7vXicP87CYhOj2ZZa/Eti5Sk8p
R50/hPriygCovjKvxPjUVsCkGhZ6JYTbJIJ7i6i5P3QV7U8u7TBsG2O9DuQ26IQAPwwuTtBsioRZ
QQAB7AjXI/HJhY/wUq9WyZo+e05wKyUiUwCYJTLgZwB6NnAvmNs6FAz7R2RxVRqlTYmcNC3MjhPk
8gpWVlW0hnSMzAH351D7zuOQpXBCALFX/5xZjQiae6zl8vi89QR4xKv3t98l1V12Nel3yI1NgAOA
uPeUG9vs5f3ocFqNSl5iEpsMGoBY35tnEscy1jdGwhf7U8v/OrXkzI2qDn1VXggezwwYBQ5aiQLm
AjTcfy8L5do9p+92yJsFNHeSesL0AR24Mb9U1T/FXuKHgtWzQR0zhd8DqkFPdi2O2rZo4RZk6jtv
lu1FXG9BjcZPawhRcSw8yzvGwWt4uQET6v/1MwSCVfGOBEsiMwAL9AMhOX01GaumqPT+f1TFVUe4
xttvVXrxr92od62ZwoHr+NEhWxYJzlMr9uNKzMd40fYs3YdzMyH6EFfRn3k4IpvNW3v4TyVxHkr3
0yS38egPvECeCECNKgUbyEMY6oUTZqhZha/o5I4L+5qTG8fsHJtbh4Zeq96+I5KIPf1m6e4DwjKJ
4mrkZtmr57+WlL8lSJj74VKpUYQ9GMMXOKMVsP3+W4s/f5e4oYT/TJ/taLzN/sQ2AJGjNHAR1yN3
WZQUQLpG6IL2/YmElQ2d9mBN3RrUvoQL2lCZ5Dm6hetoTScXWTKzNyxkWL/5PdloZXPhV49KnX8B
i92GzCZ9sjIBLB7DeuMJZXs1Lqmq718EEwazbePIE9cqcPCkz63Z08kUtdtixS5wQEN1rKWmAOr2
DVmT6TwWbmkyPhWaXnLkd+AOYTVI4goR5O8Gwc46AGdj7nk5wL08VeoMHQ0rXFNj01eb0+ZP6atU
K8e53Rv9dF893kn6CM/kg4jCeTI6rJNbUeaBjCrNs2eCVKk0/70+cNkwS3SgMdkcOIQIOnMFuIT3
2UdMJWkI86LwoxTg2FBPIxowrNU4Aju87g16x5G23XAl833XJqOSbPUDlcPXBQ79OF55xiI8zNfg
Glb8pquv9lsqBXD3LqKWLcRdUfcG5XZ63D8hF/Xoh2MwC0maQeV/vZjrNy3AGR3ymI2Cig5RCIeV
Hgys5yB9i8q+wlV9eJvVvfSd5fhRT5Xk08FlAP4MM9ErrHa5SWjBDxvNpe3IsiPFZT+X/J2V/xKf
up3NySIpnEWxF1rHL84aXBnilKiHa5g7ETtmNg2PDpOYZ0FOjPhYO9ItSxFOOcc2lkuV0cakFra0
DwgMGvW5Z/8+rsNI7scriw98X05cBThnldLLUf1wSl+R0kwZGmCla2mv4DgnnJU3/XraenrFaQGW
EE+UWD2gQIHYNC0BhM60UEPo5SUEY8xpArktGvvaAT+6wo0e4duk9YwSdIH2babPNTjPXhu57yit
WuTCgLrzBdhwH+75U9Hurj2aOaXWVRQigG4FylSdN206D8nX856Gf/mG7y/fuoig7oJ7kBeyjq1/
+O1UfG7FWOBFEKItazi49fsgpEq02VKNDdLQQc/ABwIS+ESupHrcUyV6ywXEdNynvWptc5tDtPG8
8YtdgkzBe8tsvQO5hVvWX14ieHLgTOGGYjiYB1iet7ZwJdbWYOZR21qwmwmyrmwDLvS8z1afrmZa
UASNXC4PmcVKdKcKqRe8T3H3fYFw+e2ZK9vKnFHnLdX7rWxat5puQ8pFRbSsG+RYZeK+1dqPlLgo
zTBiFKK865mw0p/0o7MtcNKsWkJEX9ekrxMWiCJvaapwwGFaenNx7s6+KygC0jG2IoQK+3le2pWm
3QwZDlKedYIuaVcSdXkmDOSfAsABsmnrG3HmgC5CEUAGwF2aCwf7SUhbbsX7FGNagD/RS705Tonv
kTWH0uCKBINBgHcBJWqUuvEh3pRqZ52UldfD4HbTXaAoPYFFlsjtyFj/Uuc6QgKgwZZt3oshZAKN
lvXqSuoSiCUd6NI2tzOjvGxKZE9dsYwqcHQMTRTEW7mTMQoVk0BIJfxyNytuXJqC8IeP03zbxzio
tEfZ8ZPhUN9K7ARpXPh2zfF+rpo6QiugfzPsqb9fDyvcDN5dIed8pIAId2rGCw1vhlI5U0YcoEV9
8j0UDOscYWocDPRomLLOZWiOqf6rUyvYqzC4ySPLV77FkzH308B6+fEEPZI9ZxJKjeegElr+x9Ma
LHvxLbGbPwyW1r5Jjgy1fTAaPBP7tNPNWuR2dnMK37aZ7Naaqvo89gUdx404joycM3mXp9xchnw2
7d8E3sYEm7mCCy5hK7ivdnC7RQxnvQwMUpEq49ge46ULXFR0LPbkTlS+jtJgqst8BloTFbQZloZR
c3V7u0iPcDAjxO97HF6cQYwie/K9hB2DWRB9AQ10MqEHM1469tCjW5LuSheKqRjbWYTPJYyI6gbr
qytliEqrvvV0IQi81Yuxh2iKOLxJd6l6HMm8qvMt2GToy8ryWh8KfhP3Fx6hid7erHFgR1GQSMXo
6U0zSOyQjZuikKmhVBA6O/v7fcYZKXKXF7lT+38tbhuUj298/RTy9WQZMI5mCYkbojwiyo26JPwj
by94RfcuFVPJNFckhc61Ufter0gT7tidVcCZ0txuStk4ZMy9JWSPW4rRWiFjtmAOmigR4fJ4n62q
he2IQX958rQqO/Hx2dg6isodX6qF1Z4DsrfJtWG/+dAJj/XB4nGoHbrAuK+emYXYISXcDz9PFz41
ncY4LF4YkrNopIiYfgttGvtGiNDpZfNWcOApf4GQhw+jv3cTPjh/XVNDh1auNYv7arQ8cmt9DmI0
aggVMRo5G/nUCHeBqPxDVK1SggUfoy75XJDxrITkttcxqw7leje5GSlGMn3CIX7T7kRJ8SBrWgFt
87KhEueE2kkU3C3D3yAcK6KGK252g5STND7CuOFoI3KG9DQH5yFHpP1xOm9DvwCjMcia/9TxmAEm
NAf9d5Qe3HOyjJ4h+F00+JW0F7amfpkMYY/yzIQvxnPGOsW9tQ7XpCNElQYMM3kL3MW1zEGsUkEy
NDMJpHcGTe5bivytPxFHmPKSv1DwRWPslcVxXgZzV9m3gl+Tt8ThkDtpKlbMY4IiysmnJArZg4LK
MXFeFAFGVtX+RajUiWl3mnkHVEcxmk1HHQcOcIQKOMUZl57v9hjjJUbn2Yvkh7DH/y0JYITlHBUC
ItuOZkkno3gNt8bEh6Ux5L2ZSLeN81f7KXVqtrfvKgtg71U4uNUoWFzkuZx6sVgGsCy9IwiKvlc9
K3xOyuavD3OU4HovVXBiFtxfWZNhLCS7+4ViTf7yno2rX+p86+6haEOl29z2ww97RBNeu57DopYO
k/CH1FRmbw5FxJ76FYHqjY6w498PEeRVDwNHrWXZTX89Ev71gtIQJ0D0sEwYCH37FWtTk8kiagZQ
QG/rbPQnvSOE8Yk+eNINHjoKumo0uQyUi64W0pQdN4L6EfYRFzBGqdkwgdg4lMrtXnPJIUa5rfDo
/kHBbiGvKYg7Bu8RGKL4nOziZU7YDCrHSb8ZC2hy1pBPls8Umnb6NVc0GRo66V2AwXmA9RaPRa0O
scAujoUgc8IJu5muKeGaceiobpX1GXEMkO6i1GLiAvwZwUv+FlhdzGRgr9CZ3c+vPirXAJF9+ENe
7/GX/O48HxmLqAE1hHll9cBBCEC2QNoouptcGCKG6dUpAZtC65MT5bBG4fbRgpcKOERmSk+n8gEx
2fTOwVXOALjAmm7c7INwlyq07nfG7ZDz8mTSvro+ra7dwSmvD4LvSVl5pUCtmzl8MLQ1hCIyxu78
CvW2YWvLNbrI2PybhDG1DgMWfdvoEocIEi0pYFy8cE0QEqmhnqofAPMkOb1PA5O9bZIt8ntR530/
czgMfEvwWvVTjzpRbQbMPskx4vggEl38o+yU3gGr+VWRVCYsQPz6VHbdxPn93s82Zvkb6HtHT8bJ
vBL814DcqTdAK1khL6LV+7hk2HL5CetXTD8lQz/dq+CeY3e0f8ZsIAT9DQGZQxJQYRybJyEJfD73
fVANe7KC8x7yp1sgQWG8rj2N1+FWj0bTcAhlHzuywxbB2FS/on20kportPps5t3K3lcDzW/7xQj0
sI/cnbRkfFdQWLbMnP6hKBuJ9qqfo3idh2LainDpCZGj1JkSt16AWvxCyAYAXaswNR+VP9mpBqYa
hctmYegTyZ7DrdxBfgx/0SVurYrp5HLaNlQP6IZOTumrtgWZloSQwjXywx/YaQRr5cq3GtE8jjTC
tFq6CWS4f3K6qhcAfEq1MF+CMFsE0Y2nwt+LtiE0MxueURptItgjq4GYcUOovw4vOo7s8fLNEx+f
d4l8TBIc6MsOhvXJpcFXQ3ubmDkA6yYRUlrbpma2UdR20f0Qe9xdLarsDKMmqUwLGxz00oJhZ9+3
jAHhSN8TPmLRRJGzaEuGqDqBmSIZ4kjcyRnpWZQwHgZKvzyrRDfsVIWP6L26iZ+oZfnIll1/fI4I
EIBbqwTRsFmv/CRUN+CAIjjoA/Z2bPfJUuOJPvjoBDi54rTLJl5aQZq4u326Jt2XrVatr0qz/cM1
HYuou4b6/4CXFaG4GDNoMqaTllMP1ZzD8rxmUvybL7BPEIdvtlYdkWOkbJra/2GEydOYKE9ILezL
knWe0Oo8YO7FoI8PGAkQ/D1XI82d3p7c6pFRUYUFBdvAJbAmKtfi6NRKVA3uUsPcTGZ/Whk3Au70
hXvIjeAlVfDe6LimQSsJOCNUCmoE18b+/X7UC0J0ARoPhChxAfN/TnttAgzmc67pGvSZ5AMXOAit
qZ6u3pR4QIuUkA7b9Uz2PnmxP4L/xOW2Jiv0WosEwWVFCTsAAws6AqS98wHc4Ov6bNHxEPZA2//t
DiNxO5KFauHZ83qTPlDH7kW4vHlupcRJLeAKMaRNyVLrUQPejakmVt6InwyDGHU9/eBrNf0EpR3V
tjB0lGI0ji+44U4nW5P2r8xOw9YRZkrocWgQa7c3pwp1NCztVPjTm6k07I7u0cVkjQhqAMUTeXgG
y+2bLsQub/c3jgYMwbh0BHU206g+y+gcoimMXVukh33A8AiCeIudV3erzfnyyhEsq0uNu7B2mhu8
y2BE7LdeENkOKarC+qPWpV3B5avp3+t9g3/AZBkLijRlxEu526jPiT2fhoJF9Th6ycuEX+Sp8AYo
EcFzeIAkRKu8nISI4y+vEYBsc95VjrC7ERLh620yePtZ/6SdflzOR5qHA2ReNvVGj0jY191FaosI
ddYe3TFld751nSxlV+0t7S8qK2lDxvgIiTFYEuMi5iTzBxEk7BsLRg6HJOK6HKCoQ4SS8wY/L+Qv
Vvu+8wJkACjlRlXgUrqqIX6YU9alDC5z367IX+1m1XUkt5ZACZdAC1hv9uqDUE3YPS9Hg/ArgHtI
Bb/vH0RoDKJze/5VI3LMiUwctWCWsrmE8i737p9QZhY8osws5BQBVgvAE9fiYkSr1YBzstiI5GOt
+6Vd4+7fyW1ZnZuzzfwfIGTfuCZTaJ9eOLr3zqYBJ4x9hNbZL9wr7htCMx22wuK4BOljd6ie0nA7
mH5tDhGiJiVNiqZniNUyjxtNebVIQ4zsaO8CxT0WnANM9GO0Q3nsG2+vCoWAtMWOCjpAQlij3rNI
eQS8fHwQPQujDTc1Thf+/E/OV1vW5shKiYi2eH+/ofGrb2bFrKMlxHYEB9zDmiQW5u2zDeRuvhhl
6AYnkSddxoeVg5GSKbeLD3L6MFAZa1a4VAOxB0TtQJcGAA3W8u2mUwf1+mBWvy/Ey7HbtwBFGaFJ
XrZcenq7CS0UzcG5n0/d+aiFiiQNDH+c8ztvSP14+JrcTclK9vIejEwpUjaVQeDX26CViAgY5OFL
SnN7/jAC9AiXn/rDePIV8ut0bobacnvgmridM4NAmqVJ3DZi/fSWS0QZ3CGobzmhjf83BJNOI3Pq
vbHzF1BpG6n4Z4uJ+u1iGjldZnDF+7ZCggTXYDR8yUlQ3/nKGaOOFmJcMFAbE4XNyPAkv3fR5hNE
9VH0ywuW6guBsVgyZkL+wMYmZO7u+GmEc24dfo9+MVEuF0V/viCfg/x7LTqRjkbDA/pGugWsFeeR
shDoLrT28k5Rr5jWw/X5yYk8qT3OLkMbElA7/WtZNQ9/tlg80xZJrd/1XgxQM6Ju5AXOrQg1erVO
PqO9ETwh38ScWM6J0Mb2PK6hDqzSDTPE0U45rvtJUY8ZU8UxSSCnhqhhYJ7fBOYwvZkYQcyLKe70
jdinWWjOCMqTxweh4efeETYLyyBuBIL63rAVnns+P9PhtYw0KFBPz1G0bhn+nb2YrPsN4CaxMppF
RWZQMrSVRadDMClZdzpHr/o2h+GDcZTacEu6xJA7CM2njuVMK/mymn1LH7FnRMfJ2tFkD30iIP1w
DeYhcDVXSKwvBBghAm5gUTL99WRvAYGicEg/UxrMSLZYxGIe6Jr8XbFFYGAtXP4IG56+VKGm6E1J
pg3v/fPzHQ5z5VWK7W9TqGI9OWPBdvVg9OrbOr8svKr2buBNv/CLdorc2v3i1PTDKAZ2mjOLdiZF
qnFsqHn0g5uqOOYuL2WFXhk7A5CsnTpOOt+XLFYPujEahy50sOv1k+Zh94nR4JgwfgtLG8gARDsY
m8AgSBA4Q4DiFBT2WWCJRgTyk5WQoYgmmEmMmbKfUwIdx4Sr+x3FRitD9tu7R7Jy04JkIHqyUBtL
VVQBBpQiBuJsf21mMvxefnnwYBWeNRZ1x+hwswgzvxbN/gPKnMWGNqPhhKHU86oStugUhFjwu1O0
x8TarZScwjv7zp9UpQeRtg6d6DnLLzD+tyC0qKYwQSGSDkrwYFyEqR8uJUERU4sYn8UGmeJdLafv
HhNSXzzirA3pf/VFE9797mYMzbJv9jDvtQtnyMrgeVHBDf93ztAer2qqasKMkSmpGIYxb3lpcgPm
xVUd5FVgKCB6q4k8suRNiUbP/Srfkcu5xL/YCTNUsJgj5RizBV7opp7FrmkKvZ8m0oKju8OxHmy9
6UymFOIhpLLd8JFXJ/9UbmEWOCPDX3N/sT00TJwEPTqFz6udv3Bf7Q+m3uw75ZrbOz5Deywr2+gz
qkftoTthdlyD5GbAN0aw+rcwBKdAzP5VBkzQX40VEeQY9o9+n5bkB8q2k5Ogl7XW7AZ5Xzf8NFHu
Ywa7Q9Fw/dWqkm8+s1qo7MrRVQsYJnZxp/hRh7V35i9rbL24S68rQBGDKSrh/lKRX4ZNSUZ578oi
Dwgyte+VvVBbSTrDf002CLcxPYduOhy9fDlIZatMbfDrM+muBQxYEZrAmNh/cWI3UpdZHgvQV3lM
UaE119owtwrusUWg7JIdlgwAKV7ijYPIm9FhC1aEnSQlWRkL719s+x/uSw4VtUIbsrh1qsiJXSj5
ImCURLrXENiNjJ9CblUOJTBIMmdJPCM56cbq9Rvfi3XQJugTblHClDt30biWaNQZDJhViz9RyMYA
HlQQv3+Fi03/370XEHRfjk+/QbXyyMdp13GjeTImdZvCWRnEDVANXt/SUrEaPOWV1B3IpzRhLixy
a6d3Z6AsRjkKIL+YiaeaIbjzVmPRIBKjMDuzPH64jOQILneiB4UK72l6EwEARRiYT8C6Wm3uQ1sY
DB15BGpo/k00jWIVTa1+Mw+ENWb7+aA8abtlFyaGv0oMJmTh/U5MbaPEtlEuWVSg5NhNp0tQEal7
BWr7KykJ8Cjl9S1Rcm3Lqk5M0apJi3WrX8cFKyTjrOTXwO96TQWox69CStmNRYKA6AD8WUbKfQxc
sG7cFeRis3yN9wLr+f19oHWSCQK3PseIQ/bAAPdcE22N0FPQJCc00zkHKx3DRtU4/CjwxqQ6dbpi
XYNoejCOdH/mb6O7TZLGTfDGiPjDEOHRXRTpX5v/HbDIJIUJQ8xYlXb6Y9zNSf9a62pieqZ4340z
GB8hfJiKBNfDgnrNxP6HRytKUthAAPRVBAOoXNMTff/J67H/vVIhXeUM1ibQjHkZaP0zkLEYV4E2
/3nqXpU+LwfWm9IelqmT2VX426ufXsD/8/tpGA5O+oBHskCzDeI1U3maDdEygGEOH1zo4wonPqNY
oHKXChum05TCY/HKEPnzYNN0rWjQJJ14M4Zz/hAezRj8ZB4WKB0gTs1H/KmOkPdwG9Cujn71rJXY
yRAuyKdGJ1rArLVEVoJplscS+chqlgio3I2juPHJ3OwBr6oa41HAVRaY8e+iPBqfCCbeEv0BUaOn
MO8AElTXdoZ1XNS1rkxCWIw6z5JcSLgLIYLc5VzC7DYmct7nyLxSL8jG0OXN6Gia22OqhJ1+ji1B
7PcI/ERu7C9lIXsW2zv4mxspVp6HHg4jprwhV1P+gQHMWbH6UhNm0NvG4hsVShebvFsr3sbSnSFZ
W7PkDCT4sQu41shy7ocr+nBaU1bG0nNQP8d8lW1wYu3qc3QOIXkjIP0bIYsak/r6Tu0F4ZayCDzh
NAU7GFkR8Ni7y+ei57wVXzM43aKqJ4gHo71i3YPaL6oUGXIWaBeiVBRVTFDPTQKdDjDFdxDtyuZN
KISLmvJXn5AGLzWQ4XZVdO42XC+LIwpnmwisUKzKnnvzD2Ybqd9lgM7I4IfVguM896ISL/xOVPKj
JXWwTmA4ZnMVQwplyT79FQOGwdAc4w+WzQs8qxzFuokmh0H14ccqKHAaxEXSvF9AZ8h4bnHGXisz
RJuO3k3W1AjwIiz3nCuuD1U63BcIz15G34auR7VWmxpoQY1TgMBKpENuFj9Z2E46ZebxOA2csQGI
CsBP1MWAWubjpYOeYdc51zCAmhJssuNZnDSxWshzVbnpvU/NXklYMkoBRJJDxu1bsVeivUjjiK7w
4pGtiLcFOZFyx0nazjWYjeGqXkjB78+lr3A518GPRxKBS75mRiwPhBA0SVr1YZ2usOCTZ0RQwYwZ
MFT+SiEC1dKp6d3J2f5GEak4hsbDnsLU0aaaILR7NdaC+LVsKHT0ogdDmaceHTqUHSZNvSENobAN
d3CaZPnjLPGZnztYVh03wxrGgnHrF8c45YKBF/EqZeRoo2pjKXvbRSSBkShXXxYz80meSGb2pi7x
YuEuk1ms4L0OEQOZdZv9thMRRGvmI0b+KJMlTEKNPasnIvszY9XO6wxw5IHfZzF1BGrBAzcN8Hzc
ZK4j7vH/nxvl52EQ1/jpUGh9p0IN+5EHC2BK18U56Mzl8TWzcoeLKWteEaL7fHVMr40Tf58Y7wxZ
OCBUZE14KIXN63pVxGPiYGJ5fzjj11EEX8GWEF3WU/94uY3tDW2jNccjbosrQT0pZynv3bmkbHLA
pqStjWIbIsrbKP8uykRmlhDulKLN+OO/NbqXxl8Jw+qXwQ89zLvMd0XshBBS+ny7gQz0CSjTv8TF
7yLswuwHfweFpTiDuT7oivZrKAH2ETCPK0L+thR8tQnRO9/Z3WKfR5D7OC6Jb5bed50slvivEX5q
6U1o3ZSaTajw1YCntAn3j0cCNs0gqxkqC5DkvGF0tSt94+Apue8sEY7qO8+PKDmCGRqjVwMZuEZj
wg+jQa6O9rAThycxBwD7WWtih4U9QsNGuuZmbXc7gFg/g+Y5mYsmGYm/Etw1tMWfVoHNv/+K3Grc
XECSHSdchLAhtN+4r2w7r9dF+jDwB9h1tIgywsmZMtW7QvsfURjs01Qau4ZoQh9I10m2G5FZYcvk
UKaNqfgSqnmgJ0YZMdYG+wjIN6c66YJGTLubLw1/ixFY8EBiYrn0KKjwAoo6jewHORdKTVf5byWq
QQajXFKNQcazaxZvqef6WNfopaWL8AdipNiTzpj3pisN7g4LHoD1/voQlqtNk58ga7KXQl9TltXH
4JaFKXHVxRIzk0o0mzG6Kn/0QAgfDL+p084MPz+7DBH2AS8c2xlPs2zKmUyV0B/+s19MCJlBTOaq
sjNOZp6UwLkKlrZvS34uiGfRCGR6N7gVbkoIOoWcUhMgxILUjsK91Yw714xeDoceQCANPyfC+oUr
ciU3Z/pUHCXDJBh70WHE+sDV5dgTsTgiLVNcoAt+okoMMdANCkLrF7MN3IDe/4/wca/6Ilwd44uJ
v+3M/XiAfghHVnl1gyUTb5TKFm3Qvj2CUxKWUeB2sSmo76f14eEAObCeGaVp/SbkY5BXk0scPIEq
fDdAAq8qdiiThqoTmtdzXOsh2YLMQguw2ZRO36JvNZQqX9sON+6RQIqHIRCau+H02Ds7zglbkPBC
8Mmj5cBOsu5/HzVdvdtViS5g+bQn1FwEr+l1J1SaCfIy5n+684nrlXwnt3yxxZbUDHAkRFB2G0QF
7m6axPZ0NKaWsFI2WGfY5LXLi8KVVDteB2KaosNN3chzSky3WZICQK5aIcvxtzEJB2bWwyE5E1n7
Wx6GYeWKPkjX45Tr9obCMaDGH93O85mJXMfkQaeT9DDbYzbiw0yl8tm73nRXqEDUj+PSnykb8rof
OoHgCG4coug4ITSmmxEQq4yV0yOlV8U6zhWpCpD+SuwbBljistqX/+GVoMCPw7XJ5vO0q3Wumy0m
/GlWMGIIeEMnPI9hvjOg1HP00m+CXLXX6VdsP4WvKtnQ3Z+0FWaO33fP1y5T1c0o9nvcJJZH4ViR
YcECbMB1C+xOsL5jm/O7/6+L1A+7d2JyUZ35yhO0RPNbCUzGkaeNtmVLN1T9jvLanCp+QFgk0eTG
PvRyFvmQVzQYFeZY0PNB8PFfmbizUp399C63WULQtw8LJNX5EfPSu6n+cF6CAVewcFZanJafQTDR
VAUrECQRT/dZeb63UWc3D1Ga3fVwh95qm+aQiBxf948Y1uPOSLXcMxtPOxrx9pvJB9/Q9c3OSYys
/09q7gIXvHz5S2WCaPwB4lgUgc4+8SvIIcqjpqPiZaVHdz6vtDPF5aj4P7nEviMLuIlCR+LAHIMx
xRcV29r4PUw6YN4VDDMoA5Y3s35DCdJ/zMwOZTat6n8+lPjuPb90WoycE/lP3zb+MfEjSAIgOIRr
sgC/B2Og+ZHrG9DC8WuVBG8EPipqHhQ0hnNoeulkE7nz0F5ga9mayKLYBzORIrOQkXgp4qpPpgSn
dfrTm4XbXN+JpHRe4vcVaeQwT9yl9Ey71Dv71HylhvTsLdMdhhu5Qz1spFSBm0abDCM9+69LAns0
1atOrwM5P5ajPCe63KE+QLs8axhoxdypGLWZD/ie8N5JuJtqZqh10JmHL53oY32SKWPgZkl2VkQr
/xZ42Ki77vLmQ5TjDNviRzPnlLA78XDidLT4xTnzja1jQexyCXp388KFuahIxypG+2Pg6mYhJfdW
OXam6eYTMVawL4jrYshUBoBSQzHC6q9PtikiPDKIDpMriwOzWX8rBuMvlTq1BuAp2S4U8qPZbddR
foQNaWSXCCPkNxi3hrTh0jSG1cHASclCly80VnfgoPxkh2hqrfCxpAs4i026fhQZEVZ2uYykHQk2
xAUKVP984En6aRtRC+JRgUKmpYj5P4OrL1L5sfN1HlMQEcrr5BiAkuXjqnnIWi28YwwwdjQkbVTo
1dUy+CXWuD/Tl6oI5kxsyNntjegUE61InXZuCWmlvcEUEstgxnrGOw7T2GMs59B5R957xChqGq0E
c7q6fb4dtN+q05iNfx6SEBnm7n0u3NEBglwQp3rHFZVHNGM7iPU8fpWB3/wjPHBbKXF4yZQff2Uo
kqpobfIaQ2g1LEk32ntQhwDvSOS+Nwu6j7ddBN5NAmkKa5OdDU+aZu8txEWc4aC0QMBd8Dx3v/ol
04L0+jCwamjgXpNfV07oobiYHGhO98XHUZ9Dp/9V/9I6eZv+T7z74s5+Ho8wcFjzJ4DSGAN7VdY/
/WudLznEjLTmbRQFw3VnSPfLoL/VbeOR8hHAL2vujYG+qd8F9DOhS8x5Xo6OIogKIqA98WZhjmsW
X3ETyWS61mqdkLvpyzc1kNC4FdTYLe0G0zoLHFIM58KqYFdefIIr5CecYReqt6BTQj+iDaPtLR4E
Eueot2Fb9JIxVy/BenrN2kNWDPG3TNEzjD/TrvW6oZU/5rLBxoKFdAHqaFVepPdmCx8NtosnwS2g
nUHHFUS4AmF17fM4pZH2HvxyX50KkDAmyIahUm15ljv2dU53Xj1ynQY94Z928O93SAqVd/VvKRPI
JGWlMtc6MHDRUO9NB56exGTM6D4zaiKg8I7BzJwJNDAWDeImTyJFjdQF4+10TiXwEKYnGLI3b6xA
CdRgj4WPaT3QeaZkWkvEp4YO7ee5SP+HjSyNuYPUjam2LBA2Ujle+r2urcHax910pWLgw8nd6ESh
oa2bR2ywp/TUtMbVyVGiL4O43ko73PYgOFdjLruIqrNzIFxVk5u6KpCYZ9okGObqo6GqdFDm7pHM
+Sf2vJq3lIemY0hyF/1BKSpTJu+06q6l+tifIFXuS3yDNAECoV477GPqOsH8apSpCRNnxbzHkpMN
qC/MCnTsltKysy6uZpo5uaDn5+WYgEoUwq4eVzh2NO1THGJer2/VletcOP3kbIqwhRKpe+OzgtvI
rSPGHhjY4CZP8oxX1+npAalcXx5GZZDjzm3dCeSPoiiujNRz3Jy9doq9t3oTuRB/v/Zu/Fg3TQwT
dVoKKfcBIGaoZzQ9CMTlrlIKVlWF55pLF07I2/Q7vJiEHlVFZhuom4EzNcnAuxs9Bj+/0PVnvH1r
0Agx3ZT8xXa45iHLk16Yrr04BL0yQbQ6B+wCIY+M7S6q4rC40vh0RogL3PWx22twJChT18xyj4jl
e1NN2zHyeDlh1VTcKJp5JVao+m6scDsBWmHd2nS884C0Z0tD9RlOlYzfuTo+qGPz1bx8+8b0s92G
MFqFm3uQMj8Ppy9GlOChltFEQaL9pFdUUQgJgMA4ytfB3Cnlb3dIvJ34ow2W5t88sQci1PZ/nbUh
Gu/u+v/Nh7mo0DJAfBqYywGCf57Jp0js54ciy4cROKOaf0B6yQkl/dYP3MCabfNywdN0bNIalO6C
jzgW9+3B72opp/5W5xgxq3hhoFadR1DPyccY2yf1cL0QKkbn9suDtYRCmux6bpBt5IgL9kAr7SLB
ke5x/7xMdv08kP5dcWzUhyFNH/zoTo5BoZrcDl6yEgj2H2F6agq/G5v7PJh6EfTBvN4k1ctRzTEI
uLekaezWxOK8VUtH1xKIpQOA7a7V5o/7MNqpC0uqoViADkumYat1MIlSjmRT0qbX6EIOcvalyJY9
4Jyks22qFfSZOSM+jJf9aW8Fev6LxnZ9Jh21NfcYcaE/dHW6KdDmH6K6OWDysNdVs0KRoFn3O0Z3
QEuEZ+JHKRUn6Mh1EpEqpQrkhTiNuzPMbf2F5U+S2OuwZwtNfKl0mnVjlELX2xSHKlfrrISm1KOQ
b40vOrmPrpuTH9eV8w77ulqBFBPuJjBno9BAy/VZ0kGClj/DABoeD+ATn2xva4I7YHKWtEfH3HzH
QoPxH7L+zangmc1f3SPbW+5vU8e18ZtL0tIHRP0AG3RQZbBSb9nzThwHXRMToMrP3qxnDU5osPyo
pgAuWIxFH1sXH4q7R7sUsigmSuAWaRXPrBz7IaR81xWUfFP8y+hYUQ7PCBR/h2j9yIH1hQnwmy/m
yO4YxYJpljjhJ5TgoQ+wZ0z2aiIJ+s9TYhgn8FYx//+JLsDjTsHkWSp/UY0exGe5QLZ7NlAYzmP0
4+rVWngLVlRH9WoebggRt+uMrtQz2Tw3374VQmgNmJTen5O+ib03jXM7IcnYHmM9e4scM+AYC2Jm
xbKquRcuhTdJxtR2Zip81/2OlUedHKXTpbttu3+A+t0BrCWqZKL1NmXV46kgvGkwjVqXK9vZTQ7E
aXRGHj+OsHZR0wnzahFcRvjHVPvWavhZbrmZHzW0H/b1D900FL7wEmkHcoA+7HQQP61GR58NEEyr
ocpWUwXOjsnUFcAeCsy9F73fxlW0jleg7X7Ifr4lM27H8E3gVbsJl7VjNE0O8NB2cTpOK/z2DwCK
aiIaUTnjmvIsJpJhE7qJuyNziLbd6ymQyl32HOF8/GHQR6VeOm+YeEQ1kd2yHpdarrnUN0HH3xRm
kshsu3VQ2T+YuWRGu5dpZA8CZbBGITbv3ygzcSEjyhFPwz1XbzEOeB/78KtvFxot7IULrKzomCxc
OEoQGl9FZI95vQnRI619ec3ahwJ7LiAKa/mjEEs3cvWomn2lChZtsAzoxgH6iH25Tjuz2Tm4eDNW
6XiDlNvcPtplmD+oIOwIrWnCb4LAQsTh7KwMZg9wRmg+pQ0BTMkIOTSpSrBteamx0l/nImzpSQxy
yE82dtVdxa+mpQvpc79uu85NaHxupHM+pmS6VsodJ3YyfWqBoRjY3QjOU7kK8O1CbFM6IIlIwkSa
NFA1cqE+6cvAbrifGkYNeIA8GJW9P86Ta6fVmnHLa3oJ5x4wk+Pr38Te6497rR1fqLXsucoFCVAi
1L9XTwhpwzeBptEx5qCeNGvBL6S239GJY0RW5U5Zs+Y0TD2tTc+BDl+eT8gSAwVRH3XH87aB4/j3
D8kjvQ4n1yHtu6stbq5uANczvPCYrVBbtMIlz0/uPlTr3miq2gDXwN/LKcB02iZlQzNIRYA0E7Ny
DjgM+yGfWCEAs1JmUq3dohPc4oojjUZRSByBFsM1r4CivY2rLl31pLTWXdANAh0mbziMNRtrbaku
K2AQY8GRF6w74zBsqj2VckwXxasaKsF7MC5aMkbkCzLyNAxpczZkYqsab4PBn78l7UeMbRN9NHd3
bft6tH4OOdcorOWoIhDuCRjqJpbVXfCGIKzgZNtA2ZRGl2sd2hV4e/hezapJZc9WI1pgwZ0w3oBG
EeJirdUU02CUCjEgJjnZazagEZ2oxDJ6OBOlnUqSFI/tsOApzUQJSwgHVoR+mA8lwT7w0bpKuBBz
WMfzIuEqPoV1FeZONdcStLmN/uFVqE67d2iFGcaZ5Kg5Tf32VWMHOKtOeMOrSm44LADrQIWVzKFw
eEIOnuXadMC1qL9VYXaK+hJMWCZ+ZcZhFRtowpnCy2lAnTnBujkESlKpfmZqRz+/Eu06VgoLmQoB
Jn1imhXQsVyXfMLpbDivueye2NulvkNWW6ftBbnd7SDrTiOZwebMeSgyhS02WAqcUlkUsBgFbjVv
VJciRGazeHriaI+p7e675a0OG5XOSBBqMBuNKCqzOcKyu0zzTyNm64t0P7u5Jb4eKfQdr1y0psAJ
rU6vi+kvRTRVAhkXZf4D9GWZoySNWaRQpqb0xbev51ekQnr+85nKPIaZU9JTZ4L+RIx1kcHw+uV7
kFv+fUKk8I0heHa0zsjpfoIWzfqsPW28oD57HS1YnReXZd4isVrN4+03iIqySGsOEm+kw2I3npj0
XpldOL+WFwlAf/BW2IGnKM+d7aQ+vhSaGGbpVuafBQ+vn1xkN4Vh5B2TryqJhbK3Foms3ICLOKRz
HltjQjQhRzI4/rmFLO+Rnnt7LU3HS4fhsnT9jo05OXph05tu3EyWV5np6LtX+UQJV4tNADEquNun
/wI/PBGvYASyUM1r1QVo+PZ25JOBblwUSqeWx9hAFmX1Bf9nqQY9GkeA91aI+x7cR+snZEM/962x
m1yv2dPaulInFsIOUrCCryxCT9jTyJWybphZ9ef+mc6UZlRSpnzgUp07dqJ76noPDaSJkZICZJ5y
K6qVKLEGvlsGaqIYsl8gt3FAb3iXZEj+mi6WnlGoerKDnck2p5Rtv6l9FuB39Os3ekaqHp0DkYzE
QZIa7MCrw3uJRU3p7l9ahiNSiaMx37GjRrouq1T8JKFS1G+jhiFSz8S7MngolhhOcCrZRD7S2kWV
xJDJLIUxK4Kzfh1DNoyGbjTIZatYPBCyzBuxlY6W1GISSb3qDuHbtTHFSk0v75bP51XXZz+Jaw0g
XRYlqtDfE28Z7aAREpyUo8QmUOQxWBQEV8JcO5Am5YLetykKDS9lGSVSgN0EH3RbqqPrqnqhruIs
OklMUYooB6bL0C3+hPL/b8xq0AOujI9adtFWdUYI+RyXZgb6D71+WevyRDa4s9sbu63rKb5Gc1iB
mE5oludDk1FUX1zwq+ddyZQhkxaGY4cOINbMuwOKj/1r/DMADlEYDSg8G6FnhO3fOIz9jG1HebO/
raqSDXmpyBG4w8G72o5zS7f4T1HOrdYMk6Pz3lCftp7+tHdhRJXmBMTuSAim2PQ9+gXMsJDngdaV
Nxcav8l/NNov/CgQ+tRH0fkqPQvwhNcoq36/WlNg/c1HCVCjiK5lN8LHGLmzS7FO9W2lOAlHNi8p
xflHS6d5UwJZEpQYRv2ePP9XnTjn9bwlWRQN42+EDY80mDGSMuV6R24gS0W+Yn/r3SSPthED/9Rj
K20ZX3CjOWMkZHCOJWxfXW50m+RoL7FEWcdxeBDngWR42Z4u4sps2dCOpS+ddW84T+oSN7GMNMkr
9CvmoLtb3wVG3gogAfxrjZGR7ISqWD98GFupqFl2I14tIVgCqQkEsaZjLE8yuWlmKLlJexFAVBNb
Ho8XwP1kVFtzYdwgghjtCJfmSmrdGhjjj3VXcGRxwfKKevnV5MR0wePbggQeiITyqWGNriuyLy/K
8ft6R6dTPxg3k2ZFBUiPhMs7CIVKGObWpawky62FB/bylFHHuAh7JaZq9WPyBTRYk8TDoZE1j+go
4XwWncW1/5NfgsYFtqroaBtTniXCd2hmZgOGzT327Ga3hgKgQ7kaKWIAOr1Wva9xguCJJ5n+5JxY
QjTKxauGHXDva1XX48WkIJmFGaCKWKDpNSwF5AxHEBiuGW1QPdNA8QAWLuJjnUP7j/FVrFYNcGmX
Fgu/QA+X0KJeH5i4O5xgyDfvnh0kExnUzanXDC/+A9bc4nXL03zqa7HdGoOAEAiDmM32yaPmP708
h9ALeNjjC+1nBoRZkVKEUuBukek+eb2dWro0RlgHcAFp4Q1HcOKflMdmJqEEZ2JOgI3/VDlRNbos
PUeCrRqE+xYJ49imM3THbaTzTagyUa9ExQyWzF97szURTid7vv/hp1FN4t/0qBedPxYFvEKRKKwh
Itmjx/wGG7iRcrXHH+VnYThEcNTjkas2UP3OJX2rDbZvoIj9u/ma2QBdkYZ3ggqU4Mp82SNvK/I9
FROsf/0wwlh5+KlZQ2Z2OhkQ6u7sfvFrFsbAPcXa7Unw6kWV/2rxSXCV5F3OebMVbmxyrUThMeYP
7UPW1UVD+WjFPCKe0F617qLD3MgHzYvZeEZTnQavq/sv7yEmKb18HU0ZGwOC8uaJgZ4SB8HJYDzD
nl9PkNwwTTDOyo2+WkJA3YLPmsseVzMED05/7z04tmn8kI2tarXNRr5vHbZUqmV40T22PpbTDxN5
wdi1ZC8ahzzajkjvkGYcaz6C1qIFB5lHMod3TGSHqkAoI6rtK646nmTLfcaSyIx+2GMPTULQuEfZ
V1CRAfRapFSDqXEkkbePrA5wnEp8/PDTS0mMmN3AOgusIrVNFdH0c5aXQzgztXiOxEul97CXZ8PS
LhWibg0EjDtx7LD0zQ8xtS8BAnaOwJoX2cZvvIWMVLbeCMEmHxFFrdZe2Iy+ujbDII4P/RNNw46w
MJH/QvAEz4clkkUA1C4uSA5OoUcNZI5m7sm9DhM9VAOro1RTOAEQzBAfF2OINW/CUIkcRvsdA78v
JaH0cz2d/lZhWYOgH7ptg3RJGADRAvwnH1Vdl/UGTEryqrpR2R/VyZ0BaxT9fDVbSA0MvtWO99/S
1LqTCttH31lJE3ke1gEjGLWwlwgu0eyxT4EmxwcBLLlt1y4NXl3UQsGw2Xby7FOQtSvgPgkK5QGA
NoHp61RwtpBI83WCLOAIvXSnzPBqaUpzXYg9G04pFibnnWisDju7ZReIazz0A5FHa4G9mbJC7Woy
GAff2MPCkx4aU1cHRZte1Fin2Pe7SfwNSsY8bwE6ftq9TK4e20mWS0ezhC75KEvutaIAkJ4hhj9A
nYf1+fXWulHZ3VhloRnCwpoPb0envNfBtEe35P5/Bf7Td0MvTEOeBHl54QnHf4LVnBnv9ZvqgH/D
40FyBW87TEud3eDgNB5gFKtpXy7m+47yU7G9xUA3Q4MTZw6JQlIdFehv0y7mthPaXEf4CLZ/indz
8xbAC8a4Xq1KZiFU6buXzTasC45htQEzZvjK9ZJ6rJwmkCp6VwvMByzpSLjSN1kUziRZ85tCGBZS
uXmF8fir3+XWgX/M/HZa+xNB9L4QoBWRdEwE+JXpGOnnJBJFC898qntZtOVhyl2FZFAOTEkFDVv7
+uwLwmM4dFn0uE2o+wvVN/aQPYxwXTEdfDhVTM6RBNWJTXa0gD/KcvxVLzV3ca/zIgyE3Z6RcHpY
3zTDrZR8MNblhz+wfPdD+PSA0ZyPPw1YqBgRCEwgPZ9u6eeu2qXA+JeflJCItz3MJQpaYGoR2Tfe
+7O9IAbjMzQoyO/1g4ibP03LWYQYd+0aJ128m7Oq52SFy6JM4TSASmCBvySnAAu4lAGOflAbFe9t
pFkg9uKsgEwOPPPhUbH2doSXjAjHQ8M8dEfPFCnrwtYTzJgqG32HnDYU7QKyta5w7wY9yVeAR993
ekG3ZiE72/3CDJRRAxmY4o+2haWQKUe+QcAMbxCJTg+yb33p+E0Pzzqyj8t4j8md5JinrPoC0NZF
9fBLIYOZcc+N/tvv3a84nMqtce+Q8aeWZool468tPb54JUPJ/tqWQzipk5l7UKE/aTQgQWW4jALl
3PLJo4BunN4P+kBw65IeEsKzWO3BOZX+KZMgsiZ7mWPW8cETbKoVGSThddXaotGMJM656nIVN4Kr
R7Jm8XiUbRfricTDBtpMTVznm/aW6YBWy3jPs0EG9Fu2+yvWuRmBig4cje5UyTZyJJSzOYcfqwRO
dUpOiTqYlrLrE4TxspwcXmzzV9LxqaRTXKSseiwgt/cBLTrmreLKorz34bq4YVGKLql7RxDa22OZ
2wIHW4Op7bEW036eSX9RZFTVPjbAwUmcJu0IX58xREw6oyw6s3gO5cv2KLhVus7XisFAYdlqb26z
bur5hYsHsRf1WsQLx5G+78FNdHlzlgbaoSntb4/oojcAoRw+H3z5AGRD1QnndsFbtd2Kchx+wm3Q
j4096UlWqYpAuQNPGJlPNgEymR3IaOlZMgDJ4LYTyNa5/N5xX8yh51KXF4hJlE1mA3SLoYKbFUQ4
K3yIkLYQjF1+5Jv88qbg/NOTDTyMSUexb2VDSZ9xMS7nV1oIItAaAodxF6lb4zgGE1olckvP5/Nw
tjse4on1XNnqKlR/gkQv33Eidc9IXhHSpx4GaFHhnWBetHZM7wj4F47YFEblAAy2MqhtivH83eXT
gTWVOQQAo4mdzeHVtmJvdMh0m8eHF/5Dje7JRq2YaXMn9sf85gKn5W71JrSMTDrCV2DQhvEx0CAe
yAsKcnowVFchK1bzt/JINIjSraX+rsB2tDGqJMjjlnnRzdldgsY2Y468pWEBxI5xgfWKPxxkMNg7
H5r7BHaw3GbKdXbOqoQU5qff+ssGxJxT0/0ADtIIyHyeRxO0BlrZWvalFl9MSpH4RYqMUz0U766s
7EoAPWNQwO34wj3EnchoDUIcpuK6kThsMQM+LfN1ub7PYnKTqSt06lbIUbORCcCJrsEdnU1eXjcx
4JzSf2zRC2BHIQkmd4LVt7j+kGDKfX6KyhBqvOdZbCQuV/fMpwv9aqak5JoUMLkHQXk1J+LSTLAe
ZNrYQ4+AcEH2eEY4q1zC0aklRJp8w3SHDeRg0m80DXnsxVnJZqgYpwisEOd0zyMrBF374R7ZQNT5
QdI38ljcpklPSSS1UIgNNRuBbWJaA9UYx5hj+wtvWLQyH2qeJJWcqvWxwphPDsiVPtobWOL1IDIL
vb6mnQMVGUmxBfWIXN/mcbG3AWLYMUe6+J2EItDWKZMfoejFaXe1f+MdTC0IqtLJGsg0GpRa8noK
YQ8wYcq0c7XJGHIaxMb92QoOdsa19UsN1gAdBywtV59q2cU9iNJiihqnborj2w/TsZizfBmO+EbW
a10exkLenjsCZtKSp85+q1SsnXeR7V1zyAULRcuBL0Xq6nS2JCOVGMY3g5PXz1un9JU3H9BgFlr8
OQfLludmdyv9S5JtosZAAeKh13LwHLxZ1i3tC8xBrMWhxkJT+MucO+B432no7c9CuCEoZ0Qj/g6P
87LXrCKAJYbWmE3BXK3/XFN6z+hEguek3sSo65BMXn5fC+xkboiWw7qNMRVHU+Oi7/ZGxJ/PwEmt
yLobdh7S1BK7E75GAHzHjLytMQ9UmEWs+klLXLed4qQp4lF0PWn52/CdPxH1TfoFYDzOMiBznRXX
kKdC/zS1D2ocvuIoqMEJKbwkUi7kKtYfLWEMcsqsIp2kRNK6RshrRu4S5/GqlagN4HHbkYDNtS/h
wGucoDaurpgzAa4z8n2HoLSxdT1npyzy50UJNdox2e16kyLHDnDLI/lAdZCI9M2hZ5DSE24G6sk1
6JG2WOJdp1xTn8sRFjHKL4cNq+qN3jv5kpUWJwj0eDl802VfQNaZDkPS+4V209TCr1kUD2rgC7hu
0h+YC9mxTSIwn7ZIEofW7vG+aJ6FC8vMEid3mx/HtV2ytsgD7hF769oHKDPD0OM45GyQyns+p08L
SxGMxy/0sx5kEKmTVCQLkGoHZ3ddgMasGY/JqPhrx/DF4DW4W3TIq1zbMlwYSKhvnjSS7+ubvBVo
EM6sD2/ITlARkOU+oUzM34IXKFB2wB/M5ZqTUKOhZBW8Ao2s6TbRWaR/efIEIgYng3HGuYnFz9Ph
8AXUA7fj2TwKAShX4Jph6VF1z7eOjIqsmIqBuQawcl5GD/tqQl16GbtYXla+L9Z2YibZ1K+UDUJN
y6WMuQJiK18R8SPJyM8T4gaCc7ucrQEK/yMbk3xLCvo0SI2m91ZHv4NnORx/uxIfyM8bWhWo0OS+
JiKwWGslpGK38SqVLttFiS7dcMo9ZJnf7eyYucWpJwT/1VadkoxTAds09V0bJPmrW/fvR7CRv8K/
aQo3LLl1KQjlGtk0rma9lE62/xFMHDkVTr2TSAR8JYzXkfYtaeel36uGFMNA5SV71X5wHmnr8FbE
BEfhNx5wWOX1mStr+khZyDii4L8401VMHSXVWhLmN0jT98pBCHr79l6zmNqZ4KQ42JVvZT8IPd2P
IGgsvgmRlZMPVpefCPkKbnDYTmBDvMlvxSoOD5Mvosg+QZghAU8cg//r2IGT5AHliId0R+z3pyGq
o1tCqrrSkrXY981ZM76UB8qCPhL3Vfl4EHg86hhyCHqqTxdmdBQ+8MKt1/kmTSfPBrausE6kWtQV
UPsdIIMPVh8AET8cV8An7HWzldU98vb2i2SnpZnWvTKPBMXakGrMxeQ3ShhlB2GvKB1p9j9IwzRA
leS5aRjjIOhcq6fOLnX7hzp2w1oYcA94WDJMc9/SWnUMN0lHLLh++UUXOsduIKr2IELQrUvvLNqt
qz5qjHKcBt5JwPZyFZL+hinRVUiRSVCXZuT+YahW1owtAGjxMvNNlSX23ua1XPML4HRfGjU2AEXe
wTbv0hbePRsB5UtPTG/a3DMGqfiEqQHR2OHjYx1YCkBwysQ7CPsaZ4iPI0Zg05EZOrarkxc8T6Uh
wqAQ9plnt7GBWZCwnPaKnY/pqQwnsyvqb+oUT5YJiV/QlvjUUA7tvUzNhv6ZzSIUL/HrJsMkc/KA
3UUVkbPmTlgqoyPIm8ZNECeVtoodrkgJeXOqxDNqFrPgIp09WtaJo1+ZekFkphJ/uvAjITmiNuKU
P2Hl9WEfd4438jG/HWZuJGxpbKnqWK+X6kXZPLILYypNdgH7PQ9hMjzWdMf0hW9/xGLr03hR5D5R
RVuCqVfkfl7Z7gZQyoX40SvbJI76cQwjH/awwIxRRFlcFG8hWmSUm7LA3y2OlDZcxqMYCxZ6Kxv+
SQLPQLZg5t+SHgXBCq11E4LAUz302N7Xmz+aO1wqjLPKtSP89q8M7J2JeGnGiT6qk95uRtecTgnw
whcbnV+MVROkJphpnPrxKrBUfiImOfK//2Yh78G/WsiPkLRhKCpeTx5m+mXToYxcda42BuPgWDdH
rF7ZzLhHb1Wddnh4wQ0hqvkBzmID00UUz/8jNSNPUytXY0EzgMSkHr1rjPdn+L/nD31OxCCylAnk
n/MhVlef5Mxfky4R6HtyL8mif3E+yMzs85pxPC6KOUXSGQrfufc8PjHiOWBugrK3LmOALPRk2fIa
834dziNXm8NOcyq++ImyuUwC2LHKe1G16xPzQdO4R2IiTAEsdpAsW+JLPxvwNmoK8jb2eVGTkSCZ
tx0rO4pwJFKtqrYqCJLhA7oBG6kHBOINyf5XiHipqiycsl8MrsJCkaE4paZZqoUSXzec49htco63
KCnShalVEE2WVt9aOb3XLBmgaDYKNkzorNbqX25B49IGS4NiRn/j/EHuAWzHcYd4du1IuL/y/VqA
UIP9jgHn0hia5urli99SvpuQ61qXrg7O8J/61BFRB05DwZaWwqn2fsNS9Dg0F3COnfjwGOXOgneO
y75ngf+9shgWpVhMc1jefVpazi+xOj7APXBUvywgnHj795tThBT+ELcn2F+Nh6ersvwxujtLtl4T
lfrsbFGSApi7vkEwyhFTNpKnSewWfuuwYgaDiBFjV8CqF/Vt19aRVrxowytjxLkVYVLrqGLn3EDQ
jjN9M7/zgeHVL3PUOtnzo3DzKzKNv0tSMyczYOfXcqWIXrLQ+s5ld1J/HbsnkgWY9QB9gJgY7jUH
EbMTLhLeC1BrnRPqtvZ+WMbxrfGN9t6hLUs+D2HvwyVAdanTAwP/SdsHppJyslKSmzKBFz67z4Ey
b8PAtplMlWZsPkPSx05HgnhCBdl4840jTqRqhNjHJe6a9WSVx+CiRm66vPgRc/1ZwMqIwVqziMqR
KxT0viVlIWa7zNjnrEQgxdKy304F0ZTHLBAKIZxK6Y6/BBiv8DvLdfsRjn5yWn7Yt0yRf/A9Tmt0
IUJ/8xkEghWH5OHGN5SAvuzI8ktlg3z56LkDhQctKvPq1+kavwylG7juMPKF9jO8obDHj13ui6Kw
dEIG6j8I7/iTsfLEsI0oq8V/NTESg/wiZ1DCydK285hU1ulj9NXbREqJousaQyWCo2eSVCxsqvsi
cnAHrfeNpjfonQigIAKZ3X8+/zZk4EFFM1tL0n9PwUNR+sIDFFo3v46jYxe5bPrVNWPJHrrtLKbL
2OQdFC0tj/Cy9cBJ7UrlwamhiRk01Jg59IQNYd66QjEFINsZJTkQB2OEkfAt3rHe7EtcuA8fUZwl
SJjrtcfD3ys63CcyEwF99UiTikykOlahcwXgq0T2I+7dpmn3GVC6pN61GLDdp/AU3brqRc/XLAaM
rsRhQNJkMFXJP8s2aVrEDSSorZtTfEx4Vh0jlZAi6kM0CCDJwo2+ksAAeN8bam4E7btyG5Y0g3O9
RL7GfHHaVelDe/iBZwo+v9IyUtCOG2SEWgs3YhrvLmZOHcsOB2nC4KsOtW7Jp4m8Db7JDD3pJ5sQ
+Nm4kaafutUOvCEqSrOZZPIhp05P6VtYLFnSFiEyJrqn1DIO4U/Z/5bBJGZe+Syz6RTiXs7tGWYk
sRYtkvn5Ja4SL6sbud66ag3lEWR16H6NIweyNFBZ/9tKvbRTiCbvuRNpTyEJBzST5dP89xyPUF3o
cGHTyNalZlRoDvuM7c76DRGRgGmFf+WCViV6Rim5I3gVsHhCPE4UiIR6SM/7qsEJHkXzsl6faNwX
TJM2KJo3S4x8DtbieWuEpZ93YsRfUFeHPGU8S2RhsZZ1AmfiRCjZgoQ/oChd71dUBQKjV14oUTam
XfivL3hFJnBeaUs/2bt2uTiZAFUAw2L4FNtX66wKc48Jzfgfwyv5VPoeZtO3mrcKfjsAuTJw+k5G
FTH5RQUYO5QZItz/tu0xGXUJ23QoYs5elc4mr+8pxPM7NJgQQUsiun7ynCTDKgp974Ra33VclovO
GcB90ndhTGwWepdcGHBA2w5Et5fcGsbNF9nzz+D704pzicftjoC6xU7iqfQIv7wZ/BmU+blz84Ks
zKgPA91iiuXZUNArwS2oQZ0vQo11SWsFZ2a2LbAgwMX8QvaWSw0jTJ6705BHHbznt2kJ1A/tURSt
Q05Jn299QsN2hLikIEV8agawmOhHSbXq2lZZDdrva5BmPZab1edoe3fm0OnOLI4Aq2B6vdzlbhtX
xKMjU111BQhe+BKw5sC/pQBPSTFa2Sus8j03/CZ0dDI3wUIxTJ5T8smk8u6J1ME+Nhh4eeoDUlPn
AKrgBa/VCBu/RPqtsGP5e8M7tck/PoiUbImbjMoMAjuzPaxnSBVfPxdYiuCE4YfxMCLPRNyIsSQ+
XyJuqcWma2meNJGzBoLeVLPCrSiJksDeSNpztU++G8/ZyZNuelZ+msmaJFUnXebI9GzRlfzu8U4O
Yd8Z1p6abi8spkq/quboCPD1C2Qe2xJh9eEwEIeb/p3HrAPLZo08mGdsnIbX6tjMnSYla54YrOwY
+fKAI5qn04cMC3cC5qJRXMnoSZtgOe0TfdT2/exuBN7GiUoR2sNoWDydneLTKK+eNGvCWALVr5d4
eR9I2u1F0gpGq/CQ7Uk9zhpRMt0wXtvnnFdMtc8mLdiY/RZstfVjzsmU+dRkw+ypGwZuem/XPkB5
EaAVfk9uWjkQHQoDofbRKfDritCxVgGSIWiZ+i1Y1SuFob6ZMGFMiM0+mR3z6unM3q+xThGjk0Z1
3dIM5B/vWmHuSCmDttt35wwgyvUbUMYu9u7BRTGM/AG/Tnrh3oQH1sAJPU1dfMRnP5lsDB7oJvbs
/+L2lGO/xN8MgVk6Rm4Lka2Iton36c7NZoJP5CeZsHKQU/xKqF0R0uXOic71fLZUIi7Y9+TZBhw3
3szyemKfMtXWfaFnG8oGjL+HcLVXtB+dkIZMz4qtja2vjXU4lu03z+Eqmhi/WMQ/z0KJBbBmw2Ok
G/WtE57yYgypKlxAGF+9bbUCQzCNqMLym/IgqRM2UcwJkoxsin8IQOrBMgmRFJGDhu6H7VeazZXx
iJt1/hMIsAyhWUyojlw00VGCKpYe0d003+laP3CP4OlyNv2W2Uem4LPShVQ251U/ptyx7W7QPK7g
hDaUvAsmQKqiAx8AqO/rlJ23yR9evxDiw4xsT2hAcTV7YWkMVMwpGuXXvZ+xiUA90J1a1qYjGo4X
YOIYIOXIhgc6zJ+5aYf4CJ+ycsr5UIes2QzBzCFdCNIgiZzgtHhcUt9lC/3DBu14UKxreM7617uE
fvG7xjJUMafl7o5Ii49DjRMbY35Rl8zs8qh5mdDbid9ingc/hlcoBXrpsF1xULggb8c2iWNEcrOi
KC2M21J3q4B7proctJGxn9UHE3ZiXfjf6BtVjlFng4xG0anmw6lTv9bZkRCkEMVxmjmQvUUqOqXY
JjGNNNguUlpDfPWwZcxJpBcJM3soudfYRdSZK5zJhHbZ8YPiaK9pTA7PY475wM3vkFPCQddpF8rK
qP5ev7EFiHRiV4qq9ZetDPn/3I0hyNTRu+DL4Wv/IEed+bd6T66gZarJ/QY97egJRDSDJIQbvTdv
p15Ptk/Y5F1NhONVy5bnb0618o2rslLsYsXgIuAS8zYBUsgUkiJ1ET37DGfiNKuEf5DIvk0amMSA
nFj9etnaUcXTwpE9c+PE+10cGEKTIZfug7YEbtYRDSfJ702lVNztobYg/7Y3jirb1DuNZaLnVx4g
c9CJ1qqCKR+9eYn2wAbrO5bRNq5VCTayx9tkhO/FDXADrlin/fkMRbCKpCVidyfffIEIPVoP6nut
FfY0StTln037ABsy7Xy4898nk+iD393sFvIGMfMdMJl61eA4NEOAh8Bq1bo4D2M7rKsWpJKdB0eQ
2Hm8UYhK/9htVS6PYebes4enL0jU83A3amhBjTu8N3pbhMO4oFBfaOKUaiZCqHzP8zUBZnhDOv7R
w6E2PC/ypVkyB/0JGTCeNjlr90cTI7fq+5w0hDLBFEkWsDIslZnz71CxAO2mVn62Mzs+BL7SvH2P
UZAZH1aZnlBjLMCyXbnEEXI6Argr9Nke798CNfZI7q3hG6Pca3IsdLvGWFcwD4Ykh//4OKyQXKGa
6lUKMxgg8QdU4qLMrv2LyjNM4VbhT1Htxpg2jXc4TTDVXMYLPxm9evNGOkI8t8Zk54rjiiOmpU/M
HYjYYymtDKhqbliL/7eNhQ6kGNAinIf7mW/JgqX0chmTHCDFLZaHPChcC2gIrH6iJ6sxAcu7hbyf
KouENIZg6+beu13LaGiseOYBFJ9TRce5V369/LeQoBAfhfzVx4INEyAUvvE+tN3FsAPHZ1c4Gg6u
/g/0IUQrt1RAmcvv5gotnVILdvau9eVEtGN4k3HfWGAdWop2aOSotzAxUu6kJiNm1X2tRdqRmY8W
OFIL9WY4utu6fzkBGx9QWBIJI4LHX3nvQQGfl0kaqWWVcZnGc9FGa5AO+fHY2fk/SxoIkPMtUBbF
fVUsMmmpi8rWtS6itF/3lHK6BOtyFmjfmGpfUxJhpQUDIPIQST8B7VsVQ5gR1Qckqu8s6BfczY9Z
lOr/54//aWyiahBFyJazvI7F88ys0cjo1PeqsVxaJPXc6accq/W+nxvD2jWT29iLAO+P6VVGtwuU
TV49L8mnRjDAyfZsLCAcS++lmLXsxmjO/O+zxiL3qkJ3mh4RK7C0dIZKqfMnXCuwu15gErV8WdNm
AATNs5VFfocjeKlf9UXPNQxcMJYxa0WlgDNr45P+R5gHQDpVvGhfy2aOQONy8G5sOuEG1sJD6z7S
62iAfoJNGIMOhDt8YBTApi5MrxQufDwLDVZPBtDWDD/UPQE4hARE97CbruoWD4q/nziWA0iW+axe
Besvoar5ERrkcOf07WoushICTDpaRyvj9OqvWCdPOO11qN3TDfHxifvNy6upP8TA2h0mPWyBivvV
NaktFJnrxdtLdH15gwLDvDMNcgpjXB3C4EWxK2nnrkM3fYS84B58UcLi4IXkR4G36rQ58CQcIE2K
pqVEsDu2OwBjz2941PqkdveHRevAHeqPuCC4n++sEBYNjFRqokE1mi7dvp6H5TT8j7z6Rjxva3VP
VOzbXcUgwx/3kEHMOI+FXWnveUrXWn44uOEEus59BwyBVvfW1n58lLlgsz3Q+VAAmMUqo3n41ZAd
JQmFddt+ddgqVtNAmPhFW9WPmHqzNl2d7Gfasfv0a5yb89HzBvmH3+PXm7G1nG1L9KBXqLiJ8/G1
MeaQYOkTrxrnrvwnlPlQUkgVjMxqxbeK5LGmfCx07rOyvXHCi8GPbEh0UHpqu7//qHxMYscHd+WL
skLRBQaTgv09Q40NneVz7sI6C7X2EUq7IOtbMVZuLZ5ATm66pe82EVJ5YfglXhkQ80ci+XDGQ4em
1Ae/+pl7YioUd5UmtO9Tvdt6aiDPrPGJqZ/UAtbg+Kx63dggiILLgrhM8EuHVP/RFZOaGUkOdeG4
+1mKOprAEFdhz524RmVSQW+aQ10RwO2OOMNwYto/JkFDevkH663N+5FX/Q6mA4/nUTsZAR+uYCEX
pR6i+jZGXSOdZ9RQZjF/248CYkrnlkTBpXZ63ND2EDZIYvljOjJAddLw+/AYAA1xe7yJ+FRVjHLE
FP9R/NIJOWtkiCakEXhK7RUgVrREZ5OCAR8boUierTONKUFuMkCtEVvhvSq1d0mlH0TrRxXjr9Sr
68GXwb+aGiVSstemLJq1SipP42RCAT9FdtF0w56DtdOK7xfW9nD6ulc2ti9anGU0kMUw2ImqL9gj
mLRW/1KEz2Mkm0XhNI7sGW2EaBLggj1QjtemJq+g6mKpv/ENRgAK7GhDBfWshqTX2XabUWrtIKNS
58ppeDDn579SsLl0HyUsIqK/E1TUH3k6lYsU3wTsZ8vr7A5tK0Kef+Jm60rA77hEU/NlPgyCsfCK
5BvyypsytcmYdNkvKMpr1hQ1muiYrhybTEm942e/K2psw0K4kMdfRpRlv20iQRlvq/Xk9Zq3+wFU
AU/c+Knfr7yzl1cr7g+gzc7ZJrTAGQHvW0e5d0Nq9dYv0sw3WjnTfEkur6T2L7wvlUxa2jyrTQGF
lBF30tiR1HnGCAKYzCMMBWX7LebG+84/P9WU9j9TU3RW2m55QapRxc4XmDWkmA/kf0oltSLO4wTK
v7DXhkw5djDaBcdNiBa0nzj9ojiB7F1c3bpHCrdkkkJgf6YBxno0FN1TBtN++8sssH4/QujECITr
xIG47xxYxLcbDwE7AoZsUH3O3LqetzuBEk/GUhwY+JtDQr5p4lHAHYUWRgaYCCNRFJJMb6d0jtf4
vd6k2gIBRqomSatNvR2QvA/JQGcD2PgPVL0S3N2Km1tfLH/+o9uuGDRyNU25Ri61bkZkucFtjbxC
8stMaMlRZmYuJg18Uy8oG0yoQb8uqXAPkQQZ0pOX8weBE76SwSe88Sz9LXt5EqtUKw/IuFfx5E6k
OLGs3OJa1V0rsajrM3QqzMq3/PXoN9TKWRBAhLzk0/GeS+T1dsXLGxMS2kHawVec+j4U2QKL/I2v
LmM00tA8/EG+wwDPd7RP7sLbRCtUGnaDWZ9PAKE5dX7IJC4r9H8m/G3GyvdWBtrrP581MGsMHeaZ
A8tUBuo2p5XfV2fLOucUt+gNpP2mTLtHXxJtiTi0h2yYW7dr+0yy/RnSjeMXp4h5PFY6n+Rrfyrb
7FjJWEYHKuwCPvaRsv58u9ZVMqFgjMJeY0IEfVV235MDvOKYO9DskGX14Bh7HeZVuu2ebwNWNOjd
0GUAFqxwcEWerlPHTA7vCpQcRy4Cc4TAHo+AEdd1H+ji1RHHD2JUzNWKOHv1RqJtolSRGLxdwuL4
JKxXAJoA77jTEdNPKxHUByjrfNsq5Tc6wl8clGCDv87RBGk6PU0i8LxThpiWXd5+4HA4wKggfqCt
ha6n/uSkQ2R/PoICgiXZBjbUzFmaFlKDehw63ALFoM7LynMGmUZBZIt+eugXk5G+c3CBxu7ajtGy
bckkydL5XS/nIdLL+Fuk1QErwXStjKYb4bsoxHH4Gf49rw633s/GxE1YrpsrBdmp39xRkIsb1pt2
toNrb9TGxbcT3l+FeeG30LL0UbauzhYbPF58lYxUE3sC7CVjUDLs9qKNqfrcbW9JK6qZQR1n8Nll
+7sjaXAKlozW6EPOQOrJ6wB2cf1KrTP6x53P21RRcFjgOX4Zvu0/vToRBx4xUUJ6jGIa+UZQmqqb
NuU+oYUcKHRnNyLHG32OTlr+x4prWz1AUTQ05iKC8SohLbE6l+F1W5lzfnR3ME7QzeUzbTag/I5r
U/coWSj+P6K+z35wezYcZDtf85NJjCiNhVkxPwju9NzYHs9eSxe2ZNkL31rzH8oHhIkA6ZDcNuGd
EvoTzqNgy2l6h3OYP07d2UOJQsALi8oIka0TZ8roI1OeTDMpZb4YE/oP+zKAIsoPj9J2BUsnQc1x
wAZQuxYOkqTtm+dKBHy0aI3v4mYD5pUxV91bmegleOwlrSVthmFpdhbkbAxHxubT62RhOjp/G5Cq
O/alwCe7ROChTuHPXUEIZDeZKV7iFXn6Z7vq92C2QZFOulPDVQgcVoWsgXzogt1YYldeAx3BAmdh
8x6C+5dRERenY0vStQksL3DJbyCZEmc0y6bGr/Mmee2Qpk5fTGxThggAAm52jb9F2Dy4WOBGDYtL
qoy0Ts0BnH4XZKhkC5jdZZOFlI+e6FNQyNE5/DMoIackwKd6U3ON+ql0eHJpoGjhHgX6ixixJkl0
/s67KkgeXhdqMmzY1RVegHQdLIqcvaDbsXogI3aVUnabeHGFmL3XfhDaerwOa3KBfK4SQIV+9/oF
JTn5fdw2Bs+J6fVF8dWZ4lJuOTANy2QUL4KPMW00J4p8lokWwgbOa87iz+IJnybbX/mdyoGWw0Jj
/UguXC1C/6Y4wMSiQ11R/8uAhGdCWhWauK9N7d4UKr5UQ8JCMfL9BMOLMQyKzeDozeSgSxE48QfM
5rwCXGryTr9LeLncCVCgr3P+nNf7Zh5X4GOydPqJfq9VlzvEXK2BckrvG+7GHp4OBstEYcSzDfsy
zYp2odyz9rLs/UWSZuSnxhExXyNoy6XWcTdD7HwWaAham1hPG5if1N6yRA6ITVR1sDl7FQGeE3UR
WytMm13SmzthPmnfwNDf3xDhk1VH1jSOhqRmGiijTwFShk00swwzc/kiD23G8Ic5sMqoKjgIMP8J
pvscggQd8plY9rUSJyvS2hIE7C7PHCwzGHfeJRHpVgqpfxoNfnJV7gbCUUnVdh4D+2hzIY08CQMb
BkG6nq6U8EiSGA6k54dsoJGaadxceAWXZZ8DZzFLQTUsiG4ZEymPrO1dis7TmTP1cRCEkm9zenfN
EzEsASw4A3XZt3sfO1lpyf0QwPfU3k7Qzv7cthgnB0P0CCOca/U2cSGqlqDQn8O4AMVf4gWdk8F1
4CHy9i8r7ksTbou3XQoejJZNNCmfAIBhdlkB6cTyHZxwlAeNJIgoN0yNSKqRRo8jSDBH3yb+lhqS
lscijauOOs75LvlH2n09GmZEqu0IYpFE9XcDgzCPTMTmjxLqv/zJ+ewBhEGNLFrTHBv/FeaqaLV6
Cvg87jCDPTNRcuYIp4o/7xH6lUEZQUveXIQEn6WYglzKObdr+eYE2E7lneTiNTjfHPHfdFM7V5KT
DDdBb3ev8oX12M5R8oD2f3EzP6stUWL1TWEH2r04Y4WmZKTBOIIgcnGCKCXglmBz68kOr2uAqrK2
LobuSrHm0q+Ijf0ihDadXCaX/pZbtpMpi3uyDeN7RhMOhjWsIvQ73pYRREtftAFf7wZp56L8E0Wb
Tju4TKVo0kIdeeVEoCSvu4hutbF/HKR5nKlRNSAsTRH5zJrP6eCZKu+XfURhuMRQr/4+lHfu2z9p
81kEM3dH2veXQ913ytGUqi46AXFBurhsUnJIEh3zp/hrmNnigLidTg+gdkej48UZNQ30r9QKRdRe
dSskMyzahr0LAQdzUYAxr2Jqf1iblBKWJEYul+SQ35f7tnSy3jQKCig3c3LN8nG/31YwpTpsnbnS
HdoB2N/zxH69op79a3+BQ94BjTurXEu5IUv0iJtIYVbELurNxiwo+1QxPWG2WwcxtBnkaBFAtkGz
gO/e+b9Icyoux58Kuz9MoIwfQcQF+mpiBnjBu8BfkV/0JvORotdzyJdhd343YuslF5eEULP/JYCm
TFqo+E1QIHawOHFeXA7+G7QC7aYx3EwEBRenvTi9S5l9OtewC1uvMzA0EWAJrcUeQqTxJ4lOmZzl
nnCHvEcbfY1TsIQOsHS9tfOObsWHQGVYGgFuP3KHjnk9NZDi5GZUI+WwXYUvTjGQCdElsHTi/0aU
4wtPVyWVl3hkaYxw5a7UeHn+4G1wgIXVgFWBUl8TKmpDqvb8+bwAFOXbbs0P63lq9S1OwMPUK0lb
GcgLEG2Scgyp8d1FM/Lefhnjr4fB2m46AKLLVpVF3qqLVrDEVdaSUwUh9PiwG5eaMO26BusH63CC
P7ix9eNg8wdczBVB7cDRP9VGgBLnTRmhtrLTqo/31s7AubVyyGsZk4v5h3ykn61I8JMdFKmRq/DF
nIoJcYQ0+ZGgyBEHaOAy63E83pxfuXkH140rgnQVVo6l8amwM+d8VgTGCkA7Ce89dRB5xpBvZ5PL
025ft5g/v5eKWeqh4Ur5W25FYgKfXm2Zqk/xgkOXzWZwlDN1WzJRZr50TzxGn00JMt2R120SbHzj
aYt6uH3HvQBoe2+E54BGe+nSQzvRuWhECMb/TXIY88Zt1go58WdE8y+ncoNNGQCGdNSMN9pvNsca
CCeeUVwI8T7n0AQlfg6EgV5NyLQ985qUoAhST7jTiZr2hKMZin4NKtDkXxmzwLKj9LQ7JrhXDP3x
PiYRskYO91a0EU7CfQCa6ozUZcBEpIXt4jqb1xEWGcSYkgjjljJvF0XtzlrFjbHx54txtFkDMR/1
48821k6vGksZ/lqinZaOB2GIWSxbvj1/QIqXeHFDrQDm397WmMbMM64A0FZq3Zwznme35gyOjv+2
+Iq6sRTmKR+5XzwWeieOG0AlOe0ZlLpF1Yg5vOfYvjUW3ot5I9ZPNyxwn10IUag0pXl1qZ+iJbcm
kK8eIe7dFvGL32SEoVAfNyirjaDo5/WevFUEevzBNYxQQrfpRzXDnKLI1yIr+BAfiWi0xB6CJ/er
NlgC1bYHIJkQoX+cFjTvbPXk8v3W2rlIbTBVRp91qV+S0DWbpkWEzAk4x4ghxTUNS4T2K98r+ZjD
F7m/uc46u925OPkguEgkQNuf20RfZa/Xzt4Wg7WPwad1xsI7VEPeMNAaSFRfolXeSKukG5G0Xugs
FiJjiaRJ0kmp+y7cwD4cgHjUwFWdLLzYcaIXPqxv7VUadAiq0ENLzwcqreEd6JGUzf5ukDl/Fo6/
QdO0t+RyCyy1sEaE1pltWtuhhFBAKoLkMKiStyL1kGCwp0QGpCcgDk5XVKOir8RolKfch9VimIM5
xCWSAxJnXQGrl0meo/+2DWho5oqp49zrL5fU2/BFfYU1knELRZFayD9x4Jl+Kv47oylyPj6nxuK6
2pa2vvHGzcyArt4OpXtaSqWYqexrjuVMGaiLNpihxwDt3c5ui0x0ynVSX/FrLZjQeTl4QNVXbHvq
svBvFbeHlaAu0byydkXkqSEHMyp4Jqba1934SI9MEvFnxLvorMG6/xDNruwlgBLT2wRwRggeETyK
sQvx9UGddE8ntyImmccGcvZ3x5ygDHYBOj+iQy8MJkkJoB+PFnO7jDcyimPxLqh0npbHkjHDrprG
GzLTj9DVxMekIR1khKVH5si0nhZKNq9O9tS8TaXWDoszCeVKEFCbWxP6lEXW5gyIk8aEMg2JTVJL
uhVZZtc60ptUFtPnrZNCTuAMGWTQFgkLnSr/JQt0FhhvG2zEZZ9gvOK8wXS0PpLLXgoxaDuXvbl2
1pkc1qnFaI5TQOGhHSB9xdOdvw0JTj7DM/Nhuw4zfP+yWhjeqE2hKYFOGAuSY80Hqzhtv+BFVn0S
pmcckeHaLGxCxmV4G4KSkrE+RfqjLPX5FFaFG4MEVgADFCleAQgHZ0gdZ7g4lj+vMpPHcHeRDNRu
p+45/K/U2rsf1u+A2GLIaa4udvJ1rugcWPqYfg1iOPLmPNtc1yCpf2sxomH8lju9QpMeyJxwULI/
0hfBFY1U7R5R3qk9xopiSYo/BOnQsAMFDjNPllEh4ujKmvySrUxuTf//BZB/EByTGeIbXrYxs3dT
l8KlajhLtBGo3tuDBcw8DnYV/TTFuN+mXgI8biaZQb71I9hl800ebGJVK8mfqHqQup2/b+nm7hrp
RtlIbSxtZJg9YAAE6Pp5l6PNBMK5jSo87d3GJAF8RXaesH5EmWFVLL66khinVEf7eAas78oEMKLh
YdqkpD9Qv5QONBgFB5e5VA9GY5zrNKyv7GP25Q0Lc3AKRb2r0M/c1VmX+bR7tPLGgRulbAftzcCo
aItW9yG2wfO+wx2cN2sA2lM7uD3MgMrSH9sXed3+cF644228PHisiDt3ARe7lfBCNT6JpoepNdYa
3nfplG3SXkgH5gD4sbRxbFVafO1TLrw4t1RVXhcdGsN08AFIxEyDIqc6FiEscO9YXEGJUhWyzh2Y
AHrthXP/PIuKS7DMj9Me0TBdnjpB9yIB+zO0mgsBK6xLuPVZ+9g06Pzg3nSTKZ+sM5TFYLaV5Rky
oSaTIh5HdziLcUhVc7lmZHlw/x0+aZXuNf1XzlMmJ/OST+4mrft5vj620GdyZjulEiFE+SuIX/mN
EsB8eHaJxxgs6A1KjWEGgL+MUOxVlNvheV1Tv/LfD6nmlZ+rC7jL9eG/H6YR1iFRvTTC1Bx+V3Yd
3IoQ85wXyvBm+1eSyL6Jlg3ZHoXj7yKF+l177xdFAWBLsctqYttyx4Z96yd/t1E+nhfH6tFJoyH1
rZBv5/NzGohEali1siU19a4FJpgA4ZsReqRmzYQlu0gCnse7D9BFV1HLI4IJbCe+8x0q7/6hpWCk
FOfBwD2WPly2nkO6VcK2s9oxRRyuHTZHnRQ+tQ07Bn+k6LZDLqsgsltyV7SWzMIHB1tf9dxxnD8U
xvvvmiXL4noLUER00CX8WI7dM0Ee1ihwLdmLLNMSCQC7UJ760A3ASDS9I2Ehs7Ijf9eEQqgM/L1J
06tJj6tErdbg1obrcy/6O5Jj6io4AJvj8/PF+1NO2tvqmRrrfgss8sxa3G4mSqZoTClcdQDSh7yq
8ZKwexLlSmcxYglI0iCiqy5RI1+PBVNJhOeIXimBSWc6ZzcGtUnu3IAqhH5IqBp8X8HAyn0mrr14
9Ql8I3Qmm3eo+Mm5Q2GrZGcNV2jxXOoOPm8LcaeC8iMN9TWy5Eo0It9O4yY0TiDyt4j2qkf3i196
N60B4BxbFDLDjzbPTTP6MRQGxMLeSeUG9esS5iKRyyteFtYNtW4vRYC2ox9GGDJ04rRli2GYouda
VRJagHiwiLMjUspPxjpIGSU44ekrbm7YVLJXOLindmNG+knLFrfspKCTychz/U2deyj9UQiruVEs
LArO64GIITxyjvwxVyT1k/XAH55hJgyCGuawhxMHGdQc+Nkn3Tuyfa9wR6R+k8A+yx/oF7Tx41Yk
rLu6uktgenxjaCdMt28MkD6yfZ3LubQy81QEQgK9kUtuivaJZNbOjadV1Wz6jCTAMcSlKuLEGV/G
kBPUSbvEo9zpUQYHctyHX6qGGFG7eEtuIWViol2zOx8lx/mQVtA53W3oqMXgGHwW/yrAVUIbJEG9
tmBuGTZ6QcahvjyZPKKeTKWrXSg5NLju46GSjTvC4HYiudq7j5QGuFUbiSR8P9tyVMGVIGx5k9Dh
QLbJeToFCC/iTIHEAyzU9n9Ehtg8+o6RIZEifJkMenUzDjgndqviqQYKK2jKhHOITb5jbbauG/9N
OIxk90RZUyr+6DAdglhaLQGtFul700FQ+ejAebqmeDT3b/BPHEw1N+qy5wl/Vi7MtxJid+YWUqQo
jBGd3a0/WeJaCxVn7Wub37Fk939xpEGOmGdS1UhtQH2TgEPVAb7o3h9Xg5OEZXGMDb6HgI5A2gSG
cOV5wJzgdtyb1K1fsvxR9NTM0XOeqH+hYaXObwuwiN4G4OuBePLEQiq1qkgdsc4bvUgQub+0gr9F
egzIo0Rv1FJBDVET4xQWCV8Id3CJ4hv+YEOO9u2q1rA6eEb/utjRtc5/O0iiNArke5j2+u9MpX2F
WlmxGC1Q5VVIcel5V9T5bF5Xpu/XoFQeeMd8+OPtwfLgQdgfWQFH7wG/jXE4Gdge7YiMrYleXNk/
Tych2Iz2zOILFvFcgG9e6cYVEYL89SjTKnNKUXPj/yUo/tnxWMJ5fOV6bvDbYQjYR0rQ7RgrWWOU
+BYKhscZrUkUSLyZQhibOd/AhhKykwRGZ43q6sxRpY/h5AAu+yLw9xuRTVqI34o9y2pFppwET8iz
gt3jjDI51iK1P1JDfejVIwlJnukqt9xA2GuqtmFEGAqxC3BojrhRCZJmqXWV+yL0CqU81Uwh60D0
8A73D1qedgNYVJyMTd5aSzaAdhSEJUaegc7h4TfFoO7qnwRjLopg9KmzmQFKpw/DTLxM9GeeczWH
8QaEcPXFV2ND7IRL2uZzv9IXtJnriswX1IfKnNxxj0ek7zn8pF4obv7BZ0t5ldltV/V6YZRV1xkF
FHcHtvhpK0mGK3lJQcj8Q/VjCPxzHzLrkg3DOgNOATqUPBQgZW1ajZnMUKtGb9QgDJ3hfKBqfS34
kMdqf9MscLFgSziZuVDVCzNTNbPkoHumQRLKptU9QMvQjJYBVbBFXjRmJ4edG+Cg2B0iJG1Q9jKd
B2S+D1/xgGgGyJGNrI2cEHLT9wyWAy9x0CKpRS1uO3FbrsAYhLbDzZ/plRipq1xiCROOyJkFTvgk
9XYnGt9A4gmc4S5dxyldybufsjGUgeCCoCo97ksEIjNQ+PuQdOczwLhA4PCTV0SzAvl5r3cIyF9n
RZxIiawx27xPySQnFWmRb4DZL4CyMBs6Hqj9OVMXKfPc/LKhoR9CjEmpHkZhPPoCBuxUIyFiQ9Bt
kZpzsKXIj15YbtA5dC6TMiLrpcanAOAI9s8bJgl6//H5IBdU/t400ahD5GmbMFX8j5A7Z97zqmVH
DZrL+nNuP8AQmH21RBx9kbTXpNyLUrSf7zoUdI+YHGla4Wu0Zv0/RL+wzyERHiIkeUijJMKDi+bQ
cnTiRtAVuCjLnPbOqttg/CvIGG8OhivM4/rnvaTB3M23UeNsEdOg1AHS+cA73IptlKhU0df+4kab
7wEscOBbLtqfgFyy/7fK7Pnjog+xps9hKWbFWE4KWqC/J6VkPW4H8ADnbt5JAwvl68IuWZfZ8zbG
D5zbIal4zizPAYVemhucG+8ZVART3ogtoEQxdeQdEWrube+9UKVqdshMTsxdzxovwomGrre6ws/C
daYvbMN6BwzRIgMMbQN09dgg9QTPGjvQDNjh2lUCeDqbJhYJdqr7K0f9Wq4AnMMNFkAHgWrMELPT
M/Owdq6qDxOyjVk9R/6KXeZLJllS7yFUKZfdo1Be5jQDoNbU0itaXIIEQ5Zp/JXYFhxiPQyQFggo
gABHOXakLvGCjpW06U5wETmKBAhN6leH6M8N7UEOUlOYdYaEHHSW4q9wQC9SsZ7MGnSJ/DAEUtfp
fi0GUGBRMYxrUT/tvHiXCIGDXxhSDeiwa4zu0fBjTDEP3MCquD86npZAiNar+q+LUjNAq74kIP2m
S7c7uvqfAXgKobbE56c06CCC+kMOaaCiEVWXxUjCdw3oNlKvJ34+ex/szYb8zXSpuOe7LYDD1vsg
j0BCfKtSsR9qjcoeVz9aEpMHHapwIU9qEuca82suD8aY5tLPR3ml0Rcc0MaCdIs9uLBFcLc/cu4t
Ja/VN/9LwEzWUnLH9wxAbEXCrGg0hV1zNhlYKR++mlCYa7Pog4+1TaYNss5hZh9XyoFRlmC2YTT7
smi/QzSgqVT1bjgITZbbJqGgwr4WLV7yubGW6BPA5128VEetjcbtWAKzIVMwJow0kTSIxnZ+aynJ
hQQ+GggCI4dWynggCka1P1nTfC+iYaIvVaAcmIpGfTqsipCPQbM1p1utgE/OnZpttK0cHoccX1Gd
hdhz9q4p8ZUsCU9k7jTt1495so1g/lqNUhSnKVyu9M5L9p+qkpjEM/JXN/uoS5iLyEM5B/psiQ1t
n4r8snc89XYQkpniO/MYy4bOzGQtSW6QrrL4PUHKI1h3J8yhfsrBqfDnqoqm85YPl5x923QDny0h
7cOd3qN6IyZzPTuQ6RpFKuBcjKnbSVrcWqy30TGRe5mOqqa0tExx4Q3J/K+7vzACcPVrWjvEcoTT
flTLp3rZJwe0GCoqpmz90cBXyx9+vPoP62RlZfb5vhCLhmxeSAbIjlAGp6L6mgba362PhiJHGq2p
lD381bbuIK0k+oUdKiZJag1U3TUm3EraYGTYu/QND/GSR5YGSzz0J94Wf7pPi/5UmLJtpWoZM0+C
rkMVtTrwgLaN4XwkI9kbuJ6DWqig0I9IFba1JngwDzmGAWBdcQ8fkVHVTjqlMNU8jSx5YW5wOFy/
Gksv8kQgZw5g00ARByt625TkgCF0YyQlKsQh/TyfLa46jVVsuRuN1qehl9ddvLeUDSmirZ32LhvX
W3/PFknEAieVV9NER+iX5AO+sXdu82wVaONM3hx+tTRdIaq5/u64McMEx4b6CCpJ6olT/H9ll4an
lXucgIEK9eAx9KGxQKSJppZD2L+MMUft6X72ZoK/iEUf4f/alYZElbmBoHTgUGmkm1stWPucXkBQ
sQF58jRJ6f8hUaBV2iN4TlxXpMe4KbSJOWr5j+MuvuvqmbxUUpLjRWAkLN3ni+LVZ/LfJQrQe8X8
mrYDWgkwTJ/CN92UMJkpGbxkhNmGfhQwHt46CbdMuRHQNtj+tnYlEUqKtmv8x1Ew1maBsTvrCVFD
ziAHpizygff42Gcl6lS3YDntIvqcq+b/Iq37+/ik+NtPQg8wYoLLcjSnHN/E1HdPlkMsF+DKIjls
TdopqmV682FSfoWRHyhvA+ngFQ6ciyudIgXjh2ED4AW2fXTllwguOF868BLorNsdVH0TRigEfGCJ
hpYjuMJjECBygyEfaFUrnbMYI7CNvoAW8xPpR2dZ6JY5wWwrzqNn99MU8SHTtCE1UlxHVLVeaFwa
4DBwgQ+4e7LbYtMIs/11qzmT+mh9DkXqLkVcDdLIIXItPLqNEyN34ItrTotfCH2jj2fD3ktc4Pgv
017nKGIX7X7h432IhgbeD9Sij7GYI7unl6H4peamDG+YwvFwQ+tMvbu9eXEj5HdOzbvzlpHPv04U
vwdtyJ+S8X6a2xE7W3Qt5JfTQK0EQY9EC4csOFEcD2YDcjFtE3T5ZNEbb5iUUnVEtnPpvFrtqDgz
IFldmGza3zhU2QE2pQ1vPOFKrJ8yQt5QnRdcLBnuJQoxaG+2A1i/2c6Q6xw8YbFQ5YeoIYyExJbX
jF3d+sTQa47qroQSifVjPc6zH+TQYvA5nA7pqCx04BJlZRNoiUgLxP4aJeu2j/j/nY+Z7hEOihoL
FJRnDy3nCqFxAVjQMd9emROi9BxIDe2PuEfc7G+i0MrgTnEy3s+8D48/JY5KpffsnvpuHhr03AJq
prTPvmGluKJL5SMpSS7q9n8I3ET7/xFktegi3WiOzn/DXHNsqzjhzDgot3z42gxOx7Z9dNnaZfnq
7BdnT/L1ZyRIN2wGrNNGIXDVs9EBX9IsKuaRHmqHkj634XbsyY3RHSIt/c68l+HeXHVEJKFljux9
4OdifeHhMubmaBsWKoOWNaX/nOi10NZUcFq8NNVTGVePuvn1PMKdvNFpCEMolHr3LAHg673WKZYr
3BmOk85x5lQ4sX8Z/bji4HFz892zmkBAyEEwbwiJUXbzsrHXBfIWhJuGwP+HSrKTXX9ssgaXuHDg
+/FYoi05FB7AwEkDT9YtOjm5dxu0E8Uk/ESTnpPB/kLmvWlVzie5Q7a3KuKgncTRGPO2X6TkU8b8
YPHxZo/4kMrfRIBn+Us0mH+84lGv3L2dZMLEfXxOTY4iKkn0aEXcUlPx9aBb3yHOMfblD+Ynjf5L
DOwhPb27aRKDULj7OkCXO4mILvdmfCCU7aHjoj6zcPcZJWcyGafHkWgtG0cCOHlfDBRf0CmL0MRO
JqnCXuG9hv4Fq98YSzPl15G930uh0mSUwbULCeoVrqHdXPZVc4Cc3uFr5/r4P6l0j6bzQT9ERf91
jMMGS3jUgU2Qp1SgRR9p+HSpL6qmfbosv00d546aP4CH32z6gzWWqcmHo0JbLBjxByL0wuv8dqDi
KVLe1KZhuUhmORoLIobxD8ejW5PSTT6CSoUmy8C4SK9i7tZLpxCxrhmug3Oj8BDgWoMFltgVQ0BR
QDp7bcTbgQya3ioDaR7qDAgUOLwVjT79djnh5N5i5W3i9e0cTjDXXn/HnTQpBcxaTDbTgP+P/mNW
vjQ9jg/SEnOsyUGnUqcUqSV+tYBxCcHqWZwJN3KcBJdnDalhtg6+88Y7CRPGMVqbDkBIswFOSWw4
VoC0Yzi3NfCJEfXtIk1QI2+X8Lzx3CuofD+JHlTVI13AkOwomgnb6N5b7TlMttcR2Funjv7RwG2q
mhSdEhbRT6I+ujwDVU8NqEaNeSpPLSJGbDFJRCnqDb50NZ89JQsSL9iDVFhT5WGc2PrTiaN9LcGH
PsXC/D/rFYnEWxuA7e8I62RHcv3Sf6oejpWNQZSxaY6CeqpEuZw7SLG5+o5IvHI2llSa4YBsWS8l
KKxF6/gdrnlA4xHyLvZx31rGtqAholSpEaK87G7hwkxdZz6smNGSCEBfj0ItYFT6Lu69NWebIIwS
0Zmjt0zJdfZpJN2lkUEOCjlRhjy0qoa7G0REKdZ2omXThrF3HUaEwALX39nDOLCJUndkL95TMrE9
WwHLWIw0HzyRsldFr5JrnFt8iaiXqgNvuNKL9Ml+aP9ybNOaane+4eMi1Ij//WKjTYlQL6tgZzbl
t76qMPMEWnpa6sKQdBEU6IjWLvtz83PoW6srRB252H3ClTA/PZq62i9ac53KqiBnvdH92GuADx+b
wGPVdKD0YUZ4YAb8gptBQdLjxdFV3lgsedxrm2PRMbVQz5km7IHsn2YdH6BZl2wQu/kXZCQlsNi1
TNbipXn9VU1FmntNPOvbVw4cpCLzy9FgZyDTww6wCPvwySzdIySEqIHn+HJ+gKrZrs/xa/Vsbxpb
fQsk2mtxbXZ1SwMwiUVlfv6SMV5WFkOV6MqNBevy8ojf6n87fguhMNemi1dY+VF7LZSrj2P7nlyO
18bdzcas+qlEcS6/J+gsYwSPdc9tolpTazqtB9zQ6K+BCbHm/eA7MPmbUQxmkUd2eaM6EFIR3G/7
+TlWxO5p1z+wcA98xCPxUTfEeXPjzJnzrR+nbD6F9v1EZSDPZOilhZvXd5BbTUopMFlrtJNrLfh3
v57pge64HbjcNhALoXhDWa6QotpW5ejqXkQYuT//rJ9eenslmxQrHQp/Y1ZYVkO1cGknEOdqfnD5
26QqqLkdGI3/7s7c9OwZn0Sq0h2lR0IlLVGyHA+5/G0SBG3uVhkk6uIQhAvfbu6GWORcFaCsbQxD
MOwVoeHzH5iBJ1kLRo4y5YZrfilgNt7nykJfthU0InabSTntuLHu7yUCSz4Sav6aRWtCc14hNuzW
jmsCyxkH51DOWa7UFszpGafPFS5DitmOcrFNmGj1P37Mara4oMs0rmoI0daJhXFtx3XsEse6s/TN
JF6X4BGu+xj+yemhKFiDvTT8ut5X48M/opLDl2hZugx+sPdg8sH85QoXh6OJ2lnS4wMoD1cO3C9e
cB+Balkd46bgU2vMALJSIvrIY7wIVTcgTpBBMOMWOrup0nBSMwUhIQpRPmOjK9HNFC/FF/UrnipA
x0H8DEPbPY4ayP1CNxCYR4CSf55oWCQgNOhkUhYbDrXi4G9JfqlmLzBaaXY6x0NZtIsYHK6UMH1R
YAS9dq2NHgksU7K7QssWR95HMOAxVdsvNL6Sw9RdfFuuCeFWRTxFy6jvDCgeuJ5ElhOZai0O7jpN
nGC8HMBYjTnEXvP/AKmXIwcrm1ZRBxknlhGUWD8f7GLU6hjj+40udvYd2WjiVAK0LBeUx2lC5Lw5
rs9NPPdLsNhckB5To8ef50QpDVJQCIIrIVygQCWggkzgMfmW8iopXYIUCD1Z04JA+FgL828JH6e/
Ed3R9Ywy/ooKE641njudd/XcksE2EI56brobBr9DnUSXmxLWl+4ooELxIwdDMQuXFf40wszSiVZg
XVS6dSO2uD5xlvr/jtV3aTQk5L1qPqDch1697QskbtPwKrQdwRRzMd7Vogq/rjhQqSmv3Z4ygsmh
8+29kGMCVORXZp1ewsXywl/ARu278cY0xwibZQXJUFYpYaT6wtoDXsD3E8fEZV4XWQgBY1HG9k+K
WKxul/BPnQ3GZ3KSCiszAdyEsRlEeeIjOh7qE/JGpM4Sq9uidVt7BzxH6orDui1cIVBAcTi1Td/P
Z/mv4rN38LFqCQp1Fyyr2A30Fdwb2v+kquqy5uLlLkfTsEWYyXHhmLURpunnF6sZCFeBANpBTi1u
9iHnLJqOWuvLxkpynN6gBJN7MAgjra6cC2cFQIA5coNDwqBgBayGn2XnB8mBKhbACnPjWPssnvCg
53q5BX8zkoT8FQwX/ImqsQdvypPsRzxsWY6nm38Fhh+XNn73NiAW+M8SevATC5eokI07cdYhNkOQ
fVJUhj28I0Dg6n53RZQHhywZAp+guh4IL53P+QrZhXH02/OJ9KNKC5wO6lEbcGf9cmJZLA/A6/mQ
9fTk0qv1Vd0tc9spsI7cqlObqKue5l9pz7rjPqcJWIa/ec8l19PI5WUqvLKY4bSNg742QUYv+niK
gIz/onim5+mNTRMEkcTzUZm6tEX6jdWx2FPuDJA98qBbwb4DNdxV7RnbdgSj3DlixqyoKYKzTvf7
/bvb3k62G81AxQ5i3U7AQuGClCAXOVHekOteJ8ukrZNFhzgFnB2qo/tmkTl0r7SKrpbE+TLICPzN
8RQFGHPEAji2XIrc6lM+oN7XS4PKfRiNIrH9FXAWG2PWS8wHepaNu12L+tAFLKKRlZCrnTXzINMK
/bX9YXQofG2xZB6yDGwIE0V42AdEtG1ruUdcTjSno0zimBCJpxfDi25NPrFwH4d2HmpA+LTK1M+V
yS1VTCHv9vu5YtFLyXtYpQLD3xlYvVgh4chInlr9RQlbs+gxyE1m6wFJGS6fahJ3A7VoP1RTa7jI
49N5240y+JNY08Bh8hURjrLCGnPc/9Ts+6gMUGRziEA7Oea62ubEEXn42iFUU5jjOA7cOou2jt3Z
jGTlyKwb9W9Yu1YGTODAWm40D79l40nmYCkQFF4TbnhHr2OElVlVtwtkkCUhgw4bmKODdmMzFaW1
AwImY3HR1ZZWHF0f54rmxdydOqy/IYIq7f2xzGC4alq7y1ubFQrsLo4adSjwA1fkMJBr4tqDu8Iy
6Ej0LPxSy79LGsCST7exwzseO4L66NsY+Cy6MXAo1iFVuGGHjj++y11chifQAKoLRpUuXLKnekBP
mLpAaOEbkKtK4ptmKDlBeAK8KrzIpL1IER7n9wscBwFWDUX/0xALEBAZmjXbHgKrKNtHCcfe46jR
SCGuoFvGbBJwtIjcVyuYSvkh4yoAtRvwWLbtacAYpD5fEI4YYkUfPrVbWJlAaW2cRW7TnYADC85C
KKwNT/QBgHImgrgQfaLtYjjsF11uP2AbrvaZoJDf7T3pqFJtRMSS7VqsVL8OnnBSotImeGubEmfD
IgKfxH5lBOiSBqE5+E3MpSWwmCrvX74vZUZkChG/4TI0dUUnDDgpeTogYNSFL9VVfRjMNvnIA7cO
sF+62/z7YQ3mFieK5db4CGw4HBLNkpXM4QWX+KTwXnPTaLdGnfF/MIPcMTbwYS06w1DV1bu4a/6L
ZY4U2yofj+HJmBTIbzAp7aMm910g/kVPlKo6jYy1r4quRgGaQZV+SzgT39DJI9rxlznEA7GwNNjW
5nmhamM5AHLU0xOjK6nmnqQWDSCJFpCgPGK7pZxfpmBoIwkr660hUFx74jkKCfXqsKIO+BUhk46U
md1Pxc/vvVuP7e2OBOasztLf06asNHB3vA8kL22zK0fgPAE7ZKagTb/LuFUcYeq9yYX80LjtKhH+
7CUVrGBuHmsZP+5NrqG25FZgUGsBVoPc3Z2f2e9ESCn5MJNs0EXoz/zZgKrlco4E69rjiTii/W5P
mB6HeqUlpKN7uWZtpPFbcgJvdZjO5RX9ajUzZwW+D9LU+W0i39hJFGFzJsxcO9XqA7gXfTuw/vWH
aOxtHumCRbOQXwaClyOvIGVreXgY6QYzoyHZsjBVLddCrEcbVZnJ2tZCl06kwke6Q4ZVpjzhEZyh
xPBnovEun4B2p5jyXwE2/ZMcpQbYifHcOr1e2fQnm3N4Rc/toU+YMf84XHww45mcnP64yjWrXZux
R6LrEBxTghrSx2LwlpjPHXvavnsC33E8ofh+FiQbBevqbNe8qTAxsGHyJqPCp51j12wlKbQlCBDg
B+p4SqVzcCTPqvRXolR7tNTCD51/SFP9KzUlbcE2PNzP5hzfCniU4qdrLXVrURrrpfsKXnK5rH1f
DgnZJdv5Ndi4sGDhNWl+v+FOYr81Gtkqeh67tcod/7+/eTpBaczoPZh7N+nGgCE6KoGghrOpXZRs
TW/ajDspha8U50DGaB53YhU7IiTj0cbIpmtik2Xp0HnNdZ4IlyMb3EEM5hjR+AIEo2kws8LBkIve
uqYcEo+BviHPu6pb324ul2JNEEVKR4/Hel7avRzCuaw6X9PsI7w61bBqL3Rz0+qXAuKqgE3yVwts
hvhz4FD/1eRDt+IL40AdDI7ZuOCMAW2fp4vfSXgv0GKcIQiNLF1IboUJ+Wk2To3pNwbhMZTf3CsY
4nCH6GO0/25tN9tC3J2T4+h0Xlk+IciSlJgVioxaXPUqaaJfFIF/xA0WLo/t/TzftP2ZU0oEeKGc
lKrOpO8ojKUmFE1FKsdJ3nF15THd8B9Fgt7IVQoD8YwqkQBcm1zP1/zBGDMJIbmvaWxTd19DMkdD
2OKOlYaMhealGi75IN1l17TSY3nBm/Uk6viGluiS7JKJCJTENpiNeD5S/yPqcjvmYCxzCLuJCZ6i
Ck8tlDFwZBd29cWWa8tpX6v8ZCAM/R6F3+do2+9hYlxrFczCSfWD5sy2nfXd1TOHlydBqegtghwx
lzMQIHnV4EOvoy62pplZiU90RY/oWn/QmuNhiVvcfc88GA4ikhJ/vEPQTg5PISZF1bty5JxvC3jG
LXyEi707aq8pNrqPplXgCpssvNojuwdUdbYX7G8v8zYvLFSJ4E4etaxI3/81PBOubvSXCuYMVYoy
/oZoP3/gVa5qdK+kdGihuKyvtJwcTuk0car8SG+D6Lq4yB4NfmhH4zxp2R3Tosq+4lXUAR13f8jX
N6oUVzpevDCg37QTTy9aiziNpZNXdM84YSwU3/5vIYgBOvB4qTOlmuVi+pHFOYwh8BMdeX2xfPYW
QeiqKVzRGQ7cIMWsCFUHlivdAsuxAYSTtULdGuXl1+paL2zcHgQqM43oVFHn5zNsScrnbWQNeUUW
MYwryfx6JV8ZmVx9cGgRfPTan4WWkVO6pCtHCJ4ZdXfYiZkT2dhpZBVmTYNLOM7MD+Goj4dUb7F5
hFNtM/ees9Qk8iIY0G5It/jyPRfZdlRF6aJZkdfo0l9f1t2QgXLuuK+Ku9hq3rOkkPuozSCakPdi
z+ODT+3xx06tuyQKNhLG818NpU8dovjXvtSNYn8F7NjSprNfSRi5Cg5ju5JLySBYBZx/33ROk2qq
4ek7/TylvulYczj9e7ME0XmH9Xmxl/P0wjQuD3uCT4rwcIToc98JZmYEL7DKVKgMCayN57OXZxJl
Nm7/HjsDGCdeDY6Jva/k0gOiuMuEraZ2QqK7t4vMKtmgwBv8o6m613fdSbUc1w4URE6bBJMZtHhv
q/6cuINx4FgkPeGm7BAtkLCUtBb+1D/mRFzk4bQONNLyr27oNRNByZXqhme/AeLyo8hqjq4Bo4YJ
iigcz9o1IOq91iubUKXLvqBrNKBZ8+H2OZ0A6z3B+hbW02UR0En6VpZSMyEnhUp3QLXJsuQ1b51T
E7AchysbI5WKUdhzeyxMWSSW695kvLekzHNJ05VZAPpLLbgkmRahBsfizRDqqobcrzZgorwejOCW
Za6o2lToHRn7bGshkjmxm3IYLgTvBLpRn7E0L8XSTc5apFaKP6M/blCUQHIemloU8iI0Xqi6f/0u
qcrMj9YNQU0i+yBoK91ujPL9QSe/KaEQvS6MpuHUXEVVADTgGv8ZgPtfttTfpOWT+r/taDH9vnj0
guuzgbCaiwDohQQrVf+L56fmiT9F2ly8qRMaHX1OyTyyDhO0jdfU/6yFp4YxdN22QSQUF17RwEb9
2kUPKXXnv8wsg+Jbdj5EwUiNn1AHODaR+Yg9AlIl4+yVMm10J9vgtPj2lTeotq//ido24RAqFKMs
PDu8+5R6BkKoj3C7AL0msCV/dFDw8Libn7JHxGRZdoQ73pYt2IlNbIZE4yF3UvfmnXn6RQNy0Ph9
uwKhOIlnp4h5fs+pGPyvMDDhZfaKhJjlUMF4z8H/kGMDoi+hZ7iJ1H7pKtR5a+yjJcBR2fVRhieg
ylXnNt8l8ZKJ7hJ4YiDDB4pqg8K0udLKZa627DIG5EHPETfCqRCnGcc6grAuQWNQAW7R64/Wu+N5
ZA9azL7khJzwcx/ZpWVGTUS+VDqioCb+H65aJ/cQ9kgS4GgEpVlD7YKhDp354OkOng6kZOjW7O0b
6/d17SqHpDyXxy6XsXEg9UXCgsnVkgW5c9SGv42qfQsv7huJxQRqH9uY7gP/cdTfN8rbC60DjlrV
gslhXlQ2AyD/zybDwsTw1Jc+Crmj22Gn5Hj17/OE9nBNTcYah1nLX/8vEh/zjqA69WV/DVawToH/
VpdCbSKnFR6P5cEff8TEOy71DpbtfywkIgZ4RJO2D37zbaHzFOXuZ/tBdjeG06F60i0s7gM9kIz0
NXb/VmEmABxdZFYMdTEk3feMEqPfOSKpSPYmUplvnQlM5Jx2NQZC/tQ2ETfQRUW1co7gVo/JYya6
ieqrJvRBmJRjspaxL/hu7bndElycPpjiayphlU/6jUkFXlslFdd2T4QamAJLHpyzbJQo5ivgBN3R
l5Aip5wdljgr+QYwJrvapMKQPY8nMUl2seEu/vodrcGOlc0Xn+t4n1INgRhEIYOH05fZiWhG476Y
aTxPv8MiTlpGcuxEFWXvP7MxbpREc1NsoQIxri0OoY9M5Hya2khOuuaPIcAj2fWCaIFEg4+Eq6QZ
tB2i7Fym2spHcz/2ZHSGjLmkwvi4Ou0g/9fc8ZnQXDyWKpNiHIKIPooltrqPHnMv6GALWJ48X2nL
tz9EsXWJnEbkQQhcQP81horFMmq+cedKESvJRxq0NtffxT93DPP9UtGB/wWXn9nqeZz7EQUfzO3a
F5cnuL3RbDRghLf0jMzni68Tz46j/iap5z3dlA1m5YQTgOKLJ0gSR3y0yZ3Elu1jBAgY2jd+2SZC
Wb4suZPIIQp9NleAZwsLOY+YgLvRhFEnSroBWg0uqsZHpNn25lloaLiJ0S9X74pVdWdD1aRTlvmr
lcjSgLVRZV5oo7H0FpYZeJCNOZQRGqo8aHmZYfYCamQaSn9QzZzdRO5mFodyYKGJRCD9+cAMzr9j
/LcY1hbxDEb0G0tCGW1ApRZaRQ6jedNvsbLeS92Z+/GRBmHHPQog0tIjhaubAElkjZ2hYjEZBrAu
pCbwys+yGrCHs3f0lQU9Len+qDFfZYBY5tIxBMVuiteDoc3OmtaH9c+39JvI7vcRAI2HJUjpD2u7
kFChEcv/GRZQpodhGp1IVo1ULBMjHUjyCWmabPfObNpEvuN7el2Q7L7Xwhj07zDD0iq6QxDHCzKS
QMUWgV8ARsDvYhiJwjoKyQ26nzbCU/atSq5qnTca4biH2pWhSMpfpDDYPykr/xmbQYAO0ZiHlnmG
9ZhITulG+vZfbMacptYF6aTbsGw/9qtyse8ULvcSScUGtNvoh0i2SaWYLYuTj8f7/Od5oHHUPBTG
r07OxPf3VJ5vaRKELZ7iQmC3f7B1T2Bsr7tJ6HdQvoHO35VJM1xn2w6p8LohWP34S2bCNF+dlj/F
ebisbzcgqIuUA27T0I2fgdF6aCo11jwEzvr7Qe3DFN9BmY+Vu+SYdClYWQ/iNUx80qooXll57sqs
l63nKoY/Zr8oN1gfitRQpOJUSPY5EfgIa+7JMp3fVnSfkFAGwe9QHhldlZKvHIPpb8BAEq/iM9io
QNiHmNM/7DCsG0cQoiaRvFbuabl4MqSIcrkO2V5NoGJR+6I012vtjDI6pcask0h2x+ddFn1Bt4AU
iKPxgLi03NUVKuGeesN711LJfDG+PeAF9LTUgBxQQWKPqxX8gHYtajzspf94ecB3PvAkFQY2L3zj
rAQ4Lzp+ehjg7Cg9B5mVNbocvd9ZLPS52XZKmcbXCYuZHub9WTgzs2ZAHI7G6zcb4YBTZSkHeNP4
z4nInPQMhV5pnSXZATcrmChEPhF0+Gr4TPeosqtGpvGe7wKSfKRrLfY6kUDGGdnzJEOoRMtujbKU
5Q8YFfZN1FdedjC3vWDRWiFFuK86+MjfPEOuB3V5+qW9EGVhy7oyHKnWtmLQ202CMAe0hLuMSfO4
CxLiC6tlafak+1cGD7ZTdq9rkC79rFSVP3ZNfOJDRQ8TF3iMu7ZcNNMZr6IIRvsBSN5+A0WLaC+I
KDHx9Xd8nULTuW2XNiMQJmbdwjWybWShxA5FNOg5vEI/UHNndbVfB40xqokbQaTexhfC3CSYzPcp
EcXrhM+Hqa0ySExUP6lidopFWyvHRnSOEFMMV3KU7M1n0/Zagfya76gmPGnZdoVTa4ludVmy+ae3
keVYfT5w2FGbBZ/vBqBYADbz4zE32t1Ko4zJQgbjzDNZqCHcTeaV9ikEMsnEMOb+0WsbzjJGGuHv
Xn4ZmIersxHOZ1EXUmLZK5CXqcYwtgGcio1t3TSi5HprY8TWVhXA2/22ZNsSVsDc+4OEzjU34o72
DoQNr2j/LnTctV4l+QBhabQcn9i9yjNHHWTx0aRrcfJESCia9eNfpYHFWI/WEV7KhRyPc4jwSIXM
GdQmKsuQ1RtuIqri1LevsuuNNFOwd/KqaNZdpsUmlq00S18IZo7Xg9dQ9uwaYg/OmeMAGs/iIxCa
Uke0BPm6b/SFc8+Qe82Xj9nsmJ7l2d3ndbpDk9sLo38bcDIMGqO/q9aRbJLw6/UWY6DMR5NT2F0P
Ed1XJZRIe9YmuaxGo7wleSmUuAmIku82n0xU2eSB0LOjvs276qbSev/oUeopaxkIt57czPOIMgBL
5jJV+5yheDGovfsYmxU3Cg1wNPYzRDjFwd8JkCXIdoXaHNiBG7VoVTJnud66Y7kwbrZk3C2Uh4ED
EF2XsaH1ErPqaQIf0uL+A7+kpul1LbYTwNinA+4op6q1OUYdPa03X1OWfJHv6yFlhj5xXVzr5kgf
JEC6fijON7ARL1Pi4pWD/XGUpIQysSJjdclmAMZ/keEEknvakyWVDQOPPPXFdkpCYOoZbTEB3RhW
lav4GSkDlCMpd4EDnR2ES5QmRN50JDcbIEmuO+amum3YGS/V1PCMeahRac0e8y6cdSXG3IZtKjMN
VTNtk9IbNpm1t4ja1528YPbpTjCq4IuptYSu38dUKe1Lp9PAl+L42A6Boe4R29ukB43XUNHYtWG9
hyD2eagDLMQ+G2TUMNsBWo5J6cllbeqEEDOv92ODeCGde4n+2lmFav4ZLK0yC/rCtqWq/J1a4MAD
PrfgW2+gt5A4Ni3hQqz/TLhEQrJdGLLJYYKTm/IXVXonGd0wv7Ao+AHdKDiQ58lCrIZyeJFd2nHW
osBo5QkWbIj5Ijh7WWJicFdNn31cdsThnPG46DE02Hf3zu78VtL6nu5XUiSFuUYav+8kP/WCnuo/
O6oChfsRtoelfe3u9Imyf25duW37mqfQge67WLzWAXR5A2qd+3E0DICkw2Z4Y24EghNtJa+un97P
1BvRj4oC8GiwIjcxZ/kGRhZbK7hmUMBjrH6GX4XVplnFhfOgecYempwQqGAzwRfEyNSGWbgJBVne
dPryxbS4BuQDQi+80pvTOJKWh/D9vVawHzWRON7jQJ2gCzDvrsV8LEVTMPE4xz52KaxR6RoA5Ojl
U8BiZ8YvQnU18w5qg278Qx/m8ntc1dC6uxMxTowJMQdD66O7el7NOcFDb3+MPy04g5iG4oUYopWT
pV9yJVaZ3OgzZI8KVccC9//hsUAh/qQoLH7wzG7P+O0TaYmUjeyj1FzP+YnOAnousUVf+DOla7VY
oAfc/k52bvXbiJ0PtaUQzYf9YbVzxj9Z1BFpHYVrsa/YDONhL0tFgSDF9WNNJ+9MnZrOYHe7KB3A
DS3htYmBqJhhVv4IF3W8WMigP7LWtZljkNP1/IbiQcRLaejq5a4Z/vSlo/MXW6A3Zs55p12X4uqq
vYW7TO0DLXI5Mom4U0tHqW7D0ptFVKiIdM4tlpa2NEFr3X2pzhWRUx021/LQBUkVdsiaSEM+UhLE
AaWn02TUt5uUWjCxBFAZyJml0sE6RUpnNNHnXVvDkTWu91oRBE05o5I5/Havw1IlngVDrugF+m+B
lOEtC1/cPAWP1nCwZyw74sdRC1sXcx9XB03eGl3s9qINZ0mGeLU2TRQiaInG6SqrKEUsL2w0EDQy
/lYPLljFVgS74CKaIbyEtv/kAkY4dL7dU5swLJ+prb8m+p3uLEkvq/g2yGkVquJEHdG2IT/06/qY
z25KvHhOVL/dQlly6Wy4JV0pKWCtRZKQ8zlxMBnoxkFwfkgtyreldgEpcEOcHNxZJ/C0V9uArGGF
LtjpBkzPm+9kWVZtybbDNbV9UhOHHp6yrcUh6mnfd0+XO3F4evy2miJ+KBI7UuCncqG0HsTgSrLg
SCeMp2wIbbkWYDSsZ3tABpcpbJSaFrDRThmduhzvB3NRL/ypu/vvIIX40vGfImQYfsMiGh2Jr29j
3P7HzbWVP+JcPvsvcPKaCYHxn1Nf9d3/jKprQZ1oOdlcQw5rLUgSHxdvAXDnkjSCYONoYcdikqiZ
m1LYiF3wFZBNZsYMc2bLMnKTyR2x1rMhNjux5yRwJGPioOJAtrNfDvF3pDWVqN6pawj5Tgc0JykL
ujXxh414hUAUoi89T0XCM8M+kFHH4i8CBMMKD9HzF3xQCig78V1aEjiIvVSSFz1DpWmUS0/Ttt5f
fGM1/nr4gPd7sJABEq1+QuQkpg5AvLvXN7lMxfeIIR53Dd6Q5okHELzQ6Kw/8QecJ+0vYI5AYIwZ
mYjkDLmDNoFQ+RRxAfQF/r6rb4fzEKIE/byI2NcCwDQF7tHePQ3/peL041rFS2ti7RDdzOHMK5eJ
y3pByE5GfkvR+woo1Wppe2XQix2fVNy44xu6dLKoilHgnTwsFdPTrhbFdQvyrGFSeKceVZUQnKYl
jpq0900Rh64ABGGSkeLHFkxGEKpFwYo1jMNplJA9Jb7/vlbAfJUsMd2JxVPYhPoZii84b1TzdMxd
x7g1Tup0BYng9ibiTvgiDFhNyz2/JLH5GgKBNozM84Zjuj56UJkxBI6Wuq+UdyQ2pdkJvsWeGZmJ
2cExNyIZrSu+B4jdWf1Y0G754qiHRyy+SBU5SkRHc5sksvZ2UROjHicylc9shxmKmybQhgZtm1S5
UbFKEdttTG+APU/rfXvoWLnIgy/ZiqtMdDWc9pk8DKkyKnvyctbZdGDHZs5sfuiUx3Jd9NpofSy2
bwtxzrblWEHefjJ57Qv0fNITMvLyftx+ZN/UaTSoleVOHyYJ8UmH0pEmvfGeEMf1Gc32DSJlwgSk
u2liJDbMcqpvU5YxlvhFDk5H9kJPb9fOO8kgQ0AnykAXXIVcHNXmdJLvdc8zr4CNrApRsdhXG5eS
cmahtZLNDsQ5e7kESZ5F2EQ9fQeqYnMCUND2zMHMNpBykZsKLjspRj9sZGUSZCepFefaUKTDuETF
oOmjQ6DGlCHqRhgtHQqEFpsET6k6wAx0+qSniMPce4OFIiP2t+yQsFS3P3FIzFKGdrWQoeaNM3eq
DHDyFPumRzcwfSsCeZip4vOjVdY1ia6oVzQdtwqf1oqmuCgouAMDqKlQCHZh2Cjn03S/2b3i1K71
gzFvjgiBEJAxFvORmBifTBGygYmPD3gY7TpyMCJph2k/GKWKEcpWRfED3Rdw04nb9vd6hsleEQ9M
+uM89TZkEiC3/Wc+R1mkMJVpao8IyNedSaXdx3K9bQg/yPvKjU6YbwENmo+jWX0YTTp7vjoqDueW
oDsbutqDzoNyCBUMP8R059NldKKPGjUl/OV9TyBRiUw7fLn9MIjkQfGXHapYEvJW4DLdFCkbLF6h
uBCaGFmcOqjyBrC/xrbjoR8z0XZ3RaNb1SABZPR+X/r8ca1VJks6wM9yMDroTrxy8PujST49+pJT
P/JUx1v6AwOd0f/xAb0E+BqYvr0dojazyUDokUPMYbEDRyQo4sOBMZPxTlPDNDs4zUTip4ajf/4F
IdEmt/ab4njCANjb/uYBKh4FJafIOXotVYUHsQB208Aie9yYWlN3DlaZS+yNbh1Em37GBjX4+443
DKiA/mgcW0RFpuTcKBWGfzwKX7q/HdEvaP/tqx7mLYyU07Cjm5V2It6rB4OXDXmKmdP2hIG1awX+
lsKO1K3a4VT0HiCmEJh4zhsKNpGIydHppOwIe/GdH1++CQG3lw6Kxrdk1c1v6U8EFM4iIOgI0zF1
hefa4dxq6U9KiCJvkRiEbbKZBzNxCNvm52fiMIGuCpX88L342vGO9K8DHBLQMQjkF6r9PCV5ChXo
HRSJyltxCdJelAiFvJNDDXNsOnWGA+QO3wLUjWK3RvhJH/4DUXzgMVvdCrTBWbPdZZJeFwibFP83
MGB5Mqq/XfFVGdX7rAOedvfZrPt+mk1Ia9Ab7+Ezm2OlSCe3iK2tfwpqhXNouALKjDpqFTyCAhqh
IKY9DGdGz+DYstMW5+VzL7TICv+9VAGBWcWNRuBlw1muZOVzX+hRdlZl6dYQQ6CljrRIFp1wAglM
NDGEkMjeAs5dS4J0wp3ye0vCMxbeRFLCGwSOcjumhGsG43KCjIC6EmOcJzc1RlAa2JXaHA04Gkok
5hCDvLmr2SVdV/2IIRMTgBOilRPq85VUWhvFs11IFkJAJgaVEPOP7CZOSkyNrtlwhHFSJm+LWL+W
aTJZ4hyOSMZ6yUK9f1RwucaSHBmh60u4NKXqvVNzoDeD9bR4tOj8calSzMenDTEfJvTdKrXuaAfJ
UahbMLSdZB6Vdp9APXwxbpU9paqgSVzhWjcIZvuAHMAEBdOr/CMN1Hnsu0x4S1auefRruflsL9oo
xF7PUbLoqwwLfzvUyypd4G14g+BRMOZI1UuuyyKoOR7YtUUqRJZJlW267ojLTVN9Jn4XIKwZpq3H
aN9tIvXh/DrImHWYYF3ql6bhFfhTgw5fZk+RXID30p3khUm6vAsKxeQjKErTe2x6cnqroy+Jr4oq
2YJkpVkHRz4cg+fTf2qYlU2GOF1U5lCButVPI2MU5b3yr7RvvJABE41Y3ruAloZUPBATpHP2CJHk
/Vz5QXesPoR/LxX708EYPukJ52MJZ+GxyiXAzc1LXQVopDrzQbI1/bYaY0fRRawlPw1/i/zrzDwr
q9/EBki0K4nIjaEb++oBHeIKlDrdoMGpvhKiy4oPYVi/ON5efHXtIQPRz+q32cgZlNjAfOImZ7g2
jHDeVhsheFPzsOpDKWFDvJlM2g/AKwAE9DwCcaawcVVRpvOJSXhekC8Dv7d4qtzrUtMB5tAMngN8
NL1cX1pUPjuA0qhjvkW0XpUbDevPU6Lv0PuhJjZeoxExJducSdAzKhu5Lwpia2Vl7fGgCh0VtkXf
RTTkRq8ky/+Hr1WVsyPFLWBLkH65UeNq6P+oxXmmjGE2FDQyL1qXE3C0mI250hA75kVbwe1r8cPb
7Hv5/jdJsmF/jg4UxbRW1e6bxQ37V2YvzZuXseYgPKm/LVYje74f0f1z4VY65UP2ssr74bWAVcqz
00aPhbY+nJihrx/9lm33nqcBL471iPZ+30UYEydTJrcW6rxT24kugVNa0HODCGgLc80/UM8bjmpf
mKJVLx5F6+91fvBD2zwmDBcgBAjPywbSU7VSJAJKIKIfkaciMG+U4y3U1gTDzVn37Lpou7lX/hvd
Sb/Nqr0oWS7kUhAJ8d5Rbisn+n2b7TY9csZuY6O/Sosx9gj8UPvveTNVqvg+v7YsOq9Pdby29v6f
jF9dBsZBocqptrsjjvz/7K6JkgaZvCpcK2UfuSn3vHNhgC/rftwXC1r+p31nDzkckwdRJ2LmbAZD
1UwlUaXiyTfEQcphhRMb2qxZ9DgR9BUkeQykRpwiNu7Le1BfWb0bGUUHdw1Rx4iRau3uRTQLaH20
L4+S0IzTIgjy75dZ2Dj91dYMtV3IoiEA3yP2kPqhhI+pefRw4zxnolm/gSw0GNtTphuhbH9p7FNR
hH+uo10xCKX9aD/2r8r1yB9e/x1+7UjXbsyS0WvU8fRL2QNujl2GHAZmIMWkV8WNFw9iWhSWg757
dsZt1fFl9usSr/jd5JA2TP0EL95dLOuvf3GH/KWZ3SzEdfV7mTvjmb0sEJ65Eb3KXO14vdkTJvu4
jLLV7XXkRFcJj2owjhmBvlx2vj54GhBwWgdmFNRZ1Lo2BwexU3oZ+zm0PxlE9N+oyS5orj+2Zp9V
cuYwcyze000DoXByiYxRIXl1pXyygtmnotnMiu70bn85tNiitPnUZ7QmqrkIWG4dooPeBoELY67Q
qbWm+zBi9VOaMAkLPReJIz8zkHLVoiUbqUFc32Pw+jNoZSzsVwPVinpsc2Zv7bJ0bVIG8lOiDReL
46cDIZpAIsTD3CfdefrhZVigUZRlHthm8Bh1xYg4yChDbKhQAdc/ZVHwtWmBEa0YUVcrGwNT8w/X
OTTBZD2ibafthp9qvjWGtdtjsR1Z3bob9DVh8wOtM2w4c83D4zUNAVN8iOr7Ppb8Ur3TObQlM7Wk
5cpTy7ISddCbevp4uXUNOoC7KkCHio8c1DFg74stgyzOIwVdzMnEelhjV/2Fydw1Bp0gBvoegPOl
x8tQu/4ZVcNTACn6RFOn8BAeZy+vgNDzcBpxmEEz90Ol903+TG5nC5Z9iFBA18VAE/xDyRNx0++3
4S63/LmFGGFJEYUB0hWxevMxH/K3NP6eU0Vytqi+KZaq398qs6gyVofNJTnoAv9fgzxjdzFBcwq4
qcF22Joi7oV2e2DXp0aTuGAZ9YVx4AFl2rep6ge7lRjKLx53qQMBj9OH1TvoVrYQjoUt+aoDCgns
lX0LwFqfwVd8mM4/zw2Jfy9/+vrMQgjVFlEo62ck45GidPmaqcoQW8wpjT8F7oRGC4C2Q43/PkPq
zzRKPIPWWdCHVTyV1w8nUKnjik67pLjUiSaJyv1NjLvKDNJPaKGh6WLWx/2Itp4+ixabaYXG3isW
9oGR2G3601dp4Y0uw69/5emjgC6bX66S9d5ZifyDJXp+2M81Qgj9IDuuY1HblHOc9mlGDn46KlIV
xidr19lXRVegSb3uYQCOVuSwbS5hzbG4fB5FoFcR0BU1tPeX14udDJr+XUE2Ddb/oSqGQBphdC48
sTfF5KrHnFT0yYytYZBuFEXbNDi7NKCJgURgIyiZcSai3olZaCIxNFAKjnN/RP8+E8LqCzcuuQK+
5J0xsewEXQ+Mke7l9rPVsVxP+rzOggC7ZqUnyGbtXsKv3ADf6TAmkMFD0bsa0F9Q4BQh/GdNITDd
Xrhr1zS8cTCneFcy+wXjy5Mn9AZrFS6GVU1ZWWAkcChAup1Qg8kAHjiExsPpeXb2Icqb6sjCwuLO
4vwWS/slAD/5xrJTAY2B6GZK5hB4vrqkD2uy6NMKp41CFBKehQrVvwePIuoG37Pf9V8reg9z9QeJ
IReI3l07t8vSsa/KvpNd70I5mroZz83kZAaysRqo4fK/Ves9xyH5sHmc6PgCMfygwmXiz/yYjhnA
CQk1O/MtVbS0X0iHjsZxZ4wfxvC1OUcvBWmGbUAxEM8e6dEvoTRBWw8ID29U9vE7YUWv0zSdbUdC
F4l1BLm7xeN6FqDxjABgRH8kAo9+zZ7Bk6ucDSKqcbefGFsKUKbMgyxkDsAk1o9oLgNm/DLLzpXJ
jrHNKAJcjBBtl+5mTo5QOwLTeoCF82L5qwgFsdXXtxKr9Q7lcpxyxIwJ23rIKuScYzu6kFaC3tHa
DEP7Krb80oihhNZAx0fGka6uzAbUytK/P8Z0VAeEG9ex+NDcKBxSLDnpGYnpYAE565Fv8Got5N18
agfsvwm93Ea319V8lo5obIki+z2LGNv71JJSft516MxIZgVMXOqTsSEtXbduDLDKG0JY3jxu0ttI
WPXnXRwqnK9/D0Jw0M9QSBhdHcPvllYgGuOHbP0Wl9L2eZHXE8q0iymBmEYmbNCQThZtH7ViWYAW
JJ5w7jX+f0+eChWi2m6JtgjFHSJTp6aw+fJvMg0UNfp1M1WdyWePrtIyj/lovigACBHbM/wdajIi
K6SlwqZgfSvx2U5ZzeWoOoKlOX4SbVq4CPFHn3vzTXm3dJpacO3tPe5sQEsV0sCq9OhokNQzNtv1
9g4RMDnvaNcrw3A6KPoi4mOgoX/dxsIzaTFdOjyZLTc6A8npMVmJDLpFimUTqWO1zo9dtaSLyzeV
XXdQpGa5G2Jk0Z1UzhlA2rdmPkVb9oBZnkKG12EHoti9AntVnNXCQtcRiE1hMXEpC1pJRmcqM17k
kc12uDEtR7Y90MZJMs7TUFgSBttKqbKzd7ppp9AjjWmo8ztQqpXIKypkT0tyhcyIPadKDCNws+3C
+Ozh5y2RP69a6ZkVUR5/hSAYCYs4prC6jDW65InEvaXhFiuv2vyu7EVFuTIzMM9fwklg+kY7tJrR
T/Pias/aBLXOyapXbvP5ZfM+TrcGNEGmjVxqaMpg47wyMqikieeGBRGBwpmp+L5mz47CxfmOVvXJ
aPpmE548b2IddwR+WKBYRcpeQP2DHjb8ey78dOiUYAb7U003f057vg9CucimA8jUFjikCDi5sjOz
Alfy2lc93jSFzrbhCdt+guT5jugZbnuKEGo3UHM8lRyk2PQzIK+X1bcZKK8deajZIHwzdlMMxlQp
LTp/lDSx9Xhe24T3VWwL2jmWay+DD68GDXrHNf/cjI8veHjjEXUeL0PRNI8M0K165amsUPDLGlNK
8gZIZimwAKc6B9DyayPEJxMZBpqi7OmdxgkJF3R8uoGMFjm+Erjlb673Zde1NJHxUk//Dn5wuYKU
0V0qGTdGY8K97exrtJOnDyQoaHObBf9oZF3Tk+3eorv7ugKv3fJr8yb8++rUInjK64gLEwOpqwY9
eUMQq1/4j541YM+m6PMIp++xhQ7nDQn2YjugeAvaFn0v+BcHz740TYuc5UNnJffGfI/kQ6hukWVW
I11O4xLBvYswJlwBE9ADiAZQfLLPZg3zw2O5v/8oTgpxnCr0tdDPTKVeuFSptKtxo5JPcGuTra9R
p0HpLg6o+D9K0iF2TDejhfDF8vJQzpPYykOblBtb5r9QcoOljla1dgdUa43BmHM2NXWQVY/C0We/
pALWOjWPr+wWqFxhAV1xWwi2ndWPX0+Bl2P2fJ7B88CotVd3QnBLUBIATghH30yYjLJre3WF9Kz2
Wn232BEHdJ9NQUUH9Sd5ZQeGhxnjBE80l4NLBPy0tcdmYxoePP8nIfFAtLfgQjTFzVICzk46l1wW
OrAp4Arv7h9A2j1hLqUm2jq3/6BrLwc/HfoN3GbBkCmGnYhBgvFy/JKMSytKLz6dCwmu+6RkvTOr
W89Y/Uc7olO6pzANpi6QtEm/nN5XEpprYIw7LZwHQ4jWrg3ncoS2pgVAdmVATxCNWwLT3Ni7R1hB
BtNwhfOYrlr43RMzRB9SwuzygSETo11Ph7PryO17D+7lE3s6iBkxBDvOj8Z6FEHWlFO0/YuYRt+4
l4jQtGEcwOieOUjEILEoem+jwtRJobm7Tm2X5MeRvBxpO/ynk4F701iFOrqSy2BElhSnNOk8F05c
bE47MNKXisfULx4JFFk12XK+PFhEWQ7PfEm8Janh/1cGSyOJgu8iMFs7SvHempJBMWjdTHTmo7Y2
EjqiAvzRzvFuzqUz61rOxWdRrC+2trCKVvncnSlIm6N4tMDrcQhL/Hdi1wNpO5vr6QRfyWPtGRCQ
kAAN+9In/9woOFr/S+r0TgGaOxhk/cWrjWuXZiqUimV+ODjbFf3ebGGZ5mlHNylbmlKmIAfhpzSS
viMIc/rWLOWRDXVp9uio1E9/DB+iwELF6m+u6UqrlGLHUNGMqhrC/9TqYBq7xcPvz5IQs0jZEnaF
O3+5E5GLtRlXOmSYtYbY3/8O9sUSrIFDjezpWwm8QQ0IAWJ6q8gXncChIblREJGu25j++zbykbAW
jD7JriHz/kRBHbhL9dkSwLHolSji9/Y/ZyPXeIV2NW9PM7mvFJDyFzLSU91MGVwsD37qkqhn1ogA
6JuhWITag6ZZZ5tOG4FXrVbbRAfBPL2HZgf+tBNFAXin/bXHaZmxZYjceUeMZge0oOcTrAxH+mbW
GXTFeUdQwbbR2dg+COmnTwZ4qZstmV6gOSMCM4k8SsNBeJZOmUWU3CEkkoLarmzooXnNTiTyFOy3
IJf+dBWj+UDkFjSRMb1KaqXpwinW4Hn6+aH2JSBO1hxR8C8pCtz12NbDlIm8muO8bHl5O+GQmaYM
Vlg/yOYsgypdPMXI7lsJuGKMTjcBxVnm5sPju57vTEs7g7gZDPWG/V9BmpzyBnySq1A8zZWZlLEM
Nn/waB1axAt6k8M0L4yFILbBQ7V1Ed+lMnBL+neVknMZfq/UybZmqAAUUm09zd+TyTHyeVvfTvxs
zx8NkvB2ANrz+BOZFsNfg9BZDvVtXOtr+4ZMb+bw/jmnTYQjdj6e3fMGC6WQ3YbhZf2EsXqxbeJH
YtX+Vx9/i0EOw3bFEvGLg1WMpOHE/tFK1D6idH+jcYNa0dUYQ2dQKJW66PvG+MZ2fYeJS6eWkVJ+
3P657nZURu1NiUmWmPcOcvSvC12qlPWo5lEk1JLdhceSyobivtmfVZBNl1q5x3/WZulf5l7g+sSe
5vsLz7AWxemes3ksAUa4kTwLHYpO5upnEHh4KSjLrZ0uw3ggSWfVQeVbvwEyFQ+etjs5d19dqZr1
sTz+y8CNTQtxzDds2RzsnpSEm5SoRmHkaT3MgTu3goiSMYNQyMtDlil1tSRw4rLZuNbRxpQLJrNm
MtBnvny+BDu+ER/UdjRLeFF6Y5i0ikbs6xoyqcbbqWP7gQG7b+V6nEwxwW78t9tjJX+CHlMdF1QJ
FAbber373WKv6AEAUJ6FjHODnaqTH41cU0fJHqkhOYBsaagxKXn2yai5Kz9MVxrCo8mk/7v81yUU
0YbMxzUARsdWSgC2hPx5s+mGIWVFJTYao9GvStIOFHC1BjWhN0akbWfyJcEzQHjKFkTDMbkTU8xt
wUpLLjrNyC9ZAfPPyBgcni0mwpckM23AEMDAXMpN1842smmPjCVOGf8W1aPMJjB9UtUaD6Ouviqf
Ml5q1K5LbwbaW8Ixmt/VF7PTLuy92hd+I4C6ZJtC3RQIfjOfdm0ps3Xh6Crt5+1qvLPVTe1p4Ozz
kt7y4kAS3QeG7WBUc1mdJA5j7VLp7N8SurPYoT+yrXsY0CUGRFXneHajOh2lg4o6g9L6mUjXHkhj
PG/7Hww2sJoQGDG7jRnQ06KFBbeKxvfWwbn1/gZ3jcjw/yRbf0YG+4pNRPHvSOYsZ3Ia6mKrgxdZ
icvlDCF7CgJF2LRflijS1rdD92o9oMttmo0i2+g21CId4t/0nHP7tOWd4DaUJ+s1WJnho924rTsX
TGEcH35OtOFKU+OhoOaASPlYO3gZ/tsdiK5aB86ZYsQ3RQjzZ9H75upzWXtESZdy3BE4cRmmqDGw
gWjU3LP6qd8mY7WAqevQ0W766Lfwf0gRGLT0v8dEf2OSf5TttHHRRCa5YBeKKwuA++jPMnJByE9G
hRvcrrzb0tdMc6gm4tYYn6INv6AshBgYt1Vp0y6D0kFjYg3zdvnF1v4F2+YQ2MtZ8jtK3m2O/IHl
faYz8XfWB4c9+3JUzOudhfDwHFzzUseuXSe+gW/hPBfnTmBsXzkiRdwNFJJ07UmXg+kj2DZGC4Ve
8nRVXUNSzJZhylDYLfmn4ui4NL/uZp4mZHP7D6WUGL2GteO7B2/YPIB+zb2cmliUNDNq1Syf14Av
s3tClIH2kehBCEa6Y7YJMRV5b2+IKPBRkY8fGj8tJEP8/oIYO8Od1xb/qyT6kW4ihIgjFmCCq6aa
xCJ3gXpIidNh0LECY5AJRMxafgGBf4kmCfiNdWnFXu80ak3x+h4wdFGAe6PLOz9kZL3f/yTP9vwy
F0iQ3hyglSDgb9Pog3sdmvbKE8XLp6enAlkMidQtueL7QFqTgZc0tz1InqVIvmIeKvKj0Z0B9gkB
RXhl37OZDdYBunGcOUIdpeq58j/a0XfBcxPtIlP+PMpsyvDFAGY0QqK6XqGpZ8RCAfPVnhZDOSu9
V7T40Lv0TDVY9woxGoEVFXEtWAcE6Y5NwghQSZUbMvDhWCP2SJHP+Yv4L5KG+7cWR0DLUomzMqYb
HlTIZsk3CYDg6ZcQUIIo49SHLhX/48w7HK9F/KvnjLwrIATUUJeuzw1MOVWf9pmiWt8NPgEEnU37
VLZKjdNJAZiKpR6Y4tEwbReDyjn5/rY9h7/Ax5lOrnItu1jG41438i5X5JrZD9QNjhqvIXUHrDbT
Ygb+Zit/UIaBd6x+jo+3R0SL26ME2CyFOn2BjlID4FBsY9jorLhA0KxMD+zwNa0nK++/ba3d1E01
vPvOq3yb0eXovozBJHyVmIaTj64sdoensEbjy72R5MTqowgtX6wtwcyeDnT+bSi7yohxTEwZaAJF
yuQM2NgLjKrXEScb/bSqUxtCmHIzOo7SNkeeZo0KlRiL1qHJtsWLnflC9WempDWeDeqvg/cCPQ7p
ROgP7Vs+v5E3AsGK8SQob9JEzzn0P2LksharCms3K4ahkgynqKM37rKhKjPoM5Az7ARVk9MKS1O5
ka9K2SyYfjLSu3SGq1uvjJZE15KmkLNFyz4DlZWkj88JVnekoAtrf70/ni5ZPPqsAlB6Ym38A3kC
mQpEUefxz/wY0K+wCzxocVZ5dinzUcB2DSGkZ/6p0Guqd812sct1VHkxeh+uxtkjbBX/6cHA3vll
jbHeHVzO62rvW8MuRQ2WyK7BVIlQK6O0gEfaaeVi975x7WtX0CciSJJK/lb1B8qcN3h8iL920kTm
+/7X9B7VUcJHv/faXxKFcedNMYrU3zmQ3LP2JHR7fAeuZb1SmR5aNDvzxXvEltMDLmucx7A6TYhb
l422+viPkUhc3J88EZ/wYcEzv5oRnaoM8mHUWYfPh2LrS1lBJRVktZ7hc4Yj8WWnxVEskkE1nfzf
/Ibkd2DOzvcHDIDKryRJoWrHmryQW5g3tNEPkmKePOfyB55wb4fGR1Bmp/gFyIWmrm9RaahPz8Aj
NL7MQhNqu56veOAahaaXxbl3+hcx47J8KOEvpWmWVwDRaXqvqBpW8N2aFHn4T65jmycoEz5Xzzhd
hfHpCO435XBJumVTSgQMhEhbvilWAT7agAsVs3PN/oGPNwN05yNAzdgyZtVwEKKzS8AG3vLb8Rvk
klHGNWJp9EoFLmuoqBYlB1YVPMVpQo2q8IJoMnY1xwTj4p5gfA0LJCVn3dudcM591IOm1wONXHVu
1F3jHmMY+AjE+RO0R37rBi+yzOoKMCCUZVIsJa9X0qvQGmgAROxv6kKV3j4iCuYu8glwxtKWM/VF
1gVzE1ZsOO76hk38/v443yqg6IStJRVZzmz8RZlIdM6246xv4y7gWaZj9G3Ypszbr+IafT+raubd
1XC6Yrh77sa29R6DEy0pb8rdKXb3G/nvTLns0ZVC+EpLzdHFhghrHS3wSKhiXXdMcRiVdtT8CMyn
nWJ4HyfgyyB1NHWy4eL4kdz0gC1EdjByClNsdINZqO5BSWkbzzO0MW0SXY9C5WF1MR1KjaBmiTiq
AVmOIemQ6E3Xo+k9F8XSqHAbGFCMavk8uqlYt99KzJCYbA/Uy20c6xpGiS4BIpDxqlQlfqD7MfcL
x1R8kLouBo91b0pK8EG4UkO2mWOpMjOQ+c9kbr1urXqKuCVhI2xLefcPkwebT7DXVbJHDh3iSvny
oL7L4E38fYSp9XHaanQS7x/mGW3JXMPGHQPZI9zInNh78bcZ+HC/nwO1N034+UC/zek9182+Nkri
A6K0ClKNRZ4rO1CQ86V9xRgc4gXqVqgoBF/X82xFk4Dkm1AcotezhseLctHJKnVYS7ETYcfJ1DCG
7q+B7f24KQSPM9b0eMFaWKVl2+WQO09i7apaLjldaK3XuYRoYn29KVzY5NjETlvYbgE3Bunp0O5e
6jELlj76DZrmu4NWzqpW4+uy21u7NfEEYV2QAJSmZ8IeYmelICfHznVLbeKydc+RMBk6nLsWdHr9
UhunQhNBJlsICmDvDe2rv4aQVhh6DWnHMhTjnWoYmpk2+yimD2KNC785yTNf41CH2LXdEg972kLy
Pf7uwSiz4DsIOQ7Oa5UzsaypIBxInftL/HJu8wJsYO1htp5qv2tvDm/o2E9elvgjOKNgnyUxhXRr
xnGHizNSz+FN1Gn9aqx1xSbUrAphKG/kJy5khnhyMZ+IRqJWkLBJI7OMZ0A6+HvXZPCtA87GB4ZQ
ZGwXZYQPJsUq2UhvzX72qNZvFe/kN+tWtMOGv5GpEzNn1JWXR+rcdwWoc6ow5TuCgcicF6ALlb06
zU6TSOnMi3qW06nyBJsSfK6IpTmGZfUDf1uNDTAtqXXzwbeGqEC6jEo7YN3j1Cbgv6I9tTq1qgfO
xJCZzDWzmE4/OtmFpPpC3ID/UOcS5DlDvtkMVUIw9ApiEGIuv8/t4wg2zOn1hZbE8Vd+KkJO1zbf
8/8Xg3nTX14rXqgIjQQ5BZYjV8eK2DEmX4EEqCs2rE/dEN7My9w65ITLbanKIsI5xPvW/6EI4BDU
zBrYrIllBlnGuXxo+D7RB/XU+xGzLx6eooo/8GCh5TQ4igDFCNIFt0sffZENSl8e7uh4jqY5te3r
LZAF+Rx2+pznY9yfjvcs/Su4MlgVKLjOURaKdXV/FMBcPvmyWTnCUMNzTocaoXY19d7wb8AtQJTy
0DfywAI6vEwgVjii01SqjV/cXrSoc0UWtYNV9qfIhblWO3rn5tfOJhDXAkTcQ0XQKEiEOJ+12sii
CZRyN7SBOpnCgvPna6MDdNaekGzdp4Bfyr7ihgkPGFAHkrMbAzIzkO9DO9tzac42cahH3WrDh0Gm
U+nuBcjPJ6lvv9ietDbNG0SA6ZJEsaSXZ3qwlCSWraWItkJMlOg8qeKyNaheexQBs0Wu32CDoL5V
HYJqr5AsFUmOV/7jqQxp8DKFdXMolkJMxZ/I6yWonIxvdgQ7BSWNJsJlXiVGOU479jI7cBYs7YJ+
8m7MP1maTqnWtGWCOT2verdMFD9xIVqpSwG8rWYLRAwsxziDEA7XG5QaKJfHjwAEwVcMugGCytkA
SGp9t6MQpgT9Cd2DB2ZR4hvkLXMVRts6m6UJjOzMtriRv17+iH8gaJCrHEOOCZju5OrfJgEqyJAV
7WxChl1bazpsrYO8s0z6guXXKqsSGne8OeQQU7nLCtNtPt0bAd/GAVA++mvOAxMqCbU4dW9ZIKHB
sPzbm81wAjeSnGwhgHwf4504GXbfAPXJd9QkimtdaN6RhxY4+hKffrnB4rrVFj7C5LPfhySywOoI
2iUYe7GELyyOVaTaH/EjVYtsiHPn2bUrLFbTVzwB52/m8vXkazOcEloUySJOYm0QdVgVPTRLlLVl
M6zOlYyhRLM9n2iKwXFwO9SI5yv5mbQ+6synjTdRxuZVbaaSWv1NbNSkQ59w48KQNh7vSTPCHDYW
hxpfhpfeRfreR/h9QHjVvjaM8DrA9+bbatu8jenaEwPIgskh60BUO/ylhx/47CJlCz31H+p7o3eM
3e239v0YyeevbX3Ag6KHuK/e1KFTtw3KY6vN0SDQb6QIUDqpNiiza4mAE2fEIY+hDWyR1GM38RUR
kBwm9pspKCKwc448jsQ+Wf4oyZi9KY/S0VlG251pzHO+URvX3kQBz4gKRYyTZffxxH7f953IiiHq
uN14jk3TWmo5pSpoNd9tkJEilDRMNEBqYdamS8rtp20i591o+9zOheZP9ht0dl8+z2C2tGqiZoxO
Mtw1kLhUCmHQwzrYS3Devoh/I/DFhaasdDExlV2861jhHa5ab4PcMWyB2bzvK1xuty3yNJGYEJVv
ksY0hKOUoMtfEjyGoxxewBoGuVGQB5NMlCdLVNsfLMZedl5UHVAMibHchE+RaMNmc7rLy1y9gKuk
0NtrMKL0MF9F8Pqjys/gPoP+CcgzckcfsLBFar1lD20ooV2CBwvVXhzDvhAXZLuo0nHGBVm/iwzH
PgRO6bP2Z8Qv+G2bZAR9TuNbWhMjZphNOuZKuvCy8CxE4v/+JSM5WxTGb5YExMB0XMzGr2WIKpqJ
7VKFRhpK/Fy+MCkPMgDizVgs/qEMdPgsGOO/X9GmhTeUr+8z9eK5uKERqcBvn/OJkMD94Dpwm8YY
MPwj9Vnmr3uTGvztsrgsu52v+af3Eu0GW9tpC9+GiTFn52sFZEOQkQmrBovhWXDCdgjIQfQMp4nR
zKmF7ehvyyLFV+6cceGiLxsxn6vSxSOCsfovOLBLcfKFv10Vhk2t3qUwu0Y4WDOqBjxdBXYM5+R5
m0mH3FFkd9KOPANwfHW5zF+aCDbcMfiEOo6/aeE9Qv7e6Z+W83qKyFWFSYgIqXvHG5LA5WcoH1yV
/3jpOUL9KRNGGhBsW9FzMb1ddzdzxXV7DmEhpusV0cYvQcHAMP8GwDUqc25wsx//qYk5lURfxtNj
3c1g2FZ+sYEbqEihP0EzB0Et/XyjhDaPIzqprJXL/gvf3gs0yuUKI+w6mC9rb9HC/o0McxjxeHwJ
skHn+HwczLqsvKrZ6tta1z4bVFVG7nZssDqIZB/Opz+aLN4JYArTW114NfNPeSTMhDCq+Dpu+Tgd
SzX4CkkH0438h/aq8WTqp/SMbwQH/cuUXAyvnD6gOXxMPZ6KD+B9Z75C1qP6/+7udsXSJectty8p
SUCVqIYwUAdVEw70q2JPv4df3VsXtx2/fKhOqeXBFFon3keEcI8fYvhazhTsmYgoZnESl8Ywmot0
BcIRVwRKt15/w3s1xRVgLuXe2PpiVZ6POltkPAGu2Evdl3rH3ushFauJ5uKf2fM82c5UBmbP9Wl6
+wrFthwck+qRXv3ya4eJ90YUo3NImGGpL8p4TUDNinOiEzPQ2TDOKfxrFNQe+KABes9H4RpRmNXk
9gpEbJMK4o4A3cqZOF6ox/VEFWBITiFm9Pv/56UVu2VaOvSLqrD+IOpqbAu39Pphkoge+WjYOfQx
pHs3HpCPw4WY4oMXRJNHZ0pxkxWxH4h4TqxIvWxov3rXg2CwKvH/SCYVRo3wcZwZ6q5BLAGesWZN
hpMWd52jlb9bWY2FBFWdwqTAl3gYem5sVLWpiJZkEPt+2Qx+cJ5pJ9H0YvXTiLGq/sTh7WlrfSue
an1b4IhreCxDbOEBpFcf7Gc2s4Jvg6mFmkNwN9TCz2ldK3TBOsSCOkhSZJ9Ww4dqgd/sPAfBWNrh
o0ulKG1w9XYJUlp740NYyIlIEIcZtS9o7VjIQZQYtkOStJWbPXBgc2xskG4U9iftBNt+NSu+5bCu
pgAKCQkoRcCRunKmtFD+fPVMMC65630sWDYR4FWgUrPT6uZyV9IUJ/NANggkKPOEc9A/sfrNH8rK
LVlzWbv7Ys5D8h71mOVXPDkZ9C5e3Hsp+MUMPCB7Xgwv30BT9hoa5c/O9+hVnXqRvqP7bJ5lRhnj
4VS5iOxNPgv/V94VoW1Qk22K/6MYjaWmwp8Yj5rcMXR39yXuYvp8iGWW39b2e9rfTl9ng6SPX9LO
ls5QSrZMRTQ6eK3PqjFYERu5X1SzhKxvnTYAsp2TtVgyWkCQRMXwpEL/0K8zl64LwI63Yi2nN+lZ
U1/dHZ2UiSI9d19VRNXy4xUZn7LvVzwRB6FzgDuoELUh1RhMNZ7q0sMlY4qMbEa3RewMOx6I6VRF
TK0n7ShQXMCqx5gp9lW6A5pjsUYtW5JZT7cgIw3eSMgMkea5vwAHtTQA8JhhTq6M3wlQXr4qZ0Up
AMApE+sYha6IFPhBoJPcyabidnrhfbccb4mnP6y/eVDuNWDOeLZ2+Fbuq+ZWH8LaAv7x3WSABExJ
n/38P85Z5Dg6db+ibAUVCIWCRmVad1wjvzjtrWVGk0RXbDXiyNXjwTwvKHBs6j19WUbyDdz+Aj7m
Nk0kqKrrrkyONgw9Xvhcv3nWKPUu6idIOiPD/z271/9IqP498PcBbMfGvThPorn+mrhn5lxTOXnI
if4EGWaTGXRUZGfUvkT3fcUcJDI+mx5eWK4icVURbas7JeKZOBPaQObXLWxyECsBuVzSn+V8G25m
H4POv06XCTSEA63M5CJYmrHEgjTLHG9MvBzTkOhh5ps5kFo3ChGbLkcnMykMB75WleeODHEVqbGF
AO3WC0vJ9NeLAkozoi5CnByiNKlehyYdudhFnwsDHPr/5YxYwSHqHvmRq8LBChegqCK+Plwuv78p
r4xr0oGHYoBgwm2M6glTD3Qqk5ak2N+q3pGVgOf7itzZHra+OPlweqQjwMHYNNax7AFW++fFBbsH
NQ+lZkng+SQqwkc4picGOxebUMUZ8I9t7RJJFGaeO6ThK8T3jYO+Zl0jPzlHnxd3DsPY50NjVs7+
2Qe9MTyvo6ce2oPg7orwDkr1KnJDiIjbswh7IOemrq+idJzbKURMue5LhDKhRFvP3QpoeQPCxNHF
DPJB4WkQiPs1LY793YJXgCXg6DlOZVI87rwxNRGcJayqh+iSQ8Tb+XPzlF4mgwI3HP0H5PZjxVuA
uopEEib/fUgINdHEBy7PZIYbIgIKyU5LQWG6mkHsvz1W0+Wxb+6K0OsKI+/oqKGAhBesJvLB9W8W
69eRJBytq0NGh4Hf2emQ4BdqbEe0VAjqqrpUwtZDIgGbhlCHE2IwzZxrik0bidFj/YB5elyXXb6y
Kw6DUE1E+qD8CVeDbfjO9EWjJQQ8/DCp7Wsn9uBZIHMFXmRkHNtjmYA6HFFjfXQzm0Fx/LL2AZ6Y
ytp/eWZV1TZxiv+YI128kPu21MWWIhXI0WE2eU5IbvqffpUoxXCSuqEB7R7DYdd/udbyRPvQJnEO
YBPWNAlYgDAP2SvHW4x5mbawAU5+5gKrxA/jIfbk3v5kMz+qL433zwK8EtRkuHN7mhhoyl68H9/X
lVL3OEcsJafetzQgPd/odE/OsL6akk+WdOE1Q6ktHIzZ73IZv2DfVgfook+RF2p4uTcaA3pypISB
sZoxguOUGLnRYIJCwxrnobolaJjoMRqafGlj2Fba4IQ6T5KPAauL1nDYVqtXWGZkFX5s9vAsYkpp
ewvRM4QjDk+9jkNfI1tHHFN3n1QcTQqZ0MkixFY9EGcJF1LffNeC+tKIt8RoRBdM24SODYS1prjy
ahQpgyqtEfxQJkjwCbF5PcfwmyrV4P3eAAqV4yuGz5NZ4NnheeHthMr8/s0mNpwXfA7rzPODoTf2
+dARSyyzf7GicdZaPt4uzHwWdmUp1A+z4pOmTqJz+hHPy8tL1KHWllyNU2lodAW6rpmaVe7noKql
YFuKfqrCrK5v+KGc1eZ6Yf8j24L+VweRlwVAtqs1V955Ycpr6E+mm+Ce3dPH07PpKPKKLKH5CuEM
BPGOIy1CWJNdy70XxD6ABr7DZnfqlZSI1lrhkPik0p5iOSsaJFk62LJSlXc7Sla19aMcepW0J5l9
ObsiuihLpbmpbk4WbqYxIf3oD78i8BM+59QlVmm3VMksicXMj0MvIZGS/NymCyOhMa5Y80KZlc8+
itkesxpvpKARIr/l/2L1uXEVHA19qXhvMqaHl9wE0djIEgfsI9c69FeZV6YFL/qww4aOMcXLn3OJ
QqzWVJdNXZffmkJTD/S0zIVghmalm1jP9BSvKz9pJIuWAGNZ5Po1MSkrSEa5fW+/B4V79ITlwMgG
B+T5bav2Gc0830xjdPDwsbXwhEvGbaXKlMvT8vzbMA0+FxFxE4vTkkOS77ktD62p9y56TyByV8qd
8oyT3mDI4+sd/5iQe+bdz1me4n7hdfyVIIK4mV2ri4tyLW2OfL2BaUULg+0Xou4Qab5AcVEV1OVd
Ykeo5lNfrnOZcn9miArwVV5IvNqVVH/rmF7vPM5NHW22v+/MwX2wY8XMIJ+UxdivMtu43g6myVYH
caZgmrNhYGOQcAL/EoRCotfa0Q1E/wIwMRT1+7JmZW59z02fPypcSx4Ug9mVoPJGPpkxZiFl32j8
YKc7cjFivnodHcDDiu/ZXQ32wL2tbp0DB/EOnNYOUjcfS/U4PY4Zu5OSCtIlx5Ba2E+7OifWxkAe
CwShzSo88ibbvZxr3mPwy5l2L1M3NjkVZrR8YcMzby+JdPu6a+HoSVIy72T115FkLMbHrspJLl7z
gclaCE7vRHe9W7PWKduL/KMCEmwa4Ao4q8UY+D6iQtHbGPFDBDV06T9UisHrNjR8i7ujO84/+V4s
GQKfhcIy1s6bQHUD8GT949gxi+av0dcJaGRElgP3990sGcIXYIagFy4LRtDXlKNzN2nWqDbQD9Bk
HlITpFh/Sxb5MO07jzO9z6VpK3HP5iNKKb/o3UHptEZNjQuLedYutnteRYxGV4MxcwKBTTiu052S
GE2jaSZmx8Z9abW234kd25yPmlR623Njd4xVDk8riRNGes75DjwzOO65TM/EGJIURp7lSsxsEcws
0p76fp2PvfaiQsnsXac6ZjU7GiUD51goAM9TbhTW7ld5iGXfmZUmtaXh5MKWfBxq0kYEHAJJ7hyM
xxk5HORDva2xviHLcaLQ4BCTK1f4V1FYL/j5aMiEiqD/7ZHuNj8mGszfghzN5jiPs5nYyO6E39mN
hrwPl60mi1Spnk/d10eX+4/in3m/lO2GVvLHaclN4Sau6a22+M2OYnItj9rtSrn+uzsy8PMuH0Xv
WXBYTC7J+4N3eduwnUNXPmtOBPAFA7g2winrkcLA4MV9jsErS0mfq87ozy/X9j/osaQbxnZPCP80
gP0KhAnA8EEFfK42m1bzDO6GR+yikyEcGAxVW0dg1+ToJsnsMonovcgEDrhL/JbTfA7vOIpItPr+
uYauT8xrCVJU2iEN0dYGzXVGSpgMSsWs4vVj5NDjdQg7MWqj2lihuMQZWgZlCMByBaAclA43ZvqO
42meRMmslQXaO0B/5TAy9U2/uMaIGtfGS5ycWr1upby+V4iyMrnF4QgxZ+JlfZRxHyWP7dg2CyMf
cYIEmayeGIVK+zP1wlK8qZjiSWmBr7oDOU35ryaEECk1k4IHpPhcgmnTKPn2Z/WRN7zTvpIdU8qJ
pa+e7J98PyygZKXOLychdBOLSoWXeU6IN5R7bDofy+Ub0v7qZGYi4iwyU/hRVm/XsCaKRBrcFpKD
lXC9J6UQLVVoKJe6YKCpfsgREeh5HTb+85/Mx2OERD5g5aJJC0Un6LKni/8s9LM/dBlC9fDGmtpu
MlHBxoNUnKe4jlWelnGkEgEf/yDk55y1X8YikLycJP2GLjEDaXj45Fy3IFMV3pFCOqZX5ul/7ZAR
q1ZwF3BDJhJU+OsbK+LGdNXi4/CulB7Ng/Qpg/fZDu8IxB5IOv2xpXsXzxeX2BcMDtoC8y/tP3a0
OaO2w+fkT48y11FdumyGIWlYHJrWlc0lJ98lqf8WlItnS3Bewau2lrLCsj3RBzAeAK5m0bPorB3D
cHtCIgwkqjGShb26yMSdu9LHlxkLR3emfFYUbNZoS1lICtChG14HlwOtltsah6yumoJtfu2TOBZ+
y26lf9Teog1heQXnROdjp4MqUSZUymQ4C9MaTK5KQjFNXynYH1TF5Ej0frISl8Ui2rEjBiAdZjXB
NbdPcjEfGNBPZHaUcH3lIOhXL8INBSZliwb/1wmn8XHRV9X5CawBttjonl6hD+4MOg7nWUzwv8xk
YWhofB60Bbael9JTpGqBpCH+FDSjejcS5L3+rz9tzUvGj6drVHug7nzo7sKtaL1RbUrXiTrkf0wU
rYj6sagvd05jtnJJplCZmGFfC4V6megRyez3vFh4QZuQJC5rwRNS9GbKKIymeHJ8pEsNznu1J0ge
peas6cMy6ji7vYwncGaoB7PMbKzlMPAFsy+oWxJdyyNZHZPh/CQG/J404OxzPAEviyusR3DDarzh
mg3dTqxq2nKWy3gPe/U8id9aLAfwrg3CBr4hSS6KUA4o9pdP3/8uUuU424OPbv9ktT6R0HNJbdYi
hmQryBpmSiFTGKFcu0Mq6szUbOP+pSpUpPpBTj3n0S/lWUukP/emo62zLL7PDsakDNH+Go2Uw/x3
8rgnYnrBDSmvc2KIfTjj78K3MO/0LFLQAJD7Hj5zIZNVdd8w8CwPLXLlvub1cGpKnlvmnFXAJrJ0
iBhRihXAm08RyBmvW2D0qko+pcRhY20NyIalRdmKsBw5wnKgdhFZQjRxe0802Ww4DeY1t1BtYVno
7atUp9iMBNeOWCCFGzHkzaGsf7AtWHWfsr169747PtGorGld79H2iv98zVlY0LLwkrbT+2sfDHVk
qkeKpvbJMKYuofIEg/w51TOWaQrcYT1UCI6uDozMD3ZyIvVytLRRIISCekZvAhIGcUJzQXCDPzJx
A9Pho+U/DPX4COpRdHRn3WKaQe4+dyE1oFRygVWpOnEUsR1Vb3vpE+MAy4/+Y3DekjbZ/VKNGhk9
8Vw77VPdQa700lt2JEGlju8ONJMxY7aiuV14eRWttJTsuNflfPMRoi9suTKrNVU4wfIycUyUEXXM
wpRbZ8wR8AjoGaFcJQYWM6AdBmugwLKs6NWtIFn5WeJvefjEGE9k5IpANZ1OJO3077qpqkI8ce+3
Bq2RPOJkuVUfv92PMD4sJ4ekvHZcHfekalQ42evX+E5PiEZC52TdWRL20HL8CW1u3Qrw9AH/lJc2
wZwtsKyjV9LzzR+QgLIr/tn4zXsk75OJiehctxgqYm38rzunf2d8AIimU6z5LBcOngYO6JsuGbbn
9dwqCZte8O40N8jyOvstM0wln2vILKsN+4GWM+Q1nhpPCGjlU96envYQ64comfljdYlpQV7xuILS
HcA4aaA53l/tits5AgKkhxm3GsKXrVkYdZTGMcJfis5rgwo5lC3rRkKXZiq37Y9IZq4v+t68r3vJ
XrK/wNf1+z2gfU/at8rcjv6chrP+uFe4RdU6NwDgkqjnaYgPWL+F5nPJYfkNcWg/dYSzrApmTV+H
S00uSWiYNziw6E2wZXi8x84/EcQVGH5NLGRqBnqjb8sC7+qY5iZctDHzBKKfhQMQZVaExCta9ifq
suXCfia8rz/WHy91Cmv2QHM3rE7GNsBNj7+DjHa6Je7aayNhCBGHM6ZhfiWl0ej7L20woXdYTQJH
2ogqooaNlNQPYRZHq7XF4d7sNI+Qd+gT0J1Y47dIETG7vB7EnvXy1XtkyyjtoG7+rPCVaEqm79dQ
0Jsf+NlZ/rfPXmYdkS4jcJy9wgWVM3q/Ew7MGVwQdNH+d19TYQGcCVguANZeEgXoxreSggYsFgPr
sMqGNSXGP7+2OgcY7vckwBnHNgCaodOeWS8/jw9XQTqso6yJaIxMyaPc+UzTSpqsLxQVYvjxzO0e
DX2rl8d41AfH0/bo1jIRQmxo/lsCztC8UPVrQjpzIMvWi4a6ed/5pNjT5woKChW3fyaURI0+/LLt
itI5bMZIKikfhxfqZnUhXisYF+BVJHCjErTYFYm0ckXB2KiapkGE+gwhh0DG4+jmVgFEj12J6i7G
j+eMvgxcuE+sZchVmGOzPrUCIaPlwu4Eu2aAZTy+h5GxFBvNK2pqSxX76OU58+GcwfYxx8TkTK9D
ZSoERSV3liE2ltaDH07iGJWqi37M8orHp1TVONH3nCPQ6neXOHOu9bkQmaSuIkDe4Hv8K9efCvyb
GAtqhG4nVfU1ee72H6DY7iKnQHf0RmHA0WyqGR+v5wG7+htamPi7Ny0NVzxe8H6ua3UXZAeH75M6
fiWmDc43Y1HdDRmPNt6ZF3sHZzfUxXrp9UWANZDwc9zjQGwf76zVXkvxII3kfIMudWddVhHO9tfb
cqKOXFeP/7aTOuOUL8IBJTIuvGFfNNZThZpkHH7BkdaBoa2E1E4KPq9MkpvWx5EBRrpOtvQn8bML
UxK0scPaxL1yfhFKEo58ees5mC10iEl2PB+PP0y3e3scKlYBNuyqP5ltICKqVLPm60Iu32GwOm4E
YnJOWZheyaLQNbfGWEcXOLXOiwxcvzN8bpNA2JacKJ0eC43A1OQrNPAFsypHAccOkAl6TCaniCPF
obpXO2Gz527DpP8FPJ8rruvB/5N6zS1buotDhW+JDHa2yuPi9HpsPlvuCJNVJLzNx17E3bs/KI9Z
sTvv4xbQfSsvFSJxHq2chYqkflgVv2ugkzvXdgca8is7BdoyI0Qo98eU4WkBPnA4XtJO8N7G6yFA
b0R9WUnrvmutoVrFhfwk6IgXn8lUlC4TFeIXcx9t9lRx1y8pFMmPXRNISUS1ctYOYwPFUsPQTd+N
vzf3/fbvwRVmZ02W0BLrLelU+DulzgE4bqvUhQuFSoTTM3uuGJ/h6aVywmWci4ERy1Bectqub+mj
Ck5Ms2K8tH1KNpBUldVINF2Gx7jWniDnNdfUF2zBCGqzmxIaZY68yCyyiD+sAmmCTahj35x7ghAK
vqyPYAhwZvFkg12aAZHV6PUYFTb7wZQcOfqkA6FzOTNMn+ApucNOAX7GqCKr19l1HNDWfKz56KBW
jDfW5scsJGCTpnkS3L7yIIR91XqGyoY0FCbCCMyePMSaPJNFLAkQm0RitmYRmW3BtcHAeAjyiXdq
7YzfFxFuKx6MOgTv2OS6eJDi6aST53GxKj/nlE89Qw0/RV5Ss+WsJaodZL1CCOaN8TP229pPCIeE
03spxSBGiICsp9duVCfYN2tlNgRqweSGckUtWlnnU2/aooDaQQ+x6TbkWDhay64qq8Yie1RwEeqb
vopH4umDPQ+FHLeqdwmijsDQk7gyX5GB1+qSQSo6kjw9EnEnwMz2XKKifTeyIIhEpVycxHs6HuEM
L6RQYi+gzU84j1J9y3xWj9mkE7NqWuP2iJpbDVHbUPfyZz+oaPnxndWSuQNRY4KZ9ItefmwW8OsV
nI7SNGc8/8aaIuvx0JfAmYr2jo7hPQ7KrabNrp0fmDUoFFgSVGukuVNs57p0Oh80YvDHKlmAtS0E
C9lEQ7t5IIMMg16zBOutFvGp1NaiLPLtF8Vp7FvsvQYLJrbQbCikbUYAILIxIdgVVCcbF8sc4eCf
/5TYOkR0O/yaZM5hqJ/3C8zcTDhvaJa6u31lQJfnfS8tlqoYU7xvC6xT3Vd+Q88FSOQjIYTminUf
ISlIpWqRSfVYtUY7iItJk2DnAPqm8B8pDTif2kspQy4Odvn2ZEyzua50svf5JSgz7nqYg5qoVNk3
vvrm5FOrewOdowPol+FX7IxOzXPWUW6aWDF00mxcYHmTJxtNzTdFmuBrmvcaQVI7UpPPGe/tvVe3
flJSDPHb4jx68qni6Mj77OpPgCWYdCLLEfa4SK70I5nT1WSEofoPHNk0FjeCYXA1zFpbmbOowqll
46ciRSwVhVfCqU/UPCgY3ykOG2ZAIDc3Vg+FjokWU2uAouS48+qbEvOivc1jzDpXkIXjXX6y7FOU
Xgjuuko8XczbgbSEPhYSubHI98lwEbz83G0p8pWARtUh6vWBZvTtxVDeG41rxQLEh39kJ64niQlo
McpZrnmfnm4PDhkYVuT9Rb4f3CSD/3tp6jL1LFSzmAj0O5N8wWXXXEn7fmxnOv65zUELsSgngj6Y
0Au9FzG67DSfAfmgB1wjI9PJ6GMTh/Tlr4Z7Kv6nnD78je0JQzUh9/bVz+DQKPexMH77K62POigF
uI0rfAxs49SvEoeOEAjXvr0ouSD2wQodME7foOpAqCQQHcv9suFar/YCdpVYEhTybkqb9ZKRIOyC
jdZg5ujoZqtFeKu2pwHAhbPaCQ0wmhRu/4JUtCLDZTivqJQazCkoxmQ2UGuo1iEsyfOUPurwcxnv
nY5NuUDv2b22praq9qw5v35mx1NAWg4OZJuWfg3FhUxl+CLQT2YDftn9yGDY/eoyFCBa+UkLAJhI
8WeVOwov4TSXrWfr+/wJ0ek4uzu96svslVNhCn6Np7XaZ2V0199L6Vb2Uaa0mmAcHzRfFrSIGxgU
Oq47Yh1asv76g8/ICU0P+0u0I+MbbyuGs9JNfpsoLyGDatgfZQYtNYxRfQASZoNjoat45DVEd7yF
64UrSqP4Hn0qOZYg6LARWPrxdTH4XMZZBHMyTk8ME6bp7m2bUEf+jJGmdaa7T2l2oy8sMyK0dQND
30wn96UFw5BqSaj+IAFzOMF6snZzjGVFY4IhFtdE0yHGzzFAFXkCw4WuSrUPj/o9Yx08nhJATQmO
RlYvBUqEdyE6UqRBJt7wuRXtue7HDXjtxFCkiH9m34/92yi/BsmWys23gdK/llEt14jEgpAIjNMT
KW5MXumw+pBwtAMEis4xaXW/LG/9Gq0OeU5Ny+SiIw8QWpNYlcfh+KfYlLalgXJe1D8n3IXHY+W9
oNscStgDG70GSNZKFzXUlzmr34qogDJiFJghnTvhA3J4FAUJd3XoEaH+lJmuiXdPm+2rkq94J5kL
JdNXCyxEFN/Yf6fuKpI+Ra7Iwir0qRztJLZxIcPEVZYJfjSoUhzZ4WXMP8ORmkUuWjIVpIanEur2
5qPfUgZ6VZRQeOvWGHQ8hnGDXkxLkqsrnNnnDolOsRSfmlxnOG/C1eMvXA6NeP/eEwB3WJhJ+B0k
idrYm7C2nF8azS2nhPMgLSJSJHzR8s/0xG4UV0ubevi/wtPJ9mHBed1/WcVyR10xqpx4WpLkSdaB
dGF7g0jWjIhhwmVDG2SNOpXu5KHSB1Xbp3cf0Qt5JelWN5CSGSk+u6zz+zihp3UYwfBIlFM40WhS
w51TsD8yet6mmpmY8n+WsfEXqYIuYUWruKojrvyMfxMcPhzcAZoTa03jXMynSrlQI3SJ+Wl5zLi5
tpIpEXld+QBa1hlLh7l77KA3YRDApdGelPPo6UZaY/2uvpVQThakiJnvbYHGZBvFnszMjLh8E38g
p/v3zhzk+lwu8U0Jv4Z7zHVHkaoc1nlZRtqYOWhw+dFOawGRWIRHePT+ncBrCHeECPLcWS5KjWw8
M7OyAbdwnO8POxLXuyipZvwlJWrPvVFCzFm28HL00kBECbc2HA4K+ZR+sownA9BtGkQpCQpvbHGy
jf3TdXAmzmk+g0SlE8fe1vaZNuXmKKPeUCFAP5V9KCOzvFBMKtGvCcvB3fwlWFPrbC4UfSrPY3YD
3wyeR6kSDs0efsALYGWuRDUTy3VTHNgTSOZCzm5/S30epazpQahuUIXB2vaGpx2h63qhb/JdD8eM
WkfqmuhJPs05S/57YFLhsiaHP/4KAToR+ghcjF7RPBpYBut/SCttafip1QezKM0OGAaIbYVb/pnc
9diyoaOg9DbX/faWKWJaKmGa8bfDDrHEqIq2JVvEkEbVlvMHJt2AmfkyHJyhyTpWwbfeWww5y4HN
Z+b3LPXyFWtmwf+FnnySzOLAxbmMrbZJMrzKOJmwoeyj/ruJ2NBeyJhzqwvtYxKOOlGYOGy88xdd
28zHVyKBr66PHo2c4//pUgDjTjnJ5oetfDOhmsfgoQZeAZyJFMCw7ryuemb48ZbPXWnyeKeRsdDh
c3FzTabf638DUAV2PN0IoswnscmjUidyJwfLWU1EVClzuBuUqb5u+pzkPEp6G0qytVE5ndxj3bmM
vfu7GctmlwnN15dyT328vKgvejUtHRa5w5GgFYvsq2rOcLshuBHx5ritgnjQti2lhSpSxMD4Gi7e
M3j4150+8+g3ypEEZ3B4Q2dxu2UfugPBsOT45EuhAZEuq8vNELWsrOgSLeGwUP+7eh0YfbEC+0af
+XroVGWO2DN/LVcBc8RfAP2l9hYqS5mWSFF/8R22dimuST46s2x6i3+BlGZ+7FQRjJszSzJPbyDi
NxLUjnZI7R2NZbc3nqdgnP7oSKYKRHfqFfNJT5NRv6iEjOckvbNfkFADlzFC+Cmmr9KkejweiJ6O
Y3ubnlRsaSDPxj5twtaKt9D8o0f86YJ+L3l0cIMNf/Q6bB+s82Xgo6s57MGpkInputKpyo+NbADg
8IjPArWuzKLqNJJ97xUVz0Bx1uRSoG8wIcRrXKl8tX72CkTTGqYOFCZfXVeDgjy95nlpflEQ8hFt
U2DufL9Nj8ZoBRdfie6Ftn5kMhNLs56/42w3d8pn7vAQbfMcHUzYG5iybtxlmSaPM6yCw1R8gun2
+RcVTwJYDKWscmKTR2rZ6nAuHwcMaMeccO4YA0tr/hC67rLPeyxWhvwaai2szt159MmWxgo1aPXz
DivKQg21ZxRXREsS2fi0SCPO/RPkHa8SX76iJmWni3LmTXsgNjIiOdL0asxcmj92YmlIXiT0BtWW
7gOo7CKZnt7v6STrAohiUcZ43vSdrSSmRuOJGsHQicS6ZIRHYyZ8RRFpb3l4QIpGa5RoCkXGkePl
BK+emOAIwrOmXn19k3+/aWeqUR1tRCuuA2MloFz7t5r6fHZQ3HonwN05NUNUnzjQnMhhwrF5dHmx
6+my/55RbJCoPKt/+JyorOqOV0zxsxI7bg5E26GnL/oOzUoJpQ17FAtzP4+QSdydCl18Ko9HkLHp
BhNML5+0aGsbjasuyI3LxzGu5y6zmICNpib50keW3L1FBbrPq4Nm/3m6JVjdtQwheEu8IhVgmbmU
2wCs7oUO6vBPq8Yq7gXUNqYnYikaAP3HJO8uOp9RCKomxXJZ5U2z/ZWPA4sXyEelk/RzJsWm5kgs
nAQpOrqUCTqdLjR5mIuFfNk9SookOy1kYfGyOlX1EBXbfOj7aL2xv30o2/jns2YG0wQhNiZMSjsL
OIAaE0vjFd88tseXtb7DDQbAXR4lKkIoqAWnwszranZkV5bF9Rt9pWO6WfCNXocWu84tc07DSFch
sGzU4ZYycuyMaxrP3a4N+kpYYUQYJr5UAVqqzMtTIG8A5ArJegVHY/Qe4izATWaFHbqtFSiCo4Xz
fiPjN6/zO6mMBE44O/ziyb35Uan+EelsHJfrw6juAVHRWGGxmk/5OcrQeXm0Zhyqr6OkOxeH9285
3GrWMqI9GwdizzHOAwrEe4rvVb+yAt2i2dAgnPW8zcB42j9r1UzeynKohYRDk5bkNkc2v3XyidTi
eoyIahafaWCfHpg7dp6nm6OWjjT/1OVb/oO7cfPG5UTVrCh1lNjGgygBdM+11wN7zJl2trIComF6
EB1Ppan+vQ6MdYlBggnG+dZikMTMVlfQUUvFgo8CCDzT2s2c7Cds7/HVqcUQ5cDpiR+4RG/mcU5R
kUeA58EzI8IiMmbPZ0I+Dp0ozQNSwqZhed6eckHAlV6pabdA3UIbzAI35Otg5VXAaPwajWf01vvO
Y9C3L89P8VuhlgAILpn78OApFfOxH/irGEhyp7/UQNDTI2e2djxFQDHopFEdlActee6O7RaU6XxJ
zADOqOBVQCqk/8FoCOuYo8pWg2NiUNiaEstoXj2l9aSHVEEVeLfRPzWyTQ9swlLIKkaL2FMUJa8H
5r4jDz1IqnjVo4pPbh6tvEQk6BgROBShoEYZK5SR0y7CsfGsEi3rRUbd5BwJ1X+SMKT+ithGBsHG
zySfec+pHv30Tpx9fJmOCriRyYvXyRVsSX5kpfSTHIztm0mwvEw5aBbLZhMULnaeKCYu0pihpOVd
piA+n32ait3egwv9k/NTVBKJYd9TNdHN9LsNw8CqjexrbUmhLKxcDOBL9kQpQRurWG63knafQAmp
vwBa0bv3QcoPhfPRRCb/omj27+c4SS8+9eCFLXTEyVdj8tZG0stm03r0fogLBgsQJgpsU0II9C7q
PiRrhITpgHg6SWRLpw9Jjkq/+h5nBt+3rh+TlJuSo5xv+I9JJMM9vcwdJwIxlTMYH9UbCLL69mXa
qiDCIJBEKBUPy5FCVteQCbgpazYfXJsi4MbAnnia6CUYU8eXu2PPdUFX++FSndPY9L7wvprD/AaP
+Bw1q0CULRm52jVs4rldjsOY5FzpaMBkMuQZvUKNtSRuQI1Fg/66sIrwBBLh5qrFQvlGPbEn4xgU
jOpv67Kc+VNEnY7Nn7w+1o7RiSjitcwV8Ar2GMZj4uAUv+CdrsTY5yHRszv8Jog6kiplewecIEqL
XccloJpm2wIqSaI7wWe0BR6gi0G1ImFwqoejQom5n6uC05sHd5Mmr0tS9FOHGjJVHJFebzHp8TTg
4xPJa1jJx5bOtuxL6RYWSQdqF8D0HWtKOa5N97kYHpVdewinLRmfWL3VdWKlQdRXmoqUOcpYJ2um
BcJfq1xSE5xpY0ioey1qeVPq7iJnG7R5aHlPoAZpQ1Q643T7pk/eis8+i9ppbsPfMJOH2IQrWhej
YnrC464aggOt9QpYGP1ikDmWEPNKOb6j4Ls+k6khuzOm5t4TnsNHaKOOs+YWXyVGEgV4aM+9BIMe
Ctgj1jISKJ89n8eYrdm7sta4n3FUvrlgPb0vvDp4YZ8n7ylXrBbzzn+v8YpFwJz979xagojauBSK
t3QyKkexx9EIXbeJdmfO2Gj1hsFNtoosMsnU7G+1ox6s5d4bqcRjiNPRtaEgucrG7+U9VAV37EcM
sLk0zvu/GOUZdBQvsNgcGGPkTiXmLV6zJXtkcSNRGzPmpAeStjuZjdH5h4ffodiK/KuhpoIeqjdh
lE1lBW4nyNNuSpnF0D127s5P9jIKM079QA6JovIKccIwvGQ76JD+egT+AIXibtrTo1t0QtdL6qI4
X5gsVWCuxmR0SGqqowYXMjiv1EwfLSDAXfntGVjSpI+CK1x8WNFWpNurDM0B95bUAhauGFQW03lW
r70MXhwZjyLzRNr437qApmmshIu+ARrxYr6XIwlYX9kkPaKleU8NFgPYNGZq2JhpvzLgDjuQdpFC
/mjhOfhLMvSvTYuiFm7R6BojhceCJ2UV34piZju0VPLlk4/WR7On41F8nT1dJ9zI4txgX1tldVJV
/krT0OrSzzkI3LO9EK1j69S7lYm5Otjj/wZkCmBbG3Y3ZYf2Rsh0h2eR0xT1EVfGCZslHNeVz0kk
enFigKBPdIn09BHZU5sFp6T+Ie/vUw/IkHi595Xoi/U/FR+WZPMEhjiscrXPpXJMaqSZxtI5HPPL
tFqpVsbotHCYRk9X3323VV5qaQ7MzufJF0fwX0mIlAf5XwWlOv/4fk9V0t++PRbV3KtRD3gZD4WO
/pD5C4B9s8WQeOc2/koYn4pvCG6A8EOYOf5eUQEcQqsT7CELZbJcWPkmW7DxXHLMAbacRvlRj5Nl
4zrCmCD/zqf4KOK1BzLVWsgXaTL3OqfVeqwToNFXcdm53ZeunbEC3ZbjqnThYJUSGdPWUf2tFybf
5rXGvTSTlV/Rav5/BKVO/9g8p7whvz0Tx4IhbMRkjKyuj7fp7Oa88tszZ+4avrKC9K5Excoy453P
am0QQxyjLwXMnKJEE6iGx0/rAZfrrHKDIVkfaD7WnsOXbvgKcuo6Na86xPBi0LAY+tVzgZ3vLsY4
/rQXgq/oa/mrLXYU/gEY5+7W2VorpbJeUfja5b7LFN6x9eqjsa550rOfe5bK9+I1HoovwEOg/hJf
zElprflCblN0eOYlivsW3NofpCKNhWHEZF+lx5TSed7gSBLTEhYMvuFENkwuiS5Vy0syCpsgvk/s
gF4BGqX8nOd5neHtxDhz9iebEr/DmTBDOIT+yG+AeLFZW948wna8pp7sW38e4eNS3moCmOlEvUYl
nnhOV62ztAlKgvRKTH0d/whmDxIWYLDWxn6XICgWDf/UOaNx0PIgnA7PnLGZ6EbRdt4Oq6tZz/W/
5isUqftUxX+cKRwpVPr+OmHKvLd6SMGwTqDncEqDetvt+WjA5YFKyeULLNpUxJnbVFIC20qM5hj6
RdeU7KY9BNKDjZ9/jljI3h2p+Obf7pZW2BtxSAjbSENachLfcdLxcZzU50xfiHwgXLwlnwHz5uZP
29E/HIAC4K60uZG9UOjBNkuepHRHGk4+mj6DC4c+slcyGTrC/x9eUSQsRZz44LZ+S/RlP/ipuomH
eABrtp02ZF5+2DzpgRCxPyg+Plw851eTvdnwWSwQq8e0fJhOATKSQDuwjQZUpMLy/m/v4lXdq2T2
2A57yKBYqcS2bh3OiMlxljnRp8IT9ViiwVvXPvYx7d9pZBgoM0eFEycbWYiNk9xl1slNhglKCAmQ
wuuGXyqC8C6XzAxYwpe2nRIr46cdLH3t8WvHnd5dFB/Dr94JChwF90iRoIrmllXROAwopUTyQ6ZU
EpM4yvuXriGPAywXxQvS/V2yTKTsybWlyJMtbO+JggAsqF9WRQJYdQ0bqGggREDfAzxryPGXIq0k
aCsoizUgawxozh0Atz3UqIIurNwssOy2pBPAuX3JOnlt6iI9ytnHBwGY/nAryxT/KLnBm6vh8sq7
1X9U+2u5heF++1Pktb45lHY6Py9hk4+VHHkn3Th0JKGBHgUOIduIAv94nCooKdSeBiI7sHaGnCjh
cwU3VEbzmkfUlpUx5Nf0x5ZpIG3rkLv81uOe3Ox9eoZ7FAi/fP78WTiOel2Dd1DR1XsOBAfL/Ddx
N4xXK/BiMSwpSdz9UB4gNl/a4pFZpMBzEwubyqqq85fuIKMO3nlX5EHlsL3dvLPVCrBNDEGVbbpr
ouM5YVc8s08+uitNui4ejq+pjOdYXnv3lP1OjEX9PtiuQ/yZdIYG4Nh4EMQPiX3xRZiEhyEHWxx7
Brphv6zukm4Q4yQTvrwYwg66Q3nmLCWOpUEX0z58OfLTUCy0FVBNnc+J8IAo9B3NGjrUZKjzYXuP
K+sOgrblJK1bJOvP3/9ImbSSPCuBV98iQ5kIchdRpER9mz4Cqi7C8KnrO5hnI4KOmKbxOEo8VfAj
sEeHYcOBksUEjtvKP82owdMUsZD6PdLk0NnuwvgbYfVwOJg25RhwCJR/w5etEWGoLMlYJQpr3PHL
6fc41A4d2Uw4jCr1vsw0rWvsrIbHLppfn+otRclFjTKd3OY5lG7yu4kw/vdI8l2smAAK2T/cpFjZ
MgzsP4ZxohARyy6CjvpOKe74SE0yt8o27fyaWvNZ5ihqvi7D7Aq+7RA7dzdxTGeq7bQSOt3w+87y
swBDI5+Sqw8JMi3dTEmrj/PClZy5HzNJ39jz3UiJxqdMtFa+pC1TDdECgxK5l+s1xB7u4F22deIq
h0jD48X1U0E+4PycgHMe0z6RKTLKSsQkrVrT6/6QjC46ti+/1OMO7GUNfDzXJmkbsM2l9FcmchDO
eE597YmNMI4Od/XTVMSbgpBfXDZV/M4vki9oTaNm9UHm1dgnAO7AoxVvU6i45i6dbFpIGudX4HVd
g8dUOGdCQjnzXEzvUTyuHowd5E5uAFGBRnOR1gznWJzZ3KAr2WlB9bgIikG5d7lnQs2VB8ABhpbZ
Xq8AlaDPL3ywwDv8gNGxt94xkxCbhuUu39GqiSpOWX32z6lnXQLvUwAMpZbQTOLtIX/sgH92tZ8A
ELBqZxQ6tKiO2h+A21Wcsr5rDpFI76IouBWJNzCbNlSFhVuCWM3Iqy8GYsh3l57JS9Yf4xA1fegX
vRcQtp5kRGHaaeR6O2RCVw2cp50zN37TrTjUG4irgdLkKN93pQQcTVTC0F6EQiGj9O++tWoQTjpU
vd5ksghlyQYVDlNrAKY5twRCMYKOw87anoQd8JtFz5G6Nn6k1dSu1pwi+IGaxhccP1ipBg6TVXwz
hGr3NwqZBbtbjHk0zD1cGWqbG87DiIxqwwrYNaM8jGD7XZcp+CmHGTG/P/lIiRnd2cG7EJGyGt32
kvWRREzmhVFOcf9j2bBT6sWa8aRbIhjURoQRibDvsGG6c0Sv5POZw6pOPidDwoL27CXb1hCu/09g
EbKdRsfpeon8GSVyk55NJ/ekAw+BJMp4CcTPoaNIxGt+xHUyZvkYMNtSnRWlYuxrcnFoQGIb1/p8
aqDII+YmeTHzAtQvsbT40g6hOoK5Epp8xd9fSnCoMS2xuZWrMar73crJPXWpVIvOgFvVbf/TG900
Xrkl/AWSP9uasQ7JGMiReJ/qdKOZeDqcgXw/EkyWzqMYrRZ2vKKqYhZqCOG8F844vH/zrHkEczY2
pOVwyAwkJZUjz35DlCBO45tRBnGHIcZdSybHhtYdtTVN7Acae3Efbgp4sBNLdOVJToOKWQfgxviS
Pcr/C0SsGc+AzbfR7CitxChQA/ZOhU8plkI7XBzb+23TMoslYOyGdfDu2YxXEK7WBogL5s9FadVP
4gJcZ/5UHoX/btlLl7O1K+Ccksp8aeKC7WcqKDeY2Iv5HryXzXlp2WGhCm4K0H3r49R12GhgsKv3
1wC+Br5J2i6/qRxz66YEbGIspbXrotVv1bMOaht7agPVTY08AgKDrQzfc1ovFzYSippfyhzglV0Z
j+S7IB8w1GbBCxXV0FBXS4SkdIKCkS7JQKaJE73wKXsIbo2bDEXvd6QVaDxaQmRehb4V1qjjGnY2
EKq/kp4E0jDZFMaewHiWBfiUJZMsZwo9ujafvas4cpOz2TSMdRSyHRV/Bx3BxA6NMz/Kk+BwGjxi
umoogRFZTFtvB2DbhXS0mDK8JJDilViVxl9Ql+tF9fFWHKLeMIJV4ob/YuPuHUs8LUrcm1EypTSh
Gg9/N1guak6Qx7lwrmsQEWVl6EskCEi3z5r+gnbOYsCRt1MUc56U4ckuek/MZeDBCpEERT0tlTZ1
zc6ngtgThrdnSoWOWgEp43QSgwJKOPJowMSnB5IQFCPpLinWPa01ZR6j8zAHozR744mP3SS5ruLD
DSyxIPyLDv6Lf8ZLbyhqA6wbiYMQs5CF262ZbPTXTCDu8VG3MZufIb83KkV/2x0tFCebmFPMhzw+
OFikgu3AClaC2/zZTnM+23WYwcg7lfKmcqoPQbjptyql/8Q/YNvWRA6uULnPluZTANvfMy1v+4Rt
9L7s+XvGmV9hD0nKFx3Y+qXd5c0KcdOFTX62CF5qzZHRH2TLrr4ofv9Ot9mhQ98CkKN1HPa9TloW
3+MfvCPP7xb9/6lij2xHxLlN3+EGon5h+Edhd2hLbn5y4I0v80iYt4iQ7PsNZiZ1Cmx8MbdHkQTL
yXTFaLNOHIhposcefIBup5/vY7FtqslYe9nrudUXYzPgE6vCx8xf4nepkN9FDc0yDB3F8iYDUJl6
gmpnrKn0PbheMF2snF2xRR1QyxK8iiBz/DdjH9Tq0sQZmhPrhVaWoT/6wn0Dj1BOyU/CfHchRmRw
AdOY2W+JFGgP6Y42HMFu9QWMR4XEuJ1PkcgBkh0hDdbSPM+4MrO4LuDiDM+mR+B1+LXF7CgPv/Q9
9n6E3dYcUTQaFL0Aev/oHWSS9qe8JUmy8Gs9y9A1uLIE5IVAtbxZxiemPeVbJKAApkZxbMvr5YQg
Kuu1eIpR7y7+wWT545ZNSbevJUQNm81gIehM4sJq4dAXV7olN1dGlDb3dgcUX7IzUJRchpl3niJQ
LjjujpfcXqolLd7/O8dlm2HlZlFu3lLYWKo44jS4Q+C+xpeZzqZ+uxNxoYAn5jGmTrButfdVhUXm
/jr8op7NXY/Z+HlL6/a1fhlsxeDBhVuSfeseGOYp0k2k7rpeG00/cMQLNyfOMluG5f9OB1T2UAUm
shu0WfHFlNS2FM206lwxpVfSOnVjBJlSqWg+UmxhKaF1H8uOjZoO4Hx/Ua2WbYj9WahxpUdRS3F8
TDco0eZuQT/4oflOJB98yBNAKWnlL/uqsT+qESBklrLPsYWUoCIFlfGjSqwZvRkKl+crCa34faWS
IFW51hlwKTtaCjmRX9TUrWowk8tzgJhm1RyKomUCDY8neAQLAdi67ev2a2zOjUc3URxAjaa0fGkS
AjAWobKN1N8A/2JGkvIDZ/FjIcGDLqd2XsGxWU6eJw+xFoP5Hkb+qF38MW+X7lgv0X1vp64gAS+l
u33rE8lUa/0tCJgmj0zM7OGSBoOs6HOcrl/SYDpT6XDdJkjom5jTCpOUvvUhjtemIr/vuX6JKa5u
zK4qJnCG1mL0GiSzXBJNlkZDKYT8uGj74AE+8Ib+Ja1cVqex4tAnCPiD7vm75ZE9zuW2GY17YCRy
t+vkU/8Riqr9M9uGkSerV8YN8IJDuP9DbFVw7usOn0w3haqFuM78V6kiASmeLICQGoXii/VnVFsu
k7qIsVXwWhBYgSt1u7rF3Tf3vGBmB+ATlaByeIN+JgNbi3Ko03111gBYn9OeCvmNO+YYjNWY8WYg
M7BTfMylCelDTjG5SfKyJaavrA873HGla8f4AULyp4f6trXmwcThw45wLLmOyd6pplTCL2UO67XD
Luo7KADm2OnpiioTp9gtyyYYexbetF4DhZXIFV800zlS21oIlOvt+85242cfiTqEf5FlbLlApDWs
nD+tKXtZ1r+O4Tosrc9kq8UR5i1kvexEg+fudZFNuPSRnPJ8AKXcCSVghRDjpSBNjXpZ8rlmVr16
oB+181YvbggOnEGBmYU7rwnU0OHjirwI5kAgVEULHHTnzdFNp+8McoRIAhptAtHxw3DHMT8KHvXc
dhq7pFv/f59AH5/KC+IFaWTknE85Zs/Jl8rsyGSVr0ogrIAKHvHKOoV/jEPTefKqY/fWFzx93mZN
5YgnuEZnBPMgu8IlsT1Ofk0hXtkNO+eQFY1Gwn2b0ruCiHHYqcAbgPYIh2xKACRdTA0/AHeehIXh
KUirf4/L+p51fPm3DxnGLD+FxprAFR5JXKafxoxJq1iUY5wfOSPCQ4BlNocqPPmdgTNzdzBg0A2y
2RcHABmAxUxlI5wjxSzc/Luw53khkj36aOkWoL2nNh9ncmv+wi5pfSkxrUkSq9otCNE7dmnW8H2G
u4VAi2hUX1mdmAVtcp8lhc374AFCWRQICBr4LS7s2x1j79mIodwJF0BU7KncpeJ4RMsMxint04Yl
1ZSt02uzsVRZ2SmqrRWGsGsVewHYqwW/sA0fNXZ80QKZY6y8rLK1FZN65p3zG7LTRqvuk1KiXQwE
cUS6l9iwwNwArodwl+z7Dh64tC0YNlGgt6wc08pNFHYJE2NQbfkmJM/yw+jJWuCBoSZ9erB3YW39
ZSZQJztz6ueVGPLKugIL3dpcagp8Us7F4hq3+2ArDfAnsFZFw966Ti+Mn0OHonwoZpFPbsUY9jpT
bHG5dnWERV0JlEr5AZGnsmEvtJa259hGYJprj7PTD6Wf99NI36iAqX9vci7WYCVaVQXVofiuUlXB
47pQr2MEp/8CwDVSFDhcbrc/bD8uQ9tM52ElTABFLg1G4bE4RkOMgKXH2GJmg42wwVyRS9x7M5Py
H36aD8YNv3VTr3wLXg/I/rGDkkruAHWFTuH95mjWUF5JJMCrZ6ZPc7U+rboMRikFtuYY9AbGnLqx
AZnfg98y3vUcU1vhV0O/SgbZORUYhN2LfoZZqf0M03owELx7wnnGvMlFdcEu2oMGpZYk9K4ZocKg
zugerkJtovMNgk15mIuhzJ1nFSvXSMOROKCGq8MfLcnqbTLHUp2k2deyzfRQVCAPmpmZZwAhnIsv
OToRVYqi/Bo0IdEwrLCDsiwUy/Vy/Q5KetKDUSiwas9USJS+3aKZdD655NE1AwFqJL4YmsLdgocB
xneRwss25Oibjth6r41RJ5h/TjWrQbuN7d9bEzThY1aogxjXEl/LLtovDb5M/+7V0aaI+0HJcSu6
MOLosfJ95QkfncKJrUjfdnyKlXtoV5g1idN4qVvnGK1Ap8zv51Ifcdaa+vdViC7gltBXB/AmyYWO
AkYKGJ4fUTf91uLJ5pBodihig9I+NJdoRxcyC1nRfd1tQk2p+kGX7jgJA/VZwVj+369WYAyYE4zq
fGg5FgJ065Vl+1WqyuAJN9pvREBMU0CHt0nUXfy8V+Ec86k+7Zvo3GxD1cXjZIbcpY8e8BgQbl9y
XT6dvRX/NDRp4oVd7ZnbM87suY8pk69iou/soZ25azZQ72mCx6M5tdbVE3kbM1Go99WuDmRuzz8X
TWMXcEIwn4htzlXZx8/9ogl13I5St9doEi1XXXRDuWOsBccrUskniNdHnlE+p888hClQ0cGq8kjZ
n3TY6PLuRw72R6pHzKA5E4mSlzesW13T75ARmg+WWsNVNHjQ67hK0b48mYwl4QzaONBSuCa5jdxW
VklQZ+w6HMNi/+b4I/7ZFheXeV+faZ/B7umo7evGbBus40+nN253MHwJ4220yKI2+ebNNY3/ID3W
u/meCbJNmUuwNe/X5GMEK2fXM5sJmtmSQIa6nsQtHOQi5+5Ee7vmWQvWoWMpUf6jO9d5A0zKWjTe
Yqvx1XQbOA3YliAB53jMG4UNSjVC7C0Ubhu1qqKdFddQZEXP0fx5GiJvhiWL+ooNQTg6jvY+GuK7
BTD9oSzqF9XDPv3k5i1StBME24VXmNRqUgShyzrWOCy/5BFQ0YRwxNhNmzvw9LqAISpp6xeo7ZlQ
+prmdJTU27dGNujqHI1vZoNmcfx5LOKGK7gJ1Js6zPXKUWbjwzMAU12KE5CGWUhOB+QAh2oZ5wJw
N0wr7HbtwSovQoXX7zO2CNiZhiakxEV8hUdKrINHQX+VrovTWIvlfRB1pidvh3aot6NNjUYd6jQ5
yAu0EFGJdH0s8sTNbPY4H3PJ4sjSt9U/Fj5nfjimB6oradUn07/9sRM4y+L92CxqYQ94WDNmbZYP
DTVpeT54OTDtjzy2fAcL5y19GiY1EepoXjkI1fdWDY9ZJ04kTYdLQn4V294Q3Eilde16pl1T9YCp
Xj61oOtnbYYfrdfI1rwy0bS3JllPxciKm6bOanaFJ3VzSBfyua628ehZ1QTZSj/f2IpKbFrhy57/
T4cyZ8QPUiO/JosJpxnF2vMgtM4yuWPy2oasj5gSq5JNPhp199Vp2iZYTtFZtRifbrfMrc616RaA
KYzdaYjGaHjfvU/caaf3u4zuGPunXrNJgb472yCn568PDhJofB4DqrXJrit6lgT92bRKcQ6VdYFj
x2uUnYz46ymfDZ0jqDJ02rI1EXSoGB2t4NRtwt4G3yynu7/Cl89Xbi/TENYkZ9/Q//rkktNUS0LX
Wh84xmerMoLF8hp8sVD9DLBFeyl7CpNsuYC9GvBjkCaUmCpFt77OCGuQxFfFT7Q34ctojxvQsc5F
yJ700t/tNEM3uW7cMxlmSfmpOgbseZhW3idJnpS3W872z950SLwUPmEoSmbBTVF5rSTkLcb7woUH
7nIApE0wF3hco0wFWmszwC0lr3ZfgTK2JgbAFuytUGz3K9C12G1FT0Msxm7jnmDBpQOp8uvzGzy5
6C1lRNj7sEzFbtZa821cljE0nzg7DmUnd2Par1l1Ydx7MpP/dkQhvvq80MdZN9zf4Ju6p4/GAQwT
jXRCLqX1ICE7DtSiwie3lZ2oyvs54chOgRQ2UiuvycKp1R249xaoLGm7Q0+54cIb8yCJuv3NDPqe
yd7OjPe7vLZZcS2XYmZFXmjUH1QUdltNx6+xSvk/+aWzyrIz1XHLio17F6tYHERHxqB4zzIQxo25
wgO/640SUJeX93BBo30+t17D6qbgc89+V7BwnnzjMCAw0msjs0dy6FzLE01aN1RzmQr9tGjWZ27f
yu1+AC0GbSl5t75zdHW2guxhtk3uRejegHOUs3LE+wSS5cJQVaUYCA3OvIsYpZ/5Fi82sW+vKwJ3
m/dehBKN9005MEhqoE/T1IiSifCd3KqZcA1kyGqaoxDu4JEjP/wt9SBbWV9tFuuD/Sm2edxiaZWH
4GoqSvvxIVrtWK0MtIWNYS40r0QUNSVZrSI4IuQOuX3t2k24GuOTB+t4xZii5KZAQ8JI1/ZjeeVV
2DMiTS5Sz8P7kJTIEiiHZWMWnxaVzAcQg58iUUObNdOaZVIfSXnSn6/dMaW0gPMWuKWE3xEfSKeW
xJOE3YBP6y2kqZ9TNMB6oiqwReqdDvXEJ4TPTn7WmxfS8FJTUEoi2wI9eI9wisi+2NO3H7AuHXQ0
T03gVFk8LfRbEpIo0hcqaarOwHZcbgMKvUEB/fAl3R05K6Xfhmvj0mrHuukM+K43qLtvxn0WmkWY
QJHfjy6QDO2Z3ScMvsS3ErYLdTmC7ToJgysSOM8UUucIt/j9TQ92dicQp5UvJvADKedfNS4J7Bgn
xXll8gexfSAm/bv4wewlzpTLrER3oo/jWV7ZQW2TZm3V4wnMhTaAw3mKsu/PRMmW/IcHZSxl8d81
ttvhL8TaAlDswUzgxoqyc0WY/T38DaWzJ3mjaFHTz+n0+Ufus3/E8Yz1/YkybnIFN93xZIWnd6VG
b+XFEEGaU44Zj8A5rxnqbboGKGLRhKes8MSVUpn8f6/fWa1iV9krG9hV1zIy5u1HtIf9o5M+9JCv
oqibClzSdraNdEBuML7wmVUqTkdz1bx7RplYoh2yyBZjVVTa9kNIQxHtLwUgerFD4bRA953aNxrQ
0FPZM89+HtfsZnQzABk8BMaaAQzHRg6DMv6jykA13WybHWvI8GAX15VOqdRx51SengOOnUEmnPGM
wBsCX1u6ABVDed8PKC2YGoRqsk5BHEoq9sdTtW7WNh7ZT28jv2XKw1AbvpIAVfUyl+2FvWtuTk+S
8o0WsaeNbWtBYH7YK5xo6EIZ33YPyvFudBu9ZEYB3lBVsYriDvqtNMWH2ZHwNxtmlw0QHx+RIeMs
H1oSElL+g2E2135+XD2FSBRWf12aokpB3Mhj6PAFc03MUJxmi7D9ETrKRj1qINZjqG8gDTzdXlcy
YhLkleoAbG6Wk0pDjH1Qae3eRT37/ugXZWc2VSWE+AVzOoat/yE0P5/WazyakezTw6MXoShmP6py
9odC94SLDs4pCAz337LWucRTZsceaphfIjJNXj7p2GQ3WXOS8WDjhkI1CLtm8EEDTlbybbbcs/y1
h6zGkgWK0PubS7r2vtj4L4lIb2o+Fu8arelErY6mAh8dAgMvNKsBum2byRbORWuqUG0UPGyQbCyl
OsjNrJ9QFKqfyQxz0Luni/gStCnUrP2Syxf/4WNth4H9e8C6vzDuugzVV8T2Xev2HJy3SUemcA42
t3A39PYTb7Sz1U3b7TAj27kf3uHiG5S18c1pcRjnTTa3L0/34sw4grz8Fgvmh0gKChOZnbuYjJvz
4rmmNhw6GEMtBxnMDF0nI7il2vVcBDllGmdkqGJcVMgaIHG/sATKwUNNCHwZJWiUQgA/p80tEe2V
RKNQe1fceR72CjjY2qRaIDe0FYAe8/2jcKpkjy8iKlP0B95euXmpE6Zs+rtoWbBVS/hUDEckX3Kv
ZIzKkdCsqJ80lRwHlRhrbgiNS4o3UKD/TV9Q6B0ioMcHyV9I+YX2DtFMQj8/gPvc2jermFjgmsif
8lVAFst0TEP1yZPPu8hYl5uzDJODH1hoVp/WxuK2vMG/wF1Nvj6eCZ855cR/C9dgQT+ugk7ICUOe
A3Z9ZZEtDg4frT1oHT2HxWItPtmyMKGSQy2AHQexdm9oVqGIylB7Bcpe/I4c7dMrsYGgN1AMJlPh
wxyrzIX2jP2H9PZfyDQaJb7bXH2yuin9yeZgeZ11+B1yji5Xoy3AxPV+qbypWAuqUiBTVWE5wBZC
FImHIgXNcdQU/MSesLZkEOGIpG+qcibJkI+OeWfNi/rIF9LG8HDRbM4SynbF+NFlw2nruEdy+BdY
Y1CS59c3RNzVOTQFsrwXZpEY6NLgkhkOr+PqP6N+vlpHUIo9eXh+7PJcway6zB6vOJr2sTXLMa97
SFBlXfilYJuhYMfGRxDd0jiDEXUk8PPsFxacLi6e5GjGQbvdpy2o/gu7/rwJ58J+gA6iEdc7HY7V
RjzPcR4b9NfsGe3y9zhT9W06+9NV061Gu/wLtLBZPREKzq1CmB9mLG/mIelikFa/FjFRoZhjBIXz
uaQX3QS1RAzrGYdrCZvGLS/Szn4BiGAoAjIl9VmDml8h9bhcYow7Xx2zqP2PSniwqb/dVzPoGzWC
+9lqXTZVqYxWRxrOmaM9UKXdvQ5n7adPzYkM15ZyqG0pmJ21+91nPVwEc84ta1herns8cRxe+Ry5
vb5RyPQKr1AxKFgLIPio27GY9TTMPiObK8logDskNSDzog7FfbC6C4NcGtbG2M5Qadxn3pMBTykR
J/Iv68IpaOaLqzHS6cNaaBgXM/iNAxOVjbd1bX8xvD9ZTO4lnxYcFeLdIYgAOatsIaKjDRj+S53U
n/WqBXF8gAKYsj7t1FWNc1BouZSmAWtbcdJ6Sb9d/brEkExq1Dh17GzKrUTvku3WCrPKGRNzso0+
irSgUzY2IScHXQbsYXO2Ke7/ftWV2PYsWQnceHzlOLSiwOLS9L+DwzkWrwHn7sRPuSm4yIuCkp9E
khMAIX1xRVmZQrvK5ldi7BLOjP8m65yiAuaTFHmXw/iqTTyxEaqSxa7dfyH0Hg3kQLwykH/kc6NA
+30IwTeDne9qc3qQEKAPSLmmrZCPN6/9SOYa4FLzCgRSvuZMJMgrtWjiEbtuDw+JI8FanAqrHotB
ILRusBC/UNvA2NQO90L2T61gg5nHIlH/R28DVKpGruwuSrTPm8V5wtojcnwuAf4zs+PSIirQKrxb
y58urY/g0Np7Xo9GIcuor10a+lJUF1/OqlO2xKmi70AZaW4PtVCBfD4u9csIN3odHhwpiqNXStwC
9mn1FGbpa38kn9cqWWS3htttW/PmRhTxri5VPJvN1TN2Ow3omWik8npUeuAYiyTaMAtZbekRST2s
M/c1x6Wup13n3fOzx/ax+0yrkZWqDVsf6O+of9nnwfJgaHWE9uJ74rrt0KM/a6he4yRJ7pl2JOqI
SU2ei7vdoZDC84ibsR9v/yxmfZsMFTB9U4g41oSP6VNncElZXWhwnMtePmkViZE8wlYSafqqG07S
6Ed4BEHt3jZEGrtIAUSq1gZlNgzsZTrwwwLo5sKv/n6mWMlvAc2t8rOlmc0VkQB7LqkjckBjbTq8
EBSzQnScwb/pIBy/FNRljoCSUEUm4d4e3efp0LR6m8VCE2YlojiNojY55GvQBOQp8VSOi6U4tUdV
32pl/457vgvUzXFMmswO71Sd11VWpJmr2+OL0jjfO3g9OommUYCxPiRUoFvnpr199NoizHHWRNse
TuCtyYVszySfgbt9l2TEGqdmqi3dzbvm49l3TuOLAGOlnS1kS8s5NXse0JAj73cS3grkVBU5CPlx
U7GtOhXc8bMhBgAq9MXgrnPIyprv6R6Qha7oHkmY+BlxPCl9UnLNeUZoP/m+GmZ0Ojy+psX2d9TC
59l085xoouqaZf9GlpuGLa2HHT3wJoW9xTfLaGYDOV4rgET99wdywvmXlRcoZSCgissLZzl04qfV
aEmVA/mqCVTAsQvxtwQX55KMBWRSRzkzRjKPnnxdy7uiJl1YTanNTGcahnve7GZpezwXBjgoljJN
Y8smRLRcDodMAUQpH8i8RI/fIzMt4xljauWOvAV2giMMPg/bOvAqp5PkBU8H+4+ZhCzda25tUPNE
6PcvzjAZwG0sS6y+A+N5LP+h2S4Hexk7Dw9KHcatqqLk+hDbWummv+4oj3BroDCQx0oFFeiqdqA9
v+RtYa3wRt1fA5HRSFZMs/qW/Mi1k4LrLU3EE242TjERw2x1NWExuJWURvV9WDI5ZdjLi7qOmpRd
bWK2ESTYsg06IYjFbkx9pvPsjos9CDfzRu1Voc/7izQmcN+93P4B49K75Sweku/BYY0TMXvPjc3x
iSMdKPzMAC91tlSmYS6Dwv3CIt9alq7f0ZB99z+y/sqrwUJ8ILRA7lFMYsYmKn8u2YNnZoMm6lWM
Z2pP/EoP4qB231GGZ8cNaRwoTeym+aVaFCE9o0XZeBapUGdtVngk9hNgZXsAEGAeQ8UOsa/TaOYN
vRX6bKEm2UiVmiPA6OOcQl9L4LLb9ucebTTd/PI6cNdR+Ejvxfhme6oZeP5qCgH9bRe975KJeTyY
oTpXi0OIOOuw6OPyCSbMR5ThDGOHJ5xhIZ7ziT2AftW138UsJLf+uKpl+gEvyWVxOPUkvonVTebO
x+d61FAiqWSChsJRZZZZlvh0hOz3u4gUsU3PsaOwUY5gkgvOZY2IXNYPNhTGHIyRNJ3mIYrFoloS
TUJKKt0YxAfueMLirkqR3hwgzh/+6f9FNyWCXYH9o+JZXfkyoPrFR4dgDToAMO7LlrYu5rY07cqS
2VRgbpK5a1Ez6yjiYNwzH+SmUI2EiXu+F8czT6M/EgEQggyMej+7BSUCI1EFKfLvNeut3ZFCHX3A
9M07cVpT0zJt8XO5ALyT+2gVVansky5wraQ+zHgfk2Y4Nnw2ohgfMmjJAsm33bRU3SwOqUxxtdfV
Ndi0QSoCa+qCY1Ao70I2sDUlCRkGu+vrEqPApAs9OtJV9IRXg4t8tt0pyTWjmY0YgDIMK5VvmdB8
kWkUTUIqh0IlrCWkQsCPPbnJjO4PjXYiq+xFT0+oMyBfhEHOYaG5em8tmwJDewv+RF5b2GVCh0AT
E7R/ok77Wo+Hz3doB2L+gkX/U936wnrDB1xgIdOSC+VnRAnpj9M6W2+uf/jOUrdCuusg5irwC9zp
ws1SZvf94QMz8WXLh6R+1NCGaZIt9E0E7vvLzLKe32SkJMcts452bfI3eHUsHGjMnrp1NEUcCQez
dhMwEi+5KziaIVuUEDBbpRJzZh+BnH0JtDsFmMAfbxvDbbqEl1tOZQ4DIogcoEj8Bqa6sjRx4Ioq
FcAn7VJXpRjWbi/xrMsrXhNHALYUKXAAp5/l/eYOG39aqDUTlNSDskHLyKq1czzv+CcS5xmiXtGv
okAzLxrLvjyxxse5Kmzn5Wj6A6yyLcSoLbU+EHbuq7OEBWWDldocjwxq9YqJRH1vCRUYYVHnlkg8
l6CaY4t8mbI61Az2tETvNcK7uLPSHvI4AyHF6aUsMQaVPY+MNgYKTMOlezUJbPTBMFAhO4THUZNx
GcshmGNdK988RT8DE8pllBDuyb9EWsEewPYzxE9by2ZWbHHOJAeVvv+rxOCpWd/hnrpvC4JPoXmA
ObS2SYHN+2SlCFEPIBKehbqokmu+7cNHcGrYhiPF0aMW20sdDZcXvdHKRTkhxsB7sWNZLVohgURQ
b5up8OyVKC4Ayh1obsLyVThQ8SL5QJ6hr08opRDCbsPwd9F1B5b6NLQ5MsGN0NjZG3kK3r85FVSm
2+SEwykRU6B/3+M6P756FBJGTPH9JHPl1Hm9qIsRdVAN76ab9zFV0UhMh6nemwBlldacBj7XsapM
cIWNLeb5r+kaJacgH+aizd2EJWSKjd3A+c/8JaKx48BX++hfOlMlF7ugRKfgy2avzUxCY+ZdwAKr
Q8g5M9yRZqvPKjzrLNmSdqEHOLqkl8/0Q5X53kcQeJWiIPZg1v8xDQSOAwmGFHvjR0EgSYqeAguR
Wy+WJdKbl96ABBR1i+4j1bwhwdnLfEFL6DFBUaAEtvlSoyboozZ4zLUshpOsHKw7MNQZ5gR8jvcx
4t4apv2Tor8zDObdVY3b8EOAq1sEbDNvQlLAxZh5CBSwv6idAUX+yH2VPzbtIFQvD1IZeAKIbiFe
GvlnX2oo4mPldukzAjHx2OhKUNkkiUSzXR33IdC+VHO7xu60vU6KobZhVMaAnEGAJ/yKsOkNe2JI
hTm7XFEDIoLHTWzVVIk1AAtODABLMXwBOBmDGCP2TdpWvitvfmJf9k79aNfE/uXkEqmPBKJMF43R
XMMCetn1OfxXt7SpblApC9W8R50SDWhmYbYBxVtJ54VKyep5Nk6aC6wXQ5UaUQIIYLxTbaP6Kd0v
NS5D+Dut2cesJe69LVCPUFPCxzj8bg3snz82wuaJ/FOO7bEtq3JbNUW604N8/06PXqZLk8/OwRcp
eDI1PxnvBDnylMMvol6W+WkhzpDDu+dGW52n8bTUgcepSzh/dGATCfBZ0RItuDhCuqazY3x4DlTr
sYHpOGUmcg5oMydrGbjAZkQQWP2k3Ry0y6ifHUf0T/KXpLnkOlZa7daqcA9hteutTofyR7cp291f
pFeC5j2yXP6d0v2sTuv4163hw014jdY8a3UgQR3XwOBoH4sJtcufad1TP3h0BxELjqtQO7Ms7w2O
3uNlBvs66bemmSNnh+D7loC36UxAAPXrECVwTDXTGQMiZr0Nge6Cc5hPJoRTocatuWJa5PnT8yyS
ah171WIydJD8iw4qzq1JqYz+6Wmhnglumj6ybOeKsVXwJTBleCS3TL8iFCl52Q4D7UuH77MPcLyR
n37rWc/JmolnjC3tkmxPktkgP6LaIZHBNo2Mm9QG3Ml6YqTt+OmGEJWrLHiLNdQ6I6zpB+POjxE+
w5HqnsJ3r7ogX08bCKd8BI1Cs+0zngjVfx5oLVoZr9fsXEs3Ac3A0ypbIVUfJ3DvRYQ3K8XRWEdD
K1XxHYmGjbYKW2e36eP+iNP6pLsQQhe33yrbQdtTNd0KiTXy/gUCYSHTNGxgZw7EuKxe3H3SplKw
E5XMgA9MPZEoMnPUji4yuOg8YeodrRT/EDBeC87HUA7gneuDKsAOwYodFCkwgfLtdEE9P+TcibWj
JKcDQn947nUBgjNH9FORAjn3nRU63GNgnGIJmMc7+mUKyMl31WZ1trypSRiJzyLu9B+9/qRecuK8
q/k40rcjELvVHCQ8futM3MzAmKD/dIDpEUvULer2ZDfctWg9Z4S1yLbNTXKp7P9M+r7HASFGB461
qqNR95VE0fIBKfxgQLLQjPDkVRGSEbu/qlNbzKi82jqNEk4DmA6rMjqjSQWUXFsurBmPG97nqUCZ
pH47b3FjPZy48Zn+3+3qnx3qxkQBpTtUN/2QyN9MVRsJgEaotR85kvwKUPUeFnkk7iB8GqEYsg/8
ITXcYlL2NO1hdWlBl1WQCAZ3yXJnky2lTnKdEpBPxfCcAx2MtpjsbkGp57ODCbNWGwH/Yjap7BJv
ZNEoA9FFMCdROH47+6nHJ5GIJCsie0PzDLvDC3ArXjZLYI08DP7vAwCiuVan8KTuqZUgnqhmn0Kr
2o0z+cHpHL4WFbLEvH0tccLMjGofbzAW4Pkv91/kKfhbNYJ67pIAKszCmNcuRW/867F5N/HjuQAz
XrLeQ6b/TXjttbQkSwymfR9dHKpmFZ9Kua0iM1PJitXutlcWVAVRmRJ3lDdpV70l+gW5LKrG/vkT
gTiZGx63cmbttuMJYxCHGaqV4JzVYEk8NiLF899uG9of7Rag9Tb7KQ0N5W7CW8ErwInrEbbGJZ8e
4ZIZvM+v8qwiteyjOVZ7+oCZ2uzkG0K5jM/ZHqWLorN+JYtUaEJzuIn+VGlkW8jJjpVMjQ/xavxg
INLK+D6qJOgVUrI48q8WF83wwlIw16Vrx4X5gBn79aQis1RBCta17oAgSPPpl40aStK6ZQKSy/YC
4GhBmTnuguOfeDymPDD6FbJZsA3vhcspU3evrhPmVufNJIBEN1+w2C0EBJaIFOkB7b5c7l3V6wM9
kkaOolDYIjpmqcrrSlUXXrpXJpNhtg38wOssn48cYWilU1HyRCAClx7kJJ/9sbgwYI8YhHtB2axX
mZZby0lbdFhJzGGCO+MPx9LfX3vxQPaiYNK+dlocKatukesV6a87vbcQMjNayRrSKY7i8NuRm9vk
aKk9QlyPJTHAxqE1wfTmuiVRYvIdALPzd8UofBec9Y9Iny1QGQs8to5TGw/xcsnXlfiuSdr47SYP
gMapGAUDmfCWfZEnHkD+rKaIf/fLFnYBpNOtrGZWMMh1ryBwvzDpofO1sYS2spruYTyVi8Z6FwRB
SzunW3Gk0qRcfgd/qyvwkXBRxWuR+4/BxVHcAHuYTQWifeETtu6i+tqpdAoiNZxJ7PUwsYuErlxP
Qds0QCTL9dkQaph3sa8dsgJLsPlOD1Ivvgms34OdPnPFMXrgJesfEOBBsEamUQp/mrVh4dNr1FLR
Ja3F5fzmPr17RL3DQZ2/jGN0rxMseG7jcBJNF2F7uVHss+T1v10cnIV8NvAEGLLg3HkEKnkZy0hw
gicAhWzlcV6gXx7D3xVLstn7WB6CqFtuZYfcy68PdvETvL9ZcZWbPzBu7x3x/DMQtlkhw88wZT2D
TD7L87UNMfNpUpyP3KSHGbHUsy47U33SjZgm71Rpw5lL5ZLnNUGcHIpRktrQiq0ngZHL+d9n/Edy
kpF32YiF/H1qUbGXTIlCi9X4XxjELzpQbjGTSJ6yOmLBWdZ1moEKWWT/V3NRJPdZEZ+8Q7X/aDWF
GcTGt8EYAo8Eb8AmU7MRrpczyg8AiURO7DtP9jl4UAva06vo7ZbN85wHPF+48dG4thl1Tt/4zcm0
E6sACM2DkkSyDPqHwcB1J/0DTDKW6t+lHW4z23BNPnR89eIELWQhsuV/pR1NwuT5K1bQyNMfdrZ1
/LQ/RYUv3A3IxulwkYaoi7jF0RGBv5QMGbtXm+LVSMhy0PJU4DK7YMer9+HHSYKEq7WPUZOQmboB
wZrc2c1lMEPayEnydDGJLRM1BFh0YddawNxXGf62S2JT4xxwEgL1o5aeEA0DhOtJoGPmKKahJzbk
Y0wq0GsFrPWJDXXTRS1y3lqizTPc7VVMArkFbupiAod0mtTF+9w+utFKHi6BY2g3yrzQ9KUtivHq
nNs7dJFMVWSohJjQSv4Rwj+zAeQ68L5IrPlkilTnHvOmH3KMhF0UI0ZxAAcbOLmx+Dvh0+irjn8d
7Xz7dGQEbZB7HS1hzQLbaSnLFPcTQIfyUZmFVfG2+ta6yhouGnHVWT6yS580uV890AUjjF7Y8BpC
xqu4W2yXxSVTDQsXL8QMpHT1+i3DyATKyOvnw/RYN6vGLoY1CSPnBx38f2P4TzAZxp5zmfbxjZCX
Kv9O++D+Js20XNO9P4A+s/PsytXTJHfZ73MnjPW/w9lyFD4CIYfJJ0qi9uDQ82Kx8Xskp8Cu5/jM
QLtJZCbAeBwWmZRpXtvWVfG0MNfK3HGDMWVfk4pKNEUq5xorwUcMRFuxaiwSSwtArIeXjzp8j/+w
7MvKlK1KtZsM0Bwc+S12g+njwQ+epXEdHWwqj2EuIX32x3Vh15wj2lw9hGdu71rOId2Z78u/OpKR
EPNvd8lAmFKYd0pbBm4aQJMlCcnTB9kLhoG/apMaYy0dfMzN3JRx06LDrQ4qo6woaSDzamvcfK98
zJG4pbz68qQEPp0w6603W6L7U7pDImtNabrrPc7MMS/FV1T2NlrDRH4mFVQ0L4ciDoPWQF4oSRt/
bdWe1G2pe0XLF79f7Wdv1jfl5FN9Oo08Rei0+mtBhy8rlr/vWReGKdRZRMO+feB1kC7DwzJFbk3K
zk8Q3shmP6VzqfiyIYqH8ReWvlGKKpkRX2udDc2d5keuHbJyJ2CHzCJu1c/6VgROpd8+N4+HNmPO
2s69XlOVz//BaaYBY4ci1NRfAMqFdvO6xK4CqFngELvV9HPwBs9blOtNKvx8cVtRSa930JvSBxXJ
t3zPZkQmntY0uBbCF/VKXdmbqNmbgq5Dw3n2ZwcI8V65bcBaWnD+FWeV8DUSPvaJvyeAilma5uwt
MQWBoHcv8AYMe0vKGGRTQCSgz9IiXdSnBEc3OWit9vCqQOQuVzUHZZbzZmrAhJmSOSqJ91rualxo
gJwGvTRDE2M3ZGPLMmggwvsG8K0h4hmCjuNkREXdD4AgSBbnMAcJ6wTfqklC7E/RMpD6aWskKgS7
bIvukPLTvjH0JdFjyMSivArnwm75uX9KSuciMtHB5I+8yx0uEtDXTGmqnTNafpefYhmkDBFuV4Mt
6lBEZ6DyLzSq+IjbdnAdwX17MBdBggznOPSQPzPHbGpUGH4Too61AwRUtPgAuOfldv+QOZ6jZFn2
R25smtL1buG0pRSyptFPTkii8PiTfY342xCAovFYWwO4ydJ7UGzRKb1nVNAcsV64iRETILtxzyUZ
haQy6Jj5Ff3XU8585yMFgDEsUsHZVW/UODO2Jqg2zkkvMm4OzGDsCkr8a3besO6MTFGiUvCZ1Xjc
mvf0eoraNvmKw0vvgKR9810Mdjd9HZc619eWht/xx2783w9tno2t1+7U/ZFk9STG9MuKToM/1fKi
2NlFrSD7T3L6wRdUdW3BJWJxLFYE2gX18AtmeNYC2LGX1fTVHusuRaUZfDswhb2gesWzajBRogxq
OF8MFJmU3tvzL7FyrwDAeUVM2k09pFImjh5POwjpeLQPy3OKrKcTeg+YWHw6PfOqD8t7ey9LGzTf
4QSgZZlxrbTFWvXimu+kMyR158qDrnmDE/jFu8RvI602V5D7OyQ51Lj4gG4D/2fmA6prskrSHnoO
geq6flJJSNZv2bAgPSSh2zInrl/PX0sZVvJ+Q1fb0wYV0vKH/228YYhP4hfnSM5SmUDu5F/l9Y1l
U0ZV76cbI0Pef6ZCvpPDz1w1ksfS3tQVHh4fpJct2mRHAX5Dl/7TZF2LOGR5lICeo98TMmE0Lnuj
hzig4XXLXJh6riDtj+Z+sOdBC5C9eRmQFH6kPYEoyFTJwcBmiiisjcZxlSBbpryfQzC9FNsrsH42
SMsstk/JYFJXMUMfqGQtQcwiCNKC61eCKhIP/xK+6n3DoSD5iHpe92+yeaMczSkdRtjPIRjK/lO5
wvBNYgYwi9utlQBqAT4bxQQKolju8Lff1OyYLs3dbZBzlo2oB9M0jmwHhKNVG4nIR6PTkn/+/Gvc
DRHv6j5t0zbMRNGhfe6PfS3BGN8aVmV0cmSMbIewny3j5w+LJV9HS75sF+q6GQG1MYzToi3N2sBV
6O2jDveHGNMdoMIhYTKffoxLGmRKVI+/nL2NY9GbhFWHh1duahjr2kyrUOddkLYiHMzXfiufgfdE
P2/wbuLV+nx7V4O7SjfQgfPuiPrqqaUYIg8qeOxdCSmBxz048Nj39Aau2SB4m3jJz1rYV4xqRO84
fp6UrTc196fBGurCF5XPWvssDE1AWKoKiqDrmeqvFOcwcL+ykOxy9ZMzAAGWr6FhuPgcYaJBTakA
2jDNa6o92UMKpzq2IDG6KGCJxeJCRdnxO3K3WQMCRcddMR5tn3I4e1zo2f7oW0w0vcOVRh/lrtam
I/oj5koe0FWfWWdBZAPtHc7hgay+YNOqN8Hgjhp4LDXtwO2gbPp3b9fe73CHYAy0aH5Z2BCF8S8H
ABckQHbYck39GYnyWhaL8cj3pzoKlNt6o4pBuuKoKJNsG1VUeoMVHHh6rP3+L5xklXHa2W58mhOB
VZ+vU1MnauE5VukZ7PuzTbPEfejoGOcssbLnrz8rGPf/ayhGDswUmnFHmf943UgqGQ+dbXjFxAu9
VaB50PGp1HyXWA1YrbYNxOq84jGmmWj9FGWzI1sNJvvWD1qZVJKa5grTXOW5PM2Unn9w+4aeXN4N
Vmm4c3UfMBCvs+AgkyIkn4iItUUtl0pr0e3fYkpJzVfDfVhd+7Yd9GQR9kBZTkifXxaS3gKvafIy
K6XtqfQF89oaFwmAKgrLZY0/hMyd9NZz8lvjZlGat0K8vNCFwQJwq1ZI+KpYPNiEZR7Od1apgIdj
YMpwtYXO5CIR/ICqt9SxJBSLSWDPZYUVzKFoNCDU7NI4k7J0LfYpHPo3csoLf7kBjNYu/QNyBxG/
DybIDy7CdJtyyi+4tB0ofJRzqTQAiwAghGfilacpdCs3UsIsyjYk0Dvez0d8CHx9McGK22dTVwYf
y09r+dNSIgiEhPKFx8UhLPr0m5AHNImW3FN+XB7TpAhUwmgQihw/pUtQB0kFz9xak+zewMDol1OW
IFQZm1ofOCZ1Y9HURiOaeQpRmh3T1r8hNbyIjzdcYtlAvqLBHnUJx4yGW9eta/gr+3cz6IdOTpDM
yN+fkJYk1LpuEpmLqtrVMfB+SgD4Ezwv7LL1APY8ZtF6m4Rovbv9NkMmctBPZthBidwRmOo6ktuM
L54K/cIih5/6zYNfdkULR2mA3oTcBvBReiFYpRu5L10hjLfmJyN0bX+NlCtIUkMlfpiFUwf4Iui3
TwpwqHDWR6r4l+2xqkPucThxo0IGofWUbIcc/qoy8mcKFaOhXuI9QIh+IauYsym74/M0/xSm3BXx
z0fGLFLI03Q+fD3KoWLzxBQV/rj7D4W72mVRSf1PvRzgdMPKSg2UVbJ2+/y3ssktfXiZ3dk3/eZV
uXMI2ZOlRxDI8MMn134IxYuK0J4Z42br2a/JNo+kQjIsuCyHEC8HS+dMspWjKpKwIVbCME3PqPV3
ZBvV9YaeVaQIb1pys+x2uUkcgNAkkzfzoHgoDWqAD7lI8sSP1Rx1rMVi+I++OOfOhv+1Zg5/c63x
tnpOFf0ut+tPydIV+ZbgTZwUMPYjFT6CRg0n1Nb/dfQP21PMyvin9RXA+7VTyD1XEwggHKVaKLPr
tdJ/BDwXaEGtlhkKgcZfAfObdhBJQ9yUYlvr1Msws3mr0glHBFRO08IaPylT1GQhWh2i1ZPG1Xz8
zLM8EEoxE9V/qdJclZ7On1KGZqTlUbpaJ4Jiax0+Q1QrVk0CcEPmA6PE5KPFBr9tJ6jcMMmKhHfO
p550Ro80201KzDZkCx7qNJXF7zJACfEcvaj1AVDRCHfrKNz5Kp2TZnsIZFwEmUJArzdSWSdlUmac
XLw61fNyvPg0sn6Kf1NgEmsWL76Nc4IYPrhNDDbKOu1inxWsOIZv6rhWJ58DIEc+e3sAbsW4R8lR
XEpdtRPdX5WKGLZhBznmh9yFbTXGnfT2uay8d8scFxmGnwA0ByO3hA2myzgDWPvEhJk3FOltEVUH
v9FmFlnabbW4yFQHugK8RHN88+VEmjuBDYX2Px02Zs+q24SEBSpUWC908CRURGVQVLSggjyQZDXW
QPs7PysFs4Zo18dsti+ufx7A7XISSP+bGT+BPnJX3O3IKw4KB+1+44lGW3WjAG+n5/MUTo4am1Ru
PGcLZr2KDw6ZzRMG8ClrhOX1U1UnWkP4JjuFVNDq/sBTopUIc90G1CK/5bgOsgDbPwYjcDZx/avr
mc8NFDYZSFNWxCHvD4hPUu4r54AySkWEWFfB4lrUnZBsO5FnQ8D6SNI12mrhUprwmLnilWEJneCs
Ubz4vN26LwKJsPoStHPCofcvCLuTNdXDjmPh2KEbtDqxtwlJhcvnoLHF7dPI6XUqJnGm0MeCLq8K
ZsmSrbuRQOHqxLYoWjvjREJCGUtjQ70ppHWDldYWSrxZgQ18ZO0RiqirFfR49OGiP5J1gvLX/V25
OjKhYNf0dJ6vZzym62NrIsNXtXk+L8/+rRcm28vmhP4nxwbaGy8o/Zw2+tpC+QSKI8NdfnhD37yE
rA4EXMz+CVhxYBo2BGWzmBt5bcjtis5dj1WBb58CcDSc0KFgBaJ8ubxCzpkLjLC0AjQP2s/OQcNo
lpsXTGKMBJ1mz1Dn3VfWBHPQglpegkwCT1Nm1OhHXRi8PSJt1987JzfQNfpSIRuh+bnnjCMy2lhg
vvE+L9oMW/wBI4HIyoYhZKzJDb1WeguQKuUPT0uWsh+sv0d4j46Chm1ZR5uuAfGXLrhA5y/BzoDK
alFey3Jxe4ryxuN3lSZ43CIpRGwtjrfGljeP6m/Bqi3m7gesVn6uv08N2YuIPUObYMVM9pk3kC4M
c/IZAltxERVw2FqJkhhLJUXd5kJ9kiJTKuxfxagKY2zQeoaZPGIlkqHQbXXRZPV4Z3X+yhtehJtM
Mcsd0d9YbpCoMjhtJDqqZJMzRUUgVPsRV/1itgXeEx34TWMwMyxy7tyuHUCQ7bafKvAG+6nEAKMh
1sTi+HOA7f9unymhgud20U/uXR4wJq4mTOaCkfM27y6EbCZFYkWXqLD5iU7IjNsO12yIiD0K2CJi
FsjmFUMNTkQDimhnEZ4QcI/ZvMaDZXsoCYuvfC3TEPcj8oQT7Ivk8yhFsKb+CrwjMS5Iv0gm5ZZi
WTw0oiSF1n5lWBFeYHmPD903hJkddcjfy/iznGexHJaNv0rI221tDBD+3N86s8h0M0A252PhaZZ6
ujyAAQv9Hs/GAWLsJMxauPGmxTEA3iV/P0sC67K5IZXG4bCDoxCzVmXXpDFJZyt8D+W5zIz04uXO
EGKdmw8OrMs8aHxHEPUFve41ZtTs+6VBL1VnNY1I5LpDotlDJkoomdcSB/NEnEr9mWAYEY3NQr7L
R8yZNJr4DzHo80b0EC9yShpWPFZqyIrWC/SU2FHe5uOF6kmgbqkylMtLmCojJ6XGvr4ZwzPuKnav
nVXZGIAZuDN0Y/+AN2ypruk4Y6FODi3HUDdLMjmGmQuD/raDCRvlyn9d8VchdNRXwOJNS568TvxQ
U3qrY5tmUqrGfLQLH5/HWs+8MllB0D2EVcVKZLyYvV0tB2U9bUU/pj1uugmEKlQraww2QYhnPtjv
VxuWFwzSbrpCHFhXRcnSUYIKka5iAfeoUbmuQcjnPD8IJzOuvm+u/aBUf/ljp655ysXodCddnlqF
/GjNbgYwVUbKFdF1eU4yJXINphIKV8P06JMxxi1bXdnc2EcHVajmil9P8a4kxW2gd/NhPKnvMGJs
zaTGTnJBL3Xo0DWdkz/AevIJUnxWLVq8kwIGCm9FXXEIuZVqR3TCDRuIOrMgQlhfzEGnkjZq7ewj
akIBLF4GQ2Nu2BEE/RzLluw01s6dt8b9fA9oQcm7Vr6VPVwDx3P8R6Be9DNgG7M1rRCg5OTrVudz
X8/TLqDo57Wk24q0CQY5FDm6YKbZW4bb6P7nG516WE7TwaX24sOmllG74i/7QG5nPTOEN2CPTCUU
fCHBw9a9joRI+A+TsgfMZplqewUjXd8ywzeeBhjCDYdTO0nr2Lub9i7D07pcNzBQiVNwdhcuKpnO
F2I8yIwKTw/ssAmiqI2nDO2kKQMLlWOahdJ5UKHltKHqIrEmkD8j++sYwd+GEiEz3Wlzd16dOaof
f/Slu+iiX9GRm+bfe5Rlb8wi7Sszrq1j4KRAcBGUcr/Q4Mk6hB6zbX9cIAXMI3hwM1/kqa3ZvqaA
XQGZ+mjXtiAXL7SAptWv6UG2Cj1TLDiZcwEx0qNG/E+14yS1QUbMn3ZWTYAxdOc93UMcJbbMfOoY
UONd1P2qnS02DJaKS3UUWVgIG83zS1GhgmdA9lr+GSz5lRtNbtpEv0PNtPMDm2TQkG4KANiYGAiH
jIIT8hV020pgezY3FQyhqqNqoVZyeOZdXsjS85ja+ioy4hPMteKmSh5i8xwZ7UGoUZOhRYFwmUWx
zEfllYEiRPXawq1B7nBThe6XL5Hlnhx/FdBVh7Y0H2wW8KKsldaj5GGkUorfYtQVshJGEiovAeRl
GmDk90L3WPyfnHbF2kbzydxA+eM9U6xmo0cKeivWZRDdSxlBwgQnxQzzJsKeoZLbgE8pXi86uRtd
bb4DiLO2dPJj9p9i/0H2S5P8VJrIBeT44e9m7koeE1jNO0z1Q1EsTntifAWVsj4/Bhv+dGxRcIAq
u3Q0Ib5AUZWKcwVrjmY2SHKB+3/LhNvN0SYCKvdgo6htDxmYdDfAHIsw6eyirwyUCwjAK5ouEswn
q2pzah7n2d0LelcfuukzhkzRzjWX04trqGR8f1YWKIPSji8P/d9tDJ3xEPIImY4I0Ax1e4NrSPKK
ameba2MXqultFstni4BzZT+Sx3b942VQbqiqHJ2n0U796B2q4ZMrNlmWzqkc+2Nz/z6PhwxrILne
C+fJTTJN8u7mj0ztmn/xLx60TOnD8Ast4HwAsAYL33pDgRbhhqNoewhAaPMlackkDCutI+Lw9Tad
kVZ2hLSi+zhYY9nI2/K4acculj39E3pEhFQs1q8iv/pT88MGogyMRPzP6vIZF4sPJ0UhyrYqJk+l
otCM20NdJcPlIyWzDOYzVLA9lrkFS0fZjsab1LoKQ+vyvRqezk9iQE7OsYfmxJYp425LYyCRNOO+
Iv8kDgtvDd1I1lrju08Q5wPRsFBADHU6aZMx0KsEd4kdAkzXk63rYf++HPcFUVAczqziPjYE5zth
UjIAo6V1wqq+Rx+qKsAkA70or8c6h45CinrbOWDDKt6yOoZjobk0otFNMX3hJTZGJdwnF436gWHN
GWZZlCv+XtaQIW3FL98VoV2RGU7J0RikqPILDDr4jFoyYGO5GEbAkuYqvXVIH8Xnno2Vecwnu4TU
ry1J6Xe/zpaTxMp5pLJAsmxAUX4/ym3ETAxQBf7xbdeaGV+a83Ub3bYrA38iipit59VQJszGuyzq
MoihGaYg09iX0IzfVGBTf2HSPv4lI3MJwa0Aipvf5IA6IynCIylp7JKA+u96q6bnaleWBxrkZ0s5
GRngfsX7cVRZAqexWVan8Phjbj1+86Muk4ZWo8wJoDi7sxwBKPwCREOb+VIDQL0biFCNXhxMen5A
zSPL9hjnzvJ8irMKfyAKfPjxwMkUc3Prxr9Exnt/amc3q8esquS4dFY6uL3SNkr0XZjoX2FzKKIR
6BqHoegyNT6OS2pvMiPPmZwxh6Sgxn8v7UyR4e9UJlCZqHbxzJQHLCVCNrO+3ZX84nU/7n78wWM0
52DUNf3LSg9QDIiB1X1wOxaiWsQhrV6xlKOe5M9zh4+fVM02sZVVf5Hb1o3Q6BjMVhhJe5dLGiiO
HV50oNns5BYkbd94mx0L1u6WlAd87d0XpbzL7ZaT7OLvFAD1IO82cGgcI8CwTl1YE5M37AnY3oYr
IPbZfqR+fRzNb9NJrCKkmxTKALPVsRFgnwXSgrrPKmyQ5gZNOLuhen21kereTyRHQPIsGBHTvZzD
hOZJViRK7CA5C6nHmSyeKjJm1tvbx3vTD28LpddAJ8I5C0UlhYNwkBCD8OSGKNhlkZQnxZHMCHI3
PLMkeW+cqX27LqJrTru82CwLWCamferc6ztnkIIQxLTkyb8NRh64m294qwIpr4TnEiTMcLRCjXQP
9vLVNa9SA8BNfgPM/VVDzrwOPLAxvMzcHjXCuG+0ZyoTtDzUpv/e2Qoq7xX969OKSWjEgFgooK+R
28iwwH0jDOn6yxVXrw44JXNmKM5sPSIKyJgVg6vGv/3YnaiR4tG4GvKcvGbDCcMCWK7UFV4zRZ0O
68B0Pw4H/4q1f0itETu5x06USKEoHZd1mWL+kIGpndaZGSeweJU6goTPi24z07yWhdzY+GRXdrbn
Uvpm44qGx87oCQNBQTNIMCUTnfppTWMcqMbwLmYq7dClJfH0/7qRmF+mNNO1+X3iaDTJZ8pmPkRY
pMOEehXy1ixst/vQZiJqtzDrkjEpOnDSrVZUbkUbdN0BgwPYIZDW8o3gNKk0bSYsc270TWwhfIJf
+OK6mAS8a44wDGOrvroU3C3ljlN/h7It1Qpxw7rJU2D42E2qmco0xXiDqidbu4Kq1/ZQtBvrRdcs
urW4bb/TrgHM+IEwG7H3eGSf2K0pL24BmouJ1PgFo25TS/naRmRnU8Ur+iUitxTKI3YKW/hIv5Fg
Of922bBX8AkKzRO8VP0nI1eZ3w+pgdsjV6svTmTzJEXVSBN2RgU6cT3WsA27KKVGW4GjhPGejM98
kvH0DWe3XAHGCDceZqLpQCuhzrBlhnKJ4cDn/tG5zpfIdi8HSmfKh1yLVCC/eMyuSvdJrHXaP0TI
RbtqX3oj4XdnrJOHact/eQ63m5DS3zZH99b3myTKTtkt0d3mEFBydGCSIaLgZhN49ruzVnmQ15of
Yzr/XECiRw0K9iK1CoiexqkNKDat6Tnzdw5rFGgsmckoFzVLLnq5dOvePXt6ECEpTTxY915/BUSx
l9LaxMC8LgueMeLFEtVmG8s159pLysrsrU3FBDnNuElWUMPOeSdkyq18GwicA5t4m0TG80GpOiQx
6p8rCqTl2w+3Tkxu7scuk2HjfVfdhlxPHutEf6jQgecdcsP9IpUpmKRJKOifGSG7hrdDlimj2f8p
FbacpCtfoiCLwLyrZHK5Zk1iFSvk8S/mZ/Cn8DIilxp8rh4FtdXcI+iaY7AZH2hLNXuigs5AaK0a
E7JuLfe8H3z8Ut12j+2Dz+tVWjkHSdLZpEyCE7/JcjVbnUD7HEdkbmXOysX2V8VDrBaqLbIHGV5/
qb/j8MKlaAmqwt3tx2IGoHcIDhFpCCtKvMUgnaCfaiEdU4gLp3cM9C2dDwoeBATvC5sjUPQLFnDp
B+llOFI5fnFRciG3sx1eGO8iV8AzdrLqlzvyhs38upP/ulKpc8xyZAPX/MUp0ej1DB0xjRaw73Eo
XkQGUmA68UkVPVuNEuRaLS9TvekvhwH/ypJcMEUnoiC5PQZdLYa9NR1UcJR2rGpTtNn2itpsIhjS
n/O5L9/G1kJoa/Z5IuL6mVMS8ka5yjw4v+P29QVP7+whX5ooW9Ju9zwpc5UR1chbgAE0OMU0tJzp
gV9dvdFS3BXRwlAq/0ScBEPqkiqMNDFrHfolELlgphvzuRR6SiFkJ3iGJnUbn9NKcrjBKpCNtJBl
fDtnVYFrlk2GeCLGggdnSlwiAc5Lcrl/VRegx8RblSm8l4BPFqYyuU08nlynXtNJRhGbt8m8qEXz
MI6fTqjUgpkG1aucxNGC95BS6DtA6F/RaaSFpQQ25EppFK780v+ZTFphxJOqw8kqdJoSXuI7rFNw
gf1I65DoNBVWukFMpZ0fea/OY7LFgeZU8hNgwsCXqc40V4vbauZeIb9SXG4QoR4AeFWPE9vQHlJ5
d5eJ2fe4/73cSkwu1bks37xEtTEsJm5LA2HsSu9Rlv2JRgK4Jbejr6r1Q1ScpQeOXxxpdBE+tbq1
HY0Vlf+Ym2uVWR12hvtbEEZ99auJYwk3z8au79n09yiDwOV5f5cdO2orsX7lDDpDYmI7oi6+EoC4
OxvcRFTnhv1OsDZWb30r/ZS/LSsbrdzkLOQxgZbcU5C/XhGgblc1s5C9L6dniCMRjDRuZA+o0VA/
B53qlfqK3IPnVZ44+/L4fGs4dCcYVYfH1R6LEsZ8akkPPB0lxALkUJ3imaxjzSGXEHasuBVgwggX
3vstU5mki99vFUOelsujvCAlR0msdbWRPQFk2itG4Ic+ljRwk44tM/AziUJra40yAmdT9Mpx7zbj
LH6zpyB8aVlk+u3Q8s67BLK2rYb2w0az5Jp3g37nPsggvM0o3Md7qQjlATmEfva+SC9ckbK5206/
swoJ8KR0zJZMmAXyVVkMmIWFZ5vjd6JDVSpArfI7nGyIeEHdqBNgYqoHLUulnP35lHcVlXvc8hin
ljHrShosD8Xt9JtexarORwqAnS35/Ko8Gg7/cNglSMZiN26B4n2XtmIDY3s2e/MLMAHX9VC5HF3g
xn88FVfzTIHCJK+2NrnBvCX+pC1ZqJkuZ0KROa52BEmZ6Do0MyO2hTmhxBsAmLkQTr3gxL2CwV67
mHm858Gc/Uuf0uz/AlSHI3SEGehPM/CKC2VpqZcwWAdx75HjYJycdXqNmdoMedr/sp7y1zsRxH28
9wP8FjLe7hQpdRMLBgkuV9vTx6buAhYmAN5p4ZzAxp+dgk+jvDwIxp/0hWfiCZ4rBvzKVa6Y+6K1
DJAnfwSeQv401vtd/viKQ2DbcUmUDuPbbMaI22Xpu57b4hqXZtW9LOuJrM4M8MYtrj3oOyMgGfpZ
J821pe1dYMBCTmob09NLd7nmjhaDsnAR4IcSg33gKubQKGIwe0nSdJPpsa182rqGr3fbyxukza2B
Wo3XU06ETGE2EwmDrQWUsyFgZNbHZyqF6n/j+iz0m5AlIG1/Wns2OB8Vk7AAdZugXiMo1vHnWMmf
dZ+sdUuMXR2FIRQ5MDGmV5W78aSA6alcVBFuWyfjU2A5b6bfubETANltF7cC8FYAFN+YXcTyzRv0
RDgsHnEv9lrbaccaDD6Lm8aQ6WS5k2HpvKEcDkNpZ8S1iZFABu4vUR0ExI/IX0yWHhWraoTUoQge
4kwZz8bc3TH0ecRWsMiHm2dQfGsOjvBz+dfPZ4+2KBkSk2deVzyQ8JnDzwPjROkbchtY5h4gbdRv
LGXAWrZwi60P6Vu4QM22YjL3LJJD1K4CkWW9GExzeXP2V+RlQIILGxdIRlfIgWGSzACJxYFBjCpj
xjBjsuuOpsDqAh2RThIgli9ZxMJiaqxRC29u6Ptemixe4oGiQ5eoj2LUA9ekc4sjsKsSREBKyRR5
x+bqI3bOruO4rijbsHBpiaEPmvrXaIibvgTvNpbLJ07sLPzwwUI2BiS/LygW2h8TNaSyQZY4rHmO
kryR/swlvCml1Q/pDjE1Dum/5MQ1VZ8hsyOZyYhj4gNLzf9IPRa8xuLB0W6zgf1uw5e1mBWu1PWB
yIIqMjh3HeWYS24jq7TaMLIvjkPEDCT2H51FI24FfXnbrJBdNk2sEePE5lxmNBcl4bmURVbvTFwm
tnaoVgt1TH0HpK37n4L4o5zmSifrmrsJgHJCNu18PtB01mryAVS7ggM/dM54CRe8kYswzwtt3qWw
+odhgncnTvvmoceKpNnPO0Y7xPZhsOQ8IejrfYrrSxz8ollZTwv9Ny2+o36GDmnyJKsEl3gSvyAJ
6eUEFIvYv1/YvKz6gpNinTtonY85/PsbkgqmNoKYdWhtP2OtettlOPPlXCj2kujrlkkIHEvu2NpR
LV9VQ7g4L5w8z9sjsO0P31LghmX8mRQ3DT+h+onEtdKM2TcOK/YorptPB42XjHtcHqFfoZDr7rN5
r9b79IP2DUMGpSLGrJTRQC8IdUoAv7PYvzF8cel++9So0BMnYsiWVHqoNYOlBtp+aRZ9AM0xf+GE
jGAkr4FVeHBf0YxzLjJKOGqjJh+yr2wbH5oFYo8ni2A6ckhVzAQ7PfV5wJop0J5b2By1hT68pVZ+
xlFIMAUKpflVZ1d7bj5fRFe7MQ2IXMplEk4onlu4Sk0pVhfALsLwUwkKW6gQ3PpL6ZUeXCu4wxeY
uPFHpZHlpGWetRAmqMs3fNZjCERicGO9EJ9vI+jIeZR65w/gfpWYXyfgCSUYnPeFBoYvruTl+dt/
2rxAIpIa0QCrkROcdo9HjENwFLm0AKFhKNULBNNbRIeG7lJYDOMbGVXN6hhDJqKfcAseGF5f1NgT
MSFK3F0hfiAdXxwy+/7TWVhEL80T4auEh0EhPI4PKsH8asUOZgZ9sl/yBU0f1nuxJixJ0+LGGUIA
6KoGQUv02s7bz3AG/QMFyBdTk1xoD2+r9pDaF1jqGqmuQ21VyzdwFvF7SlCfOKQza4GN5F8/wkVS
HYHjy+6HN/gRDpRbCwHgIVyXmJcDNmEZPz0Ouc5cL70CjYwy+2SRP6iGovSQqAHgc8MDX02ib3Oy
81lYbKg5Qhvjq8/47opKChBzi6amrRF13IycjFv5rTNSL0hooJ3/PXbxjuon6T2VEkXtpg1LbGtt
c9ukr84cmKZTqm1JoPk5NPdjGNrQ3yNnF0Lx8nYP23Et2yZL1JW2e64ClCULOVMIoX1BRIPuMW5m
iL7LIlQE82TcnRsm+8X1yq8vfPRinKzM7cXhADdXz7SPqtFWSnljSszMk4aQlS7H+pBixGV4h+t7
QtXt3DkT8ucPEZrVKzyKfgegL/k4EvbUy7UpWZ4C7z+FgdzySVaOouLqKI9QrmOmSrN2BXpGf6pZ
Q5E6NBgSR7B3Vum7tO5Xrf9VOZwtSfitKrMjMgOePJhgHrxYjw6fDl95qCZFK4mrILYchU9Fb1HK
VEo2LxrFWeGgqCOCJa1XiQhBGDgORX3TZHCWbng0I+jSPECCn2K7oXYuIItbrCysdWl2rfoAzP4i
V6JuqbILNhRywgiXRGoRmDOvf3yxht8wfvcxCfPLtEzCwG2pidGs79sO9EiqOLjy6NNYa13Lejzh
bB5T+G4PbFaeGGACoj7fh1gdMLtYVI7r7s8Ajwu2sLmFloBuAmm+hcJeVPIh/FI0rIv7l/eQEYtS
x6DMW9lX5tmo/k+hsmboG6dRakSXx3aqbx5mes+bvTq3qzss0+2e1xtqKauNs04xDFgUMonD7p2D
1yb5fHA3hIa8v+OV8CUK80T4/WwngDKWRp9IH73wB6w0DQNcPKC6vFAQ7pbJVmsdeQhMQZloANgN
k+jO6+CsBSaf7Nwnk6Au0rUVhXoh8AVmPDFI6N+vRoplLsq13sgwS1T2ciTTRu41l2ultQ7xpA51
ZrEDZSNZ+3hVhlZWuf1h40OObDc9/Y6Sz2MHWkOYArcbrwg78o8xH/Xom06aZn1nxxx/AJ2y3psb
+GencQ68NpYTKIqBUFe65w1EmEuB37dqLY6WmjDZ/iMojK6CiPyjBGmSgsEN6rAb4PgoUgeS5CT3
6+Gy+R4CsRxhQBNn6bKyN0KtZxjmXejzmQdU8kCBT7x+FINcwSHxmoeZCt64v3soyQAc2AupsziH
VSYIYzbg2U6ezT+LvUeJDfZ1uUn5ZaKrT56OA0uU2M7GbEgYmW9UXDROLuwKniR+/HQrj74sFtPn
gZ3RBwOXLFZoOWUmlEUEiiHfdtHi/UGZyKwyHeBno9SRlJdJg4cQw6v29gGLnyJGA0AVNNrJox/u
H/gwSVhp29xkHO2FiKQYeI2mqN7U6tnTVYPdfOkS7FypIOgvBqbtgsOIYyo5JlB1fAcu8oMVkoiu
VfXOPee265K5nZr3gfDb9/r3+OtGSFE5qubDB+BisjlNXR7ZHOtlOKznW90O0iHSMkFJ/sa20GKb
joCvu1OcByKlAOUscF2O46UbsXIgd+L9YyamYjbzdg5fYrf8VN66o9UmBv2ckw9cfvuz5qwjMNN7
Sz9SZA1zBbWhohSApawUBTzlDyL6uTGjpaK7BtEjLV9sBtLCcRSZSJp0r9+b9x8m2ZAnKXeLNoUR
UOynHztmJtw/0DXtK0khVeeq76B+N4IdDEUxtZTu152ywTsJUe55HZxW4UqR67P4w6oP4C2z8Wr8
aOBLuxjTwOe78bMtUVPexSV0tGUYftgdYEJAbKGH9AYKfRPNF5Nzk+vACjZ4niyIBViVvvl9GAov
jLWmzpiA/qzTc/4yJIBbIAAuE1R3g4tlOF26sJM5dC6oj1bY9imN4jhqk4Dr7u3vCzj5GJb7Fklc
uFf+ZEmiuAAD2kYTL1yWo76RM9Ea7rJ9cqCHq5eI7e4B9O+1giuB0Pc0BzH0aYsq/dF70mdbczvG
mTxCoWZ8WbdjNhQEkh30fsYVRamcKkOQW90mfottU7beVFlko1vhIvpkx+wD56qyJnGnZLSX5yDq
dDjr3qKepv8G7E6+hk7Uc20UlVyJqBxrfy6lmtimYaq1TSj8oDISUzy17sZFlq4CiUihyAi02GbV
Lo4Lur9z8nvwDcHL98kLaVWqms0dIMazbRW5AvOKy94Pwsq+XSLyKllOtikPJU4FuKz7oZyq80hF
aGNO6DpCwsCYVDy1YCfAE8C5/MquTKs88JyFjtw8cKpU/nQQUayPP7gfUzZDKtjy6H4KMnDLXr43
ey62sGW8WOdhP3mR7/muPfxoaOsAvlIetp9KtE33hMub3g0NXo+Lb13TmAhEOqYV93z6ddJqo+4K
i3+QrMv5mMedGXCgf4edPD45O5TVSdcWAhDn7TKpNiiLNrgs6aspYm4QQPHFA/oxAZ8ZU4r04SLS
pOe11KCpdoJWzZPHRcNA204GSu1s89tLC6GSmOP5yTbUKhB/1+Es5Hvq9n5XAzj+GuLI69/VpKzZ
88RDMJNZh5igY2oQqC4Em1xTplhy8C5yUBjFoVv0Y6nMsVioptk7QzI/oeDBqTQHjaBd8azHQejL
Mf+moqS4sbbNHa5YpitEpXmggN3eOpga+FlUQceRRQYIcjzt98czsVD5WjN2AFXGI//ywb7XGaYB
XKqxi8uQTnElivE6xD2OLys3+Jy25g1OF0RsE7fozKHJwrbLUdkfDiwKCUSwkCf3vKqx9HjUdd58
4xn96yQM+8afZGwtYh7md5BH90iht/KRDDwfci06a3iy8L1ne+YaKVkdTvY+bEutKkKMjwpGCZCu
w0IJL/Eq2pUSsS7N1OHPVu/Ja+n+EXBzkkpo2m6NYv1ZDy1XVbLzr17+JYqB+WcrXn13mCmINs43
AykgR7ocT3fS7GyMgjorFLRPLDy7PUSPh8QRhQLBwZtDPJA+QCNwz99kIwZCSbzV9Sc40GQkH8S/
/sij7uHz0Ri8b9VcTWPATmzW8GuaVKT3jItwJwhQLNeDUWMJUBQhY7vb8mIMSqJdEGLw1rWR0vTW
zcCN5WdApqKd6iIhLFzByRrdBWEd47Z1I4+/53fJTl/wPhLIo223dQX3sHUJEDzgihHj+1FS9jSB
mZEC3dgWHIqXgkkve4gjebTxbjYWm5Hj3W9q+kcGNZlhF2Z73UMQLqfxHio3XC60x9Utk5bHj3Ie
c61us1yFlzt20EkN2gP2rngoMhQf2wtXvQMcUbJ3U2UWXsKG0Ni10BZ4K0Y87gSJyGaQAsUWfxts
3Ur1WMcLtG6mTBGNx9f9oXiGEVm9jO19y8e+IPupTs1SQ+cK8ta43MBHZedvusgTImmXbKNotflF
QcDbzMxVyCZe4b+Vt0izRBfdiTS26+H1wh3UgTn2HkDHyNpHV+2RUBDLAiHP23TbdwnfyIqsJL7h
ht+F0M/3HAD7DQG5lahnXkV40fUjgNVMNBORrMq4LoGMJKL5Bqs7vThH9NBuLcVXo2a9SzgH7GLY
P63NsnKDAQ+qfjMZZiqjFLed6IVM1gVX8cZUuec/SRcPQeyp53UGTfUw8KZTszUhQp9Dttoj68hO
gUfrt3Q81cJCFTLAM/0M2rfhO0EjeEj09+Pr/p9Vt4Wpkz5qt0DCZRbDWQXfk2VJBE36euTbjjzl
id5enJL8o9xssSHYiq5xVCTxAy9NIMTj6fWsyPWVjWn+f+50pJn8rYh6EhcSYkEZMaw7er48yAc4
2SZbMcmDsOV6JRf/a1Blb99oXv20ZfGp7KyrfvoPQ0j+DqgvEeTFXgX8y5PGH22Fi+jHyz2/M5c9
k+gpTXNENNVk8okpSK5l9PaBtzYQvkBTBLTLhGMn0ozv8FCntsXasGIsTlnseazzkyLukRusmxuW
kYruI1AaaIxxByDY51d7uvNLwxGa+SROCHdtMHu9n2Xf7ijR93NML2DNMUwqQSmaxV+ZUZ+SvLhk
Bw7+aohPJUg3es7eJNa7CNsCwu8OSWFfkT4oS44kNhdTmpv2r0yOmY/fDErjPX2oKpx2QKf3jU8K
Vl/1cNcGuOApb1jclYloF+ymjISet4IpbUiODrLw2TfzPviZoA11IIKP4GxDjSP8IfmFw/I1WrkP
IIgF31gcMP410HW868eQnSSBVHpcjhatfeOwMVYIPO3bRfDERFEUnjSY9dxk1OhJhRfkmdlLkU8a
HNERtRNcTFlEoBylO+kpKdvxbR75wK97bnS1ixYc0mZ7MK9l/SRWy/F74GUWt1DrIDBw83QoYHrb
+ZLNS8ZOxEilvqknWjVco3WI+zzwBlo5V0BN/u04tVctVSHqrJU/A8aA4q9GeY7K8wTPZXv67P5v
E6VQMXGYc0wPecX4Dv4A6eMh8FlXk1HD1iagYpYXTKvlUcnxlj0X6er7qLKgocUVSkTis9n9VeIq
sUb92E/0pYPqZeFHX6+Ao/QF9UDcCKwaNP0KE9nrYl5Z9M2EOMHVI8rqUR5F1RSCfmLNnOaUQW4D
8kZYgW6dzG2eenG9xEWkEV5Erq5m4/tXWtQYPMoNgqz31qRdiUOhWcj+qqW6CSg0cqYgZyEEFiSP
eS72vpJ+srqItbgiKi49mdDjKjwOhbsF2ilktt3/yc/oCiUDzoOIuukBbK2f/pcD/TDjhiRI9AkV
jehk5zQKqmCGfVQFwivadxRqxCGp3zhhhmTJjTkMo+fIRpy/LWir1cfluNrRlv7UggG04ssBakWU
SppNc4l0+quRivjSADJmUnCweBjd8PuVxyJ46urgHg7kGf8L2wrW0qN/GfPP/xIZoIvVClgMeAbu
/+ThJ93fYCY+456i7ywkRBdaiXjJkk0Z0+6UJJlzL3vIYkgEwBnvbcooWystUxcPDbDKi26C0kUN
tAPTNTTaGmNwXVqAwPdP9l1YBJWnoyWhh0jgSeaSXnFiyuEulQl4ZNbQkJsXNNHdtk7ReCEDW4js
pQevSeb4HUTJggJwJhbuJlbHET3ikHzDOS71+krG4LXyoDhEpbX/53sWJ6RAsZY92enMkcIkn3+X
CPQwGBVj1nBt1ivUzqHdIyMJByJVuQiVvevWwhnEw8BqSw4cYGyaQNvaw+/OJ1ws631f3SzZHn4e
sqmMthZGdxZDFeBzG0OJk2+1EG1Fu40rm0OiNLjdqR3Tae20EGyCnOVOyaSavbBRrjkzrsvg4CJ0
ZuXFlM9fAWNOfnUtdqoNo74HbvgWjI4QjxMDBWuMFxUVIBd96QVO96yobp2YAqJHX+Hh8BjMUj0R
LqqH2pmovbw3KV2MKqZeYl+HovZ/OZ4i+fBkrh3E/2WFBK0emsPsK3T3u5uclqMtlw44Z3WbLa6Y
aCYQUQn5aKOFp5H1a9HTYqG8ihE9MEejvM0flwMSbH6D/wICBOMDMNb7JBW5wtrTYG/0P4UhttkT
5qUwHR9gazxxHb5Rib95OnS9N7Zc/76zatdqG74MKDyFol+vVj3GocS1QDbVQALV9/mV14V6jo2O
hX/j82rF9+1NwKB+IPmErJo2qOq5kUjyUneftzIpIZuPuLFFg8OgrVGxU0ZUbfNiPkdsyfKhuPgQ
4RRj0HijizXiDQW2Tmqq19aNLjpIm9WUyZieJyxpdvUM2Pn1XiI2WwuJM9Alnm6iPjD3ilnAKHjs
4bFvTHobH95sH6VOj/YS/J1w72iinTG6vE3CWaddo57wdfgW+9ORrTucjqJUFKCFeF81kW7WK1xd
eVic5/GUHF5Gp8W8shII1XtIioonoD1LN6mPBV4b4zxeXfROGlxOBbNyQ6OcXI7VuMrboOatuftf
E9H/pBVTrvFcYOkiKDJ9MKVKdbNClilG7/aD/OnyPXAtuSAP/frN1pn84Twae3yPzSrkIF5rdgc9
+pYbwVmaRPlF9fcs4wisND95qJcVkKE3niuVQsBSRYaqQ0Zkhy3S+kEP3Lrm7GnNL9SFUhI3BCtv
daBQqLxb9g8RhsdaFYJcoKASGX+aoZu7H3EEM9FwvwHk/MEBximlxz9elKs9Y5GcrePtJNwUN/Zo
NDgxVKfIIBDznMZ4OXFWwfLhi3ePWZSkDm97Ux/Jisu3ZL2xlzEKPHZGQs1vLam3mmbIWroPgj2F
VtPiX8P2BAsjxiCjE/Aeag4ljWZE9xb8MVAxisi69GaGB5jVZ9TKrEKSNrEhwz3cR/bhx9SQ+2Yb
lwAzlHJZhAEa3t/p+u0zVqpfkvJcpnFLiKxH4bnP95eYlUSP8ioDf6F6lYGJSDCz1zAz3ORUVKUu
E8DuoPRuraXtPQQmRS7W8yiJIo9Kg0NU0yojRh8et1GanjCwjHnzz0KCRRSOivtAf0wyZ9M7B49C
VsedsG0d1U0JqHlPf/I7yZOm7chXWwJTZ5AhcyGqb9mCYNq3FQRqxBuFz9kEe/uWLLqL7FI/Vlob
xJ84ZmYu3MS0ncuD+oWe771XKuQBNjT6v2XNoR9CcTnRzwbVTN99YbKkeqskOeVcB4rL6DIWbx03
Pl3vpZrbP21sZsphfQb1V3UD5XeroYQTG+W+p8IUdwHqntMJoKkZ1079Trysk3e2hJSx0HKjtoLN
oMuSRCsbANgZ09DG5Z7NOdFLeK/PxDP2SLifIHTdiP4kt0knf+DFAf3Y5hHgB49GLSzmclGR4pmP
PLdjL9vD/IZD0JxGbnTtWQXLmG+X5UAldpOjfPUOKrIDkRhCIWwQ/Wc8WPX40WWCUBxciQkley35
eBFzerSR3kK5MSUb+e8rYo+uuR7e2FbGT4f+dhEz9gRHFZzUEVux3Mg0ie6hJ4HQ/JnpDzClJQ0v
7qV5nmmCQKuFmMkpvSRjXg8GWAWEwDZo8bY049k/NNsPy4fMcIAY1BeSvgqQ3YB3Db1ImQF9gcMU
Cw1D72Rz9xOpbbXkNfwxeAbNga86n04HZPKVjyxzk2QuwYOYv0B0rZQa1LAPR+H0tFjJZ4VkXDs3
JH50oBfWSh507bdRZroq/WvBaFzLNQkmIM4JwffFn7fh5UrdmXsg3Ikhbf1BIgaNXTCxNPXrg6pO
o4Nqg66yIKT/mkoyDSl39u/CsFcinh/zIv1m0HVyAEXhVI7DU+q6fH/6mjjR1fLg5wam0nS+gCVk
IqAXFTgnXgP6o9J9HMZU9WXKaXuO+NRMyun/ZS8AIOlumh7m/ua/Xn5LMkkF8e7aJxn+Rnrj7y47
ONrmWYvr1ncCCMy6LSIIAjZAsPtkb1BmXeNymWQ3w0Kh8lkc5LQuh8spXr0vgI2BsOA8djHsxSD+
45Gq77YiYcC4ELbMAFlXpcnNPn9PNCNFfTlkIjmjXoY85n+GQEGfhzz1bYz/APzCiE2idT5WgHHO
0czLVw4etrlK+9Bax4axdWGpBLVwiO2wyrvGU/jEgGsLAq5LN+VnyMNJRHCzjkVHW3OVVr7yV4DJ
fEhHoyCer/rMKx9HSZj+zDUEFh/k7cbhjfeoTqGBxiGBzHR1vQWW80i0P0DehSAJg6OJ+0zP/VRd
SU+lQeWF9KKLSauT0MmfbHqMGMI+sDEHU9BI48fA+7rxmiMh9D88MbKMZODkMApC+jCpQyssee5f
4AIYTdAUp5tRXbt7REgNb8Q8bwgzDYd5f7jL5xTPaIWp9H6+ik4W6htVHefG+YNSxSzjK4BqiSSf
wqK39WjgIqTvzGI1XkPzJcdCq0a5cwQbKefwsPAIBpZEMUeYknXzfJJpWtg9ouT1CeL/dPCC/FLs
xrSg3Ue7Zxt3qgG5OGrnSAZVlvNK6dqAzrIJODKZajesMoShlJDXJcd7V9IziCfB1kDIGScC2S0/
YHkNPK8ix0hLullCMW25l+iD+VNEX0JKAquFp8jzcItUiZj9+kfPTHsCCAqwM9qnBIemBjV8R3V2
vzON4CMy/xM2fJjs6E8viu0P5STgqpxgCPA4C1UTgRsCrB1g6wIK7eyDjtiL7XiIaV0HAE4NSKV/
f0RHozBAA1YsgNjNsDVqUv/Hl4m15FKNOsnLYAiJkm2ye+b7vmDFTZhiBH4TQWqR/o9wfBIlBbfN
v6Vr9MUWygK18UEt6XJZodVc1oYNIZoBjg6JiSfCgclTlK9PvT6qrBw71P+ZLbf6xBJdT9GOE86v
GI4GLhdyFdxIgxzZZ3oNhQzc2kNzkhEq5gM5/KKOdCTwbAg44SRxwRvY5MZeKIC82EaacwwmoC2s
4BOHjSMMX3ODJicRinE4OCv7J8HImFHERoCNMOXNDkA1Hte20v/hz7IbHuEBlVlLM+fU6fpeOcSF
Wyt3qpNlsSWKHBoCY2QcwmG0PCg2Lw8t/I3x47y3UAeM41OfxmZYeyRqo5zrtvbJANWF2V/sLHCV
RRCuPcUP90vEobrnUnAQqHxk/i5dXCpsMhOJ3n+kaflO50zCF5QUSVV9kVQqBkIeGdVywbq/TowG
gx2J91o9/fXFY0JPjxTLaKEv3aYHmMDRSkCGBN4GopwQe3CISoUBTJcXBhp9d12UuAwnhxylCaly
V3/7uuYhcNnIZ2HRieblNHRuIV36FHPmOf2YRAbAqGcqBTxIHkPJUX2ZmCxtsvXdEF55oTgtTtPC
+9eli1YkHb4czqY/tLjSykbMKAdBd4rivEJT4GmbJyBqo34G0PlUGPyKDL/wU9sWBETlDeqGF8Vh
j/qrKb/JQA5JNsayQVTRYT8ULoG/AVqUBLb3yMN4usd4IjvdywYTpI2+B9J4WkT8UZmhR2ULoNA1
+NDVJp0jiAHANRaYfc03MJyFAmvvgPHJG63BVIXRV9Zvrfvs5ycMTeu3/LW5rE9gqHhM4NQ0pa9Y
BJTkiDvQLCu2+9ZGjVRmkOm+PCWCCl2Kuq3DgB/UzvAW62uBAHtXrDEj0ufhyElYizJGSii2X2hy
l447K/ElufOy2MrVlpdujbrDcu2b6aeb5A0w5tfNrIn5ZWHhOS8C0nVhzcMkwI3Me+KjRpG5F78n
uTsa/ARfiKLUJLil/NERukHehDtkO0PZ2WxGJemmGqVRYqH2JZNKxVk9S1IaKygb3Vs2cN+MaXll
4Uem0gBaJFIWc0m6DaIuyFVicDfaEDzaD0nXhpU/CgTIpfz5sFT3rpwiY6rlnOHza5b7lX2STcgV
pYp+i8wjIQh07pJ3iHLdWs1ScF6CH6fMZX9z4lT3EtR9gRh6OiSjq6PoIiBG7P8Nt/ABymOG7pp8
owfi70xWSlGwM/heyXxIUxyWu2zDEWxxFRzrcyt+qC82Jke+awy8hi1G+QeZrs7wMFsZTQJUzxcI
218Doc0LbTztA+I5/8YtBeoWZKQtkKkMlDZL3nYPQq3UzwCzq+xw1/yH+aAbuUfBB2OrvG8EX0br
iRZLrPbBjGSuHVcZ6UU+SEK6hpo9cgpLI1avKok8sJ4D5UShasgeWJwDfqT3nrZ7ax36xQa7roN5
vg9+rjEVWRttn6ZS9gUgv1w1VKoncVQRQ+YSCdZGlHNXfQhYVHVGh3RyPdOnacK4SSeZkmsjGWyP
oSyduMu+L0dfBRFdAFNx9Uq2DXjNjpud5hbCm80Jhw4q5a64ZJiZ9ZPi3ClfI72ZFuFFP+vabE1L
t5CUwLXun3X4fal/sYfH3bJbC7p3SlzXOy5YlIPzkivL7GrtUvY0kfFew7SVz1DqatOr50UWPt1F
MPJUDTuW75OuJNZEHHi+PVUysK6yAysLzsweIblaD9ix6TY+zfZxYNUX7fFqGlt+5z3ZAvhLG7t6
e7PChmRfadsVIKE/TjFhfZtOrVyh+P02oONOGgr09GyRRvcitn/3jPRo1JEaX+/VzAcBORfpDN9M
Oer1f8R/S8n/UMNclc//eNUzb3O66+VV1WejrKtgPItPlThTJvmYh3B5e5M8U/a4dM+FEk0nAFTg
XMVSzL161EkElfktXjW+8T3hvqFwwQNSRC0JS3z/gMQNgGq2eBTLKROaENyeCDWLljuyzqQgnWge
GNsEWtW0PIIOmZdlArd3hQ52/ZeAMyJJj/tYpeOIBzLaHDLPnd212vNQNyjYLACuQuDyUwScKtn+
b5LiZ2D8X0ibCzG9y1H8tBqr6FSfBno7L8FMa34j9qb/b2Jc460I9NPlcfMEHqSTtjTWznGST8Bz
iYeftalI2RZRe1ktDSeoimbwdJ8kmOi+lsYluLGGB3ylH5LWH+XYqEJBsKVPn1A+6DAgg+rhGSsr
p/d/uat8ZpRU2DlyfDWZGsX+GCSk2RwZO2+gWsPwR/qgU6on7U6JNILeUbVjXH7imIoeUzzbO42F
7ScWawBuQb0tE7ae7iQwKYY1cg+d4xejmKyPL/gD12Lr/bawvAHzESvelxm8qNOYPO+XQg/75FHz
YSSYFXRkNBGynUS3Fp3sjv+B9IwrDwPkpvq8fVhVZCSZmyXAEYxPdfrZ0NCLtH2N3ROHpfYXlgms
ILUwanQSER6+WM7OKj51H/K9URzp2OjWqoovMWJ7i7gFD3URclnuV6umJhZJGF3iblZWIxVPIB7Y
a6ZaM7Ds88li5P5pPMRLKqWpz/X+ubYpX8E+zxtyOs8EMJo/KQ/xP3DHiytJTfUztPARBEu50Iup
JLFwBogKBne04Flu0hhu4fx54v0GwNQZN3wWZnuoZNnhqkmtN0U/ud3dJChy0nWFXa8O4LoBoUnZ
FeM4L9jyLIihYA2HcbQMMu4OcQwRkXBACb/sxmoNFrL2RKQdoAEAvZ54H+pzmWEMUjq20eb7Knix
jbYPl1JTnMSWGCj+bb4c0pfff6ZwdI1bf2abPu6uDnii7F43RfKu2pEYvm1EmNVJnY9ycX5F7k46
AiJL4ncXaAcL27qxnefssKZGngjel4YDY46MlpL/mVilp/tqu06yMXJ7kOkFgMr2bYHrQkwc4ZJw
Ym70ly6wLtK+SKPxRyePME5NM6pw+zuCmw216cZwpiwE0ATZuoz9O1mPzEOt5SHSukTgLREv9Eud
pZ/U/S+K8mZ9WZr7yFy949BXywBr2jI11tGEKGiz6yX0vzn0UjSRcwxiqHBczudpTOhShBEf+pUc
aHxMXpQqTHnX+3sFaKLFXL8VRsVnWtyGU8XdjUMPHXIJuLd2tVMAkOQ2M8C2s+j3AQ0fFISsHZ/2
1s/MqSDUIul6HAQ5oyzgy+IPmIviq4EpQUB49oi/DPsPLWjSNasthxSKWfdla1aDEqjjZbqOKOhf
GcUlfevC6sOfdr7hhSEkU0+opfU/ILk7lal5xa4+4u6nwep/Fqc8I1QJPpRRlis6EiV4a37TBiQH
xLNoNReqMkEpLyH6eV0ObdTjeQEp0ljE5wXy4Abhju3Sliadt7TqyUJB1j8HV3MTFRczBTjVeVq6
3ZQmdPYRdT5b5xlIPA9VpoewezYXaMcFASLbq3aiiCwZsyXf2iEThn0tu59L1WeBg6+gYIVrhRBr
0ccUyD/OoyEm6Ta7yzPfFVyRepWmWSmXGgXstRYK+/d8IoAJSAInqRN9uFUnm1e0VWtagQZifBeg
FxKh5UvTZ7kdizOGF4LDoHyCoNsC0BPMPL1cLJQNdxfjvLfxgU5Q7Pfc3jJpYJWrRUcYtt/TEX5J
UfX0HKWiyL7TuEnf7NijtOmXSATYuPNo6iRbuS0bwW+K9eosHQcNYB0sMj9tw553thLMDD/VWK5R
/uJGJ4cGB+jJV67z1CdGMciApioWMskeOmGujaAlLa5oaWpi1j83fTZIu5Rq1D/kIIS9zgycZldo
ICZcw5d33qnUKF7MkA7FCqrZPF/bzts+yrDpBkf3RL7XF+gf5eM5/JOUJqEdxdVL/+Cw2bK/cJ5j
SR3f4xVhiUCiKi7XeR4pPIhYBVa0YaiSnlA4xVOB41Sl3gW5VWvxbct4/oaBToQ1YYuF13Liarj9
C6JCI7grzzGGMEv8vLIcRncyx6Ncurd1uN4p5v3U28Vf5P4X6sYu2rbEGpVxtqqC/9y303CSEcdj
fHPuGOfFV45pz31P7Ye98I3Tz2QZw4vMpBhGeBI8+q3L1FM4fw0qYQJLYEuxqy6aYq2jAG/l52CX
LjjT4EFYcyM6QrOPt9GGGuKiCIrfW57hpN/uoUU569QfU5B2KioGnVNbJ9CSF0YyqpJ512x1LDt2
Gw6sqh+VGcsWk9hAQ4U/i1eKhHSLwwxMB0H80puW6Zo6kvEllLzFveV9AgAXBqQc4gruMsub1ZkH
UACttn3p5DKL6Vetn9fX3znhk2TZ7p11ceIuDCk61RY187BUC43XILnTJThTpoh97pI8EkF0Gzz9
cy9ADRTg8IQ8R9fCfbqt7KkACgVQ7v9S+yP9W3ZWHRLxcFwCUhvOrnWeHZMNIpBxrCI3m4kRqwnM
dd54gb5MgeQaYZfuSQQ+/A8nTi7purgLf/ynYuD4gaPRY505IE4tHFBGGMerWfOtAvDYeSndNBm1
nADkOtOFZK4wE//J4AuiuYxVjA7KgNlOZ/LNx2SPmN6Zd/x5wzU+0lKk2Kd1Brf+7DbJokpLbOHz
hXL5aaeWIwVqM2WOzAP3uqtn35fqx/GKVf268YRHGdwyA1ezPfp8BpfBUoUy62OqHD0WqYe5bmks
gxVoGe62EY5fMomYQjLK5OV3GZSbR3lcTvtNyZlomyB0OoDx4KZhjAoTrCOYGLK+faDdjOB/hRch
4kBIi1F16TKhWCTt52zjv7DofqPjQK9O742eIl+fajv7KjdjX492626BuhAdiNrEyunVwxPW7obX
7gnZHm9OxCTdXW55JppAJsJBLebKPn57CYQIVi5tLHmmY/NrW6e/Pqf6tZfJ/JA1ec5VduLPkZ5y
W3Uz8s+wYnFTqp+accy+Pn9wU6mR9bi1CgP8ZhbDtloPgL56dX5wuze5gWpdc4wg8VTUoYkZUt/B
kZ8UMfxane/EuZMJ7O3v6v+qcW5j5/a1dLWjZwRV23L/VejpzmSD5V6aS81rq7xpAwZDUMSe/YfG
NghGkpNK5yzTpoPSCsx/MiB0EaqFRWLRsGv0EQK3aow3dlCIydG7sK5F/XzK+Ulc4o7KTB1EC64y
H66M+nWQvCf6Gpg86clnALfi6URnnve2o/63QREDPu7pro46ZmcLq81L2RJsGhiGlx3yRbGIiblO
I39E44ARiKHX5iOTjZlGlu00q/FA1o/+wfq2LL+QpkxKcXTRgTJqaYMvf4bAHs4f85P2Cpz2/+ap
WHTDNg/bpDAKGVPut00sxyBkKah8mvQEQOH3uVOOe5FLYaVG7AdEgqMUlMa3JQdVZsLiDn8gQUgr
JY/e/UChCUq/bok/Leu667XnFx52wlvXxQrO/IYhnmCWOHmFKbY53UKDPWjADICYNb+QyPCyR5L5
D58TC5hWR/1qMegxo64piLmyjbxZABzWeYzc0ClKBAj7NtmWEq0HvwNo0zobo2rmf4z2iJ79StKr
aIgpX3v8BqOBQPtE48EYjVXO3s23ApEUrC+ir4lI1Bs11q95f7fAsa1r+DfFwpQW3KoRJC4zKTnW
H3MTG/vD028zFEIWvAbf/narPhumkntpgvm3Dc7VmYSwww+VNpP+m40JYovF7LdpJ1prbsKa8/oB
WHilEeonDbYiYI4+XyfJtqCcYy74v1Vs6F4QgNpOrlZWlIpgghRBAPbhacBnP65/BtrGRQ5JclID
EJpuAHPd24RixQ0anddEeA+/O2Imogr2g78x5h/efG/eYgYmHAzO7nn9YbSq5FIUHLBd1CPu9oIO
zRHN5zmO5S3eWXmAkiRQmmwz/vnwKSnYUZjUdNe84P7BJdXU3kqjF+jf4D/Dn2SU2qwRK6BydCp6
CfY86oqVU+lg/U6nTQ5LgbOlXf9boXb0botkGgo8f3dSPYcbVSjm1nU+goj3IMuTJLFbfY+zQd7j
ncHPWdarBqqva4u+QECWibJINbn/eo1KDx7AihPoLTrchJ2DbMUABpibGQbQzDNK12E0OVinJP1H
Acw0gQ7HOZqDq3zIOIA/MQuWF4QYpg/W1fD9UZdh1ageTEEJWhKMtjBcxO1i6M7FqxFIeQm3IE3p
/yh3YEyr1+5K23WmtzLqjBxQCeqqrLfaar9Trt0PYmaR8/rDhI425sN2qjZ+HYZXCRLkL9uHa3Cx
ICo9eZkOGkpJGCL+F0k1Y3oZQXq3byVqu5L7inamrOZR/eIF+elMLv9N8sEP2recDg6aeqtkWYmX
/3Gcpfpb+A33sMyRwkvijy0XoejZY24aEy+WuaTdpyN9jgomrnqt+eSGH9VV4NkKARSHgdeT9k1m
F9NeXqrXDeKEy7DD2WZCutOjB8oSA+uhyMIRJFFRVPE79dZPfpXxmZu/dFSvl4KqRjg4IeFX5s/t
jjag2GQ7ERbu5ZWMCQKeHU+23AD8PFUAi3Y8BZi0uLbr+q2EdpJ7nUfbPOFG1cNAe7srrtH2OO1e
84Gjhpn8mbmheGDbbg01FULOqQP/VzfUdZjv5D4evLDQT6eUlFztUKOfaQdQQKwe0iwtYN1S4QIT
121OmCoxgLc62P8tHqcxiEBNMnj82aLDfgdTTP6cPBNnMKnKViaMmF4JzAO0GHhiO3RiL9s2adqf
vN5St793Y5lMg6i3oz3YGUdIqx9hdoKGoc09d329KyYKhHJ6W0WVyil5CL11uGeAvSHCEo3gpdVI
5MYuq+E0xOmuys3flAWl60ilYNxhgPGBt1xGLblK4KUqqEyF+PuxduP+OKBHOIW/qFl+gqwm/rHm
oWalCBjc8y98Ok/jZNUgu7Uogv8cFI5RTYFV8KMc/o889HGBoyPqebeH29gwrM7VYf8IbNfZMwMf
VgxBTSW9/dZmUNpHMKaZkSDJ9f3hys1EaKxKvGKnPT7zh+++u4Wq1EDW+ftYh+Hi6s+NY6TzdbWR
ht69bbWdnIJKvoq7/20IJT6J59SV96FTXeCtAoJpdKUf+2gN+YjJC7i8+GD2lZxUta1mrwBbL3gO
eOKJ4p6qn1bMHbSnVlKbLwohLJfaUhR8iWeOGpx7Tj3zRMamFVbHsbPeV55fi9Z7QvTkHWmUCMEq
1BGnstSR64RwXmSlx1xSUHbcHbBxV1RvqPpIVj3cQHpLRB79Kf7F9O/YpkCbbQWCpJ/6rdEaDPrG
2WPX2YuyRIEVu81RonYAb9WZJrmZs3Y8hHaHDpAcjKILz8BwtqSFUomqrIG9v4wFNiKl/CHXnbCS
+HEawxM2qJZJ8FhjqaHWhuU2qWlbRnn9RCXHYiCPk83t1X0UsdcOqLrby0F+POMqZrh5DR7BvhLl
c24VuE/CgJfhy98n+8xhcZQpKH5yx3GtQIaQNBFkjfpTZnzc4T9+4+BBxehAvqedG+dSPCYgLJE0
+uOULI2Htfsw9PlBvaGf5YfS+RpJWFKW75pEQtSmpwf3ZX3HOkDM4D+szfDw53DX3TBk5Z4YYTT8
skzruiQ4QOavb8WKEQ1SYLhCvMvBDUdJOivSjCiUNyUOvaxP798Q+hgZE8zz4WqEOwTAOb1Q3OhW
zTDEdlFLW/BlL91fXqUE2eIuoJsIKnZDh2+bIM78NlvMkDvgnfUY4wk63Ts2Zha0zj21AP/5PVjO
h/Qj0i74T6oqYED3n2wLoqmuSV13WBlU2I85V0wSPtNvlWbWCnThHmremhtJTDSmNh9SDrXv0ET/
8E21/JyEl1lEmkIaOBgC3mVvNnUN0wy7tudb52I7Gqts9S2Ody0uqVnud3VacahhEnRlIYWKQyXO
LyHWINCP5FbrTKR9XreHXTsd+KfFcynn7Gn072nSYECzuzsuWv6D9YPP2fWbPsnAa20u5pIv2n+f
DZ2hBeYpFgh3Rrh+Zegpzw9o1Q8M7Hhv/elOYK6Zv/mi7TyjEsscoLFyvBL1vGKLAqo96sr+FKeY
uw18ubWvgemrUrVSd/maBrFqDJYryfXNam5bK/vYVrRzt2ObDNhPs4QnZTM4HR/AJRlyy+A38f2r
sFP1FTiHbdByS3I8HTnesJmH5Iwzu/u9n6uRe619k/+bMYopN+9XU1UfECqGeG4jew1Tqd4EAth/
gddJFS3YnA7Y1PYrYUnuxN5egTtuQD7d04Vuby87NyvcnjuvSGewrs59J8IM4aRQ4rQY64EGnack
ghJ7xt7ROPMb6f7OO6VZgwzI1/5fh2Jg9e9iwbYJu2Oec6kwQn0tqd3lQBV7ljtZvTEOFmYXILFc
KbqmyM2RG2FwO8hEIbvBOFVEA5Fq/mWaMjs6oCk0ujblhCh6uSPzgloPaJXtGRkzc4CSNI9WHyEK
msft3a9T4uBh4WHK9FsiG9cdw0emVoJx9gQ21OnFSrXrMZUwS949vZS6TgBqsMCxjPAy1LfnR1+C
TEcoKw7Mp9LH8OGu5zfW+lwFZo3Nqz/7114ahugSaVk7bRLWX2G+hivSjoYpGSHuucYKS4rBL6f1
yN/H1vqGaVRxvSqvgzyOylHdheiQ+VErIL39vPMkRqHymjR7tthulS45v4XaiKsw4ZkM0Am5H2j3
FWMUjSF53Xnilz69UTHjGGl47tPYlFdWTRcazHwkCHcj4KgGajeLM7afTO/W3wC6tYoqRKKcerMX
9SjEEyUBDyiYUTg48G4GI/+M/GACG3Yn/HsaIiJiqZ3YyZZHL82Zxcf1jHSSTevPWEl4PiN/kfS4
AV4+cJdXpkwabOqUMX2gCMnomWmoY68l+LSsh5+iSMTwk8byPIFjyDhd0uWmt8iYmr4n+38wyBM7
64suxC7LpbGKa1gNL0vbIoC49hxOJTFRrSlcvdJtzgDuF+0qn7nqbiJtRdqMs3b33ereR2fE5p66
mvzBRSeo5aG4yqp0udlos5oVEgHL2iMDvlODizBiTXaCURYsXdYcMHIy0NyyV1GSz5yrogH7FfNg
5bE7PifBoQN2O5tFnbdLrVIO/OePf/bbQ5itmPYnBaDgxf3MiZ2/+yt0lzdFc8y8wGaeSgIFzFOi
vXG7Tv3NCxRxlMHaUMdakmJEb8xnWLCFokJERNbCiHk7D39+waR9JsmzPjupUlZEx3WaRtFYfYAw
gMYUF1AP9xYI8EtCgYou2nsgcR5kdZC5cy5MI0HxJP/qB/ipbFqg44InDBFKrU+6cdmU3iKajL46
5JnJ0DzmsQa/8481iEUaPV+d/8V/s3ilqq7Uirf33b9iPdiLI145HPrakBqOenZb7fxZBq6mdeXN
KnJjpNiqnzkNeNY4+hOvk7H3hPdI6IcDV6tYdlgdvBZc7HWyWTm/LwvowseJIhgJkoSCGPoK4vdx
VaaLBzJ0i1vQnkdzErBOMweAlLsiljan2XPteAs1Gu2XzXLPjNr7JzZQwlspeyWGut+LTsUd1yuM
N+hDoBa1R5bV+JU4jRvR7D7mOfSdLNhM1LpfR/f1jK1CrgMYI2tG19/GzBE5NuH2fE3iAMfQ6CPe
/dhsjLroyfhyDOOMMWDxVPlcZzt5wIiPO8KOYSpFupKe3MwcQn54g+845a9gonks2uSoFsZGZ3ON
UXDBE2q1jPC2CUgkDrT8kShy6J7gDrnnHu5UDrvf6KHccp6PUy33pMw3EptGuFQAsHQZrgxTJLRT
5766ohNwbq40aI4Es2MNEOU20mh/CJPyHKhUaixEzpKNST1Lrp2nj4ZzO7wRpUabxXWTl624DXO4
qO/U7Nr7Lh15D47VUguiMhtdCTGevM9JCFRjrbllrwXs3dVCsYr4OaOSTgsbX3nz4esmnWdq3BM2
kdTa4R2aMYTg65xwd44Ct3ueQkkAYsETz3QRJuEKxOvQ+gj3KUPL3x3FHQHWYIUCe1bPy/vo0WE+
KTOF4s+Pp2zFguNwdeSHVoRUXfEslOhNpJj0kBLBgIosMbiOM6fmCL624OHObpfhKva6OCK+28St
H4YQP9W8Ozwp/XhlV78/c74txSRi2OWZ33cu5VRk95vFyVMxZETjQNFF6gC8MT51sbYuQFet7yWm
jnrXSeqZayyHX5nuTx7J3HUj8qIKzSsX87LwUvvZSqyjup/15XHxyPuk8pSllLmlYyD8Q72nxby7
F6A9esZ1QBCXObXZRll/YD8yVajjJizaFUSQXPlBO0Gn8DJdBQj9x/ggC3ospQ2WoKrd7ZwKouRL
ToXBfFdpNXiXtfhI0fYBZdL5UXpbVVsPsXE5nV/K2WPk+EYxA+IvQwXHIZd3VR3Zi5RUv2q8wB41
xEzOhzLm5xeZ0/eJjG55TxmWF26Ha6I2EzVqjK9lkz+HXTpyPbMUc5pRRClwxn0/IweiMgel++sD
sZQob5YQb4RKuz33c7JrjdiQAlD3qx7IyH7GaysFm33IlHwwTaFLv3UcIMhSOa0EYzqzI9Fh+tS7
Ke9FyVdoDBnOQbaZZKrEhf8nKHmIm7PXDD751+hrQvxmqLR4BZ6ElpMOQA32xx/UYdZk63cEaXrC
mywP1SnEQ6kGoFDfTEtFh7nPOZUQfT+h6lq2gAlWw+RYo34dd8xbdvkXtk9NTROVVMP+OjKpbusq
csA/2c3iuG+o5QTuIIPP8sky1hbhfbLW38EcWGDbpE6qTNouwQhHwl2MmOMiRhYJ8xeybHMAHQV8
GYQNb3cbPoKbT+ZnHfTwONfuBgoGPZUonmFr3DAlYU6HF8MUHlvmXTYyvtTNzrPIWWb4kGMbxZKe
RUBghyNx92nghDHvIAvgitjzIf+qMWIiRU4ReDZb/cqbkG2NtIXZMcN4I4NInlTEbGQ+6J7xMnpy
yaK6OyufnfvgG+ENW5eYohm9hAB7wCxsMOH5N+vMP5SL9AT7859VBO1Prqlylt6pLxUQxCn44WxP
71dUAHGIgOWYaiKqGoUMfAoeaG6AHfuQNYKsPEzmTfXYgwFZG1mlMe2HERWVbQEg+qZogLTkVrzY
GDw8hSySI7VZPd4qCbN2KXsETY5THYTwkeLzhyYLiIyYilOv4ooJ/BeIEq1A6B3pskaJmGG51SEF
BXNkrwOCDlMqHKnM4NB8ldAlciw22j7Ff6upAtS6nTk8NB9zHXQbWy4bZhEEyq2rdxqV1TSXDqta
CcZ8hWNDXNrofrGExsxJYsz12xyy1lrTyAkrbRY9OjHs999/gxodssVLiwPQquYby9QOxhK8CS1K
Myn1QL9YB9BMa7MJHeF03I7fO65bCukTCvqe1GnnMrcOzGWpPuhl7P7EGthkOJETm3eZU3L5I+UJ
wCdgCvR1lsZaJT4FSv33kEYujpDfl/9WNVkOPr8XSpCQQCGO51P6vYwoswpEftc010ghjJu//ARB
kLT091fwRldrvNm4OseO0WUKdr9bjgyI+TfmNYGdPuahvUiqKtypN7pWoILwcK0bb3IwbbLWrga+
zPGcOTsB5ZuK/mYpqHvXjWwDkV9QqVis7xfFwxk2Orxy8wOK2bNjNV/zjva2aNIsJafReg5/pRbp
hJbuJCI0DFLFTRR5LZoIZdzhoUwt7xe02W3WoeV51IsHMZNPdNHddohC3nH12OrLtPwoS9L7cn9L
DWRwNzUnkYN+Bix65I4kl5JYsDlsQvgoQanh/J88gxhRl4eNX2Iy5/jg7cBTY7ktiALyHVwgziSg
dnP3rN6CBW6pp02M8/BgIKQCOWlKa7Lj18u1I1dSudbQ0YCOWebq6uxGXWFSOH8zHwjPwP9bllzt
ryxoFUoXWJaYskiGpIGRz508JJOFzwNTWToXI1+wQkn97rOH68KQnS1IJyyia0plriuUrVM12PoQ
juUe8OIyy9sg2tVrLUjnQFRMSqZMG1qYGzkqSZ0Rrdj1ZsX/Na3ETVmv8oFIHibkVC59MpZCcKuZ
xU9tyyllJYzNUkJf9sbl4sRI7NgEufhW5CpLpNsq+xwV8nrcYN3KNfR87PWikECcHVAqoZL2TrNV
wbDE2SPoDQpkUMwI20T6b2eVMpgmWC1rtPR9Y7B+nJNbaBLzqDWkPmW2Bd+DgWZY6E3G7TzcbX94
1i6NER6C1LS8a79lfeVDHB+w9Q8CAyl0ci6rGPm97TRVxjDPe2qUckdaQWxDDWAFZxBifpo5agKg
4uyTVn/Ip/PlqX7AbCDfZxFqOPryXNfk7c/7+Eg4vctECelVaTo8emPd1dvVLtHhlcWoTueY2+g8
zha2zq8FTa/jOs2PV2PbIy6LTbZpQ/cOkJ9nTE5+JyvnhzgJNEBKWay3yZncJ2IRGng34dZ1pQB0
xAaz7kvZOqLjk3ozkli2TILtXe0IrNqCRg27seG3sTg0p7+lXulv4LWo9ZZNFSj0/RTn7qvnTQ9b
9RknepmDJqODNWfIFhZezDJdGzN0E6aucnCEWOdJlPyxjLV4PWGcgx3S3MpvgwWRGDOWoJqDHMj9
BmQ6ulN3jBRlctsfoN5J0bi5XclCt3tvzMnF04d+aaGeGJkaiIkymKNgUsWMdLtuI+sLRZnrxvhF
Y0CAiACYOiz3dgWnHVCkoEeQZKNoJIXKf0mcvDKOwnKf8cjqJ3XNk5VAwToFIentcLINxJTDWnX1
Bm+cM1rN0NEsjTAeZvX69h9mFdfFAXjrbErblYyuUVSRM53jA+cCNHM2ZdaME3/MjEUjUk/jq+En
s2K/uRDj4iJPxUieXJJd/8VPmt6C0o1YNz/dEq4B+oJYXXz2NPsWKFmZzj5f3iq3p/G3G3McoroL
dBNqwSCOuc62dMbkR+CLWipcyfRrc1Wt1mogaMcKf67/aENHMLhiGmpm6yWvv5cUY5x6kSCbACWR
mt1UXscY+eDS0pisZr4einBJ6o3bisuwLkJ1YUI/gXAFPM1+jJcBlMaq5PeXL0vWJ9k0FaTTMAEk
maZ2gRXXV9uDHfOwdhKAt51SiXXRJpCc0VuRzMl9icNaB3A4to58yojxlJCdvUs53AkkUT5Ax3bK
0OGqWxj9E8UgZI8F5vRHf7iehOqPuUnuT1XZjtF1bZKiu860izG9H0xCPPeCZI7nQEa2fQpr7sfV
oML0JqJ3D+m31al+pZ/2t5i/xM7pR2AKs5RjwVBOod+192xlMhIU8BhCJlejGRXMi/6ICkG7kQEs
E/LLo6C1MBfCl9Y40ZWFZXCKXNJBy85r/IjqAwxhYLydRv5Ps2QjD/Fp0Bx7KUzUsH4Gh591jIJD
DcZutQgNUgAdPDL8j60GC958aCEa83JkvAr5h5/NnYtwbRCe5HA7rEm3pFYyo9QSBsBywR1Y2HuF
iT2u5gqcPczDNtcUrHs3VcCj1/I9hO2mgbjwiNsW8VrQJ2R+NQcgQKDF/7ekhD1gUUKVGqJKLFmR
plQKwSBqahz05dv8Tq8sYzA9fNuFGS6agOAdWHrVL2jl8kHB5k1kizIcyh0MPeqLSyLMhBev/A9g
2prx8VKoqrp/ruIOh1tHL3f9+63LvJ8ZGDw+9XNfxQBrIBzAqAefkQgFkCAtswLrInoWUy85HYIo
9q8NzlyIj24XXGooJAapE839mwMV9T+HSOums7eFXUynL/7HFTMmImjAsV47gl1VJ12J/UDysTCK
9qOxZzJMbOvM5DiYkm29WMNz9H/wFEvpHt+Uq2DAzaUy8PcbaxOJDFyHaGl9PySvFVfLvDElZLIf
abPWKUUbmOeB4QS98pU0AR/IEUplnl2/X3R65Ki5wujRIYrioELJHKOka5ORIWGUC4/X/RcEXsPW
CNbFrbd3lxdrPREqoGHZh6vdS5zy0BbAkL17rBZluVJ/ggmGwlegZ1+ASjLOi2lyhCU43KbOSUHb
WXy0vJ1cC94zl1UreDxxXc+qrE/ySfrJP1NJTa/wMg5AYSytxXmK6pwKvZ39KyNkenVlfOkoYkG7
heD9/fy4Jlw+g/YoJFgODFdizqvF4wftKeNJFnTWg2WDjUymOUxzjzCQdwcDcr8cNNcLVdoV3K27
sn+fl5Axtb1uO/JqRJ9TY2Z6qYSDVP3pYfxs1fhpB9BtXHkT0K6zFidPCWuAoFVbOvH2HPcnQm9C
7fQoHhyqxd6btqjVP0ofzhESVUJNqybd1onYi5waHtyTNr6psSAHv9b5pR9ZV48fqihvFo2I4/9I
qOaHL5XAWQ6Sh7Fd8OrBHd3JFoB0VzqisI7y2S32HgYQCufz8wltdohJixFlEKUPL5h3P5jUbTpc
cayuKu9QtI+QBnmbMJKz5SkCrSag+leZqYF8coifsHe8qb71K7sA2Ovw5rDYRXbE4bCIfbk9qgBj
A7aMHySMrpJS/yyJLuutsjO8osa31gzUx+6AUcl1cVAQDmdQj7vZT+PG88lOKxyWswihJmt3MuMy
8FPGQqdN5bE+ph2bAxWstjoMdRg2F4tewLmRVb5cvc12JbtHndH7H2AH50WSW4HJ/6p95gZ1rAnD
+2C6spvpJbZHZqHwnX4f1GeXYU+0+rEom/oz1wrEx9MLkYSlNEGiWbudyKBeNQ5/jLPir3EBTjFQ
iPCHHVu66SX4B7ujket/x2gJv3ZZ2r1qYIqJe2QgRrNk4v4VWVxLTqGKa1SoKy6cXfDsNg8gaXGS
KuaigkPKZFGBvWxe/iS3ZPd1y/8c2hN1n/VoeAGLrMguZUApAtZNUBOpxTx1jpgC0RRcBBnUsuDq
9+fXZ/dPrgqVWSqOBWUv0rrezCjNBe5YDLoO+hlmwvIE8KoOcT10QkSFRymGLjSb8PRX2U3jNuIy
C5M6JYsPFSgFMU2bdo1279IEQWkC+XF4H+CRjHyMlUJQzBc6h3w+6+49EiJvq48sjD1cP12+IMCN
zNusrpd4f9CCs17EsnfjIj69W8YQrDTCEXMPC6FVgfm8NILSL/fRCRlfzfy6CTAp+6MkVK4Y66jb
9fTgFJrTHuZtreRPLfRrGDg8Ci/HW5XH3jLV8AXqnl3X630c7L0WTV9meGgp0EelYCyZwl1XcuSg
4NSnz/97HdOHssfLWKHz4y5s8ZrLaixogWxyLjWJwrCwMk0qKXr9t/A1/qrQNNidQ10HBBL4iIYx
xTZEAHLwpxxwkGosLQUuuwyDgOOkJBws7AiNWsyze5cqqPQM56Tx1VKiiJmCdR3fEV61H3ZUhtHs
gkky5jmMyEetiLcCQLkxzKaTLrww31FePmRaal2h5RZhdxcrXHGvk7e5VWOxQw5EL7VdbfXJMO4s
sf2rOfCQdgj9/h8vYEy6Kg3Yhx9icGZckQqVYOnZZpTI64Bfzbsow72UJxleFkxeOsP8l8NC4mDA
wvEsW1fLuLyZmOsaDxr3a2GpKJ6lPf1Q3QDT4p4KIyh+rKcllthI5SsoskPv6Ic3+JW80CVCed5P
8uURf5Six744ZVNnxdehqkQT8EAaoXJ6IBiXvE98GPTiGW6TM+4Gp3MEZ8gt0snN6EBE3ijg8Y14
6YKt9XtMCMeS1239twA/mrV5qRUzEtX+74ttM5die09tTw+eqCmrfBVSzxef4nCt1BYd7PaBMht/
pzHguG/3lpVdESDRhEl081wuxmQtedCnyh6g8HuEnzL1BHTU0dp03kVwUGN0bcQHe0zDyOs9ByTJ
Nop1q7Jl6PbXaBO62lnejNhAax+JcmCB4FMrgGi7n7OnDn1/92pnNwK4bWvefvOHLzVrP6whEqbe
s2O017KEit5KkXbHXpyIxEoqlvJ76ctAuSrm218/+jc6oaRU5Ewt+vkDNvQkNOF+nvQyp/BnKgIK
gVE7L7u8FJNFoI6mE7EtLTvke0pClw2opq9dQRJ6PxyHi9iCYx4U5FMqvd7g+pg0C+ivmZWCBfCE
RFtde+TxpzU3iAfFIaFPugn46stmzBFCCUamBs6r1ebWoZwA1Xi1Kq5/OdL/HnBgNjLA84vUPMp6
mAOZjE1kXbKGixyIb4IADbvU+Bxv5WWWam2WSxdGUFFSI4z4GB+EFOtUlociIIRc29EW4NMnXzyW
U1wWy9MZtRpo9LAeFCwjcIT9APErxKkT3XWAVK1WzofhQ2sjM05gh4zYbr6bOYBTewkYmqiCzRvb
TOgqnts8mY1O1b1avQCtA+BW4ktKGNgn4Za4qL5Oc2q+3/30EVcxxcwQSIRON8M7/26ops7pc7Sq
MmCSBdldsVog0DsYQt1Ak8JUSOWiIvmWW5CSOjdYRSWDhfL7IIYWjA0YJjeVauGa6+Mx2MRDYW4H
5adVDaqzOMjOilBhvOWUu0LA4kOq9/6YC6o9rwdoCszSPrOWQmQ2EFnCdwBlVqdV3lY3KkTUiFaL
YSEa2N0oSnFDey4VLtWJidcE78ur2UjGwUBTtlWTj89u1WGXbHgLOTxkW8IDayLQX06VdZKy8K+7
mDChmg+ekirrUaepeYPrBchQXcy38rPM/a8TCzi6sjlC8wUQLR3W8TSsdSJRTp4659Tj75paWG9E
mY0MJVy8HIMPfDSdF/pxL7txcBnGweCvZ9iF2GkoaUPmNwhaOQhiVlkuWMJzdeKyOZlrAGQCGeQh
8ukZhKuzpbM/jhIV57hdu64BGpUUyX7bSm3vMp/b9jfcfjF1I0cPzKe9Ad88MII+m2izueLL+9Ea
UCGpGcONs88pIzIxiV5jZY13TafT3uSiIWE57YLWeqhWqmMYtWA8WtQZ6H49ZEAjlfLEFDKknZ0v
Utkd62AJ+jnmFSfIM95tGo6NIMyZ8BRvQXyrd76v9tiErkAQyKRfK26lH7F1FgGlgzD3K9mBhrQt
C6yg9s711PRXWUjmt8qUMzNmKYBxSPnaX7/O6gC/rlwDydj0ot+L8cckd+oQ2K/l8oXuYzUvVP8l
wJ7JInjROZpRCn0RxISMSNoNzPrCZX6Q2NEqMwfFbVQJLtp/SyC5Tp33wHD18axSJ4HhU3Bv0CuS
JVZhSNCBKxi2rcOXHq6wmT79HsYL9MpfvKUqQIe7kf0K4oBWZcVnnAsWOPph+DU2inNnwOWovs5N
CTH2BRGDLsxRSK/0SMMRO2yJr79OtsS9e4TDNHz/4OvVb9Wxuki5udQGDCOixJ0Bh+LX1N9Agozb
QYuJvjj7ivsiGgU2erokd5CGGSabHcxoFCFgIuHz9j85Sqbqo/msxvsXamtxSrrmMv9ocUKa6Z3t
RoncCHvS1RxMKIVZg44D823Fa5aFcd34SH5TPFX/Xe9N2vMRj+jwUObmga3sYYncA1r3M9BvFTAg
16dcOLj9zp0mb6yY0Ezb2Q3U/Lzry4YVhDDmYKpAcg0eMaK7DTfIGBRop5qVzQPda8jPKG2fe9j9
l9PpjphMpCSuNlyUdF2NuIs9hHyPhKMf51R9xFfzLYfrPq8ZeA114oLWCfK7IBXddI94I325mBr2
OyJTKjgLilOwj1k0QUSVViYLBmH2Od4gIEkGqW77j9EiquZxd01tCaFqAjEeRFtRuxvw8uHbaJdW
JNZwjxBgn679u2nT7Wv2QtIHP1eKHpsqVDbTXTJPekdBSYnSAxQPsGVOjth41lMm3wnbH+NmclYY
TFYmm2VOaCxwj6YqeVsT34q9qp1RDj39/jK+mCdHATh3q6G02ixpfJKppsl4RCe0/QNJuQcpls0t
oCTXgp+5Gdtt51J8q/YSDZT2hxChdqjFlp+iiftnxTh5tvGfhkNmm4k7Ei0hoD6sYAF7OC6pE4Fs
q+cBawuwKgSLBDyXTgb1+KcswOe0IminCA+yHboy4VfS+BG7Z/uqBni2SCtjrX2YRoEvdhT96ecm
SThsztG194iwx/7KQq1Qm4jsKk5g16XaT17JGVmBE5FOFfjrN5TBMx5PD0oVG2Za3jL6dMC+pyH/
UTGdWDqzjVkhpA7YCl21gIjPWRUvmD1G0ZAQpY1K1Tl6kETU7fBe1F27e7CisILY4vhV9+OCje6N
kK2T7R6y958LdLaiD5y5CRSgS+HbkWA/2ObmdlrleeLbNZksuPmY7v7tK5CFuCiUDlmdNVzriESr
Aw+oTx+Itpq/UBU3q8ZuTRray8DOIAs26Cz4RWtLrLQQ/PD4jkaINBAL44k2er9005rkMTXx4Mj6
lDi/yBBu4QzM/+csKmiUj+P3NE+sHnoG81kYLDWEfMPrL3DFFlaqk4FGeySqa7aQUcnmCAwAV28y
FdXk0Dy9w98zhzb2rkF+S710GC1ryoWjwb4n5WCRncV/Y0GJKgjYxr0gngiZvAo5oaoY+nPTDsTr
jJBVj4vjLD62uRzBu/n4QcMvQHCVhTJZJAyHF/WsIPrEOkjoBJW7ZTRcXzAmwiiU4RrUt6RcbXdh
wjO4ZuLgmuGYJH+74wap4O+tugFLsDnhWqL1DmIEvPI5CNcSM9gkTHlloO5/rM1C76WHt5eejAhs
lHntf9dYGUEKZSnfLlGld9+vuY/hBj7E9bu+C5U/Tv9HAZPetIiO/xkKkcZa36fLeRiy9xSkh846
G1tiLUy17rMwW4n8qWtX+pih4KsJr0bPGNbwFzyUJFJwj6P9rgMCZtz/6y5OsVKsqMmVbsi4aChJ
Io8MhQ910BuN90mEn/c86DniXrMJq0HR/kjm5aVUOiHfeT5UWIFVqgb5pP0JzShYbaXwKjlchpCA
Bq9LFofwRmA6CauPatPylX1Awz1dLCfVBXfqq0/1E2LJ4eRLS5Zip3KRDOgXDNf2+qQfxPtIHPNW
OyiULXb+GZb3gjz550u15tar1sI4EbEZQYledoo1g/WcmFumhG3HgNqg2wJKGHf14Xzy+g2xszWb
nWJijrVC2D7jgJOL/qNKGSl8wpKMIorIgaEmDNs8q1zWlByt2aRzmw3OuPnU/cIXibH4tfYi+a1X
7wB2iJIekw7RDM02JJ5PIHIiKB2OoUAidV8JiLqtoL3ZvwwQ4HXChA7SixMMVYecq71T4qsqMi+R
uBwE5GDpuGIUU3SerxmPRqXY2gP6gGdMvW95meSZ1rVfbs0f8AugrBgFnAjaBVOPhH/j6eOurCii
Z/T6mW9yDLmu9ZduxBVeBSke1lQ12z0wQ/z9xL5olSzzNHJTl1mL8LKGV3ldtIUj/SSmvGtWOKCZ
Hp9UtIhCqZmt+D72zizUvirLKEc36JsNr/0he65eZ/jsNPcvg2aXVXMM3xKR0AxNim50/Vmxg2cZ
flYDWTNae+kzCFKqy4NxOAlCcW+sxUoArccxoCRHMnHC3AH49KqOyZh9IyfPeyd/DVkor1tNAwfM
NZyqiUJpBDUkdGVERpbi2fVEKficEaBFQ31i7DVXanDWORnQDK6R1MC4zf6Km41TXL8ba3GDpXK/
VVup0bCqgtEEFjXRelxjP/a3FgY5WBCHWmf2hXc39X9j1j5bRNeHRBfPz+t3d+wascmRspsZPyAO
x7eMBRNWwZSr2j8rHk4MQplMjC4tFb0cogVn2RIpw1pDMh2jc7NvuYjiTIYEF/vpforFxxwZAQ48
+Xu8M5f/fYAaqz3j01jN6TldyfP5ns+IVk2L/XxpZ+BlFXopC89JluryfJXEd112La0RpaavdKns
NJ05IFghvmWrwbhCVasP/rHyOaQKmi48j4N7hiqNw+rkYhy2ejQQ9mYnMyAWpysTfpBx64GUtx/Y
etqV1TUl9IfA2unS+vfZanYlQ7sYaSA1nyBp+m5ENawgMDwWrrZQ+c7BglDDwKi0AbFpHBT9t7Kj
OSgwM+0puVwbx+RkPlwuKErW82/W+4+5WcEwk+vM803kp3ZwHm6CgEyi5fb64xzYHigSbXIVERbT
3FJSfn4GZv6eihZz5BF5Ayv3DIVRjTcQINp1kpDBR1hGfahHx0UkbGQxHjEqzHYqfB2ffzDmzQ9y
gkgXlejCPKnMuwLwaQqsu5tDrGFReXW1VO/zsRVXTLFlkgktsr6UTa3Vj4r6fKh2H2LkmemqCNWW
XsoH52q1mzZxn8XyFB8av3hupqJNbDLrDffCRLf2qsN2jjrpe9iy28IoBxMHkTx7gkIpQOrM/n1P
8775BQQdohJrjOEZdP4sviZWHPMRzAvdnP36U3KOTNY+jKbx571O+ZyYG3FuJkSnMZs45pBh2fgw
zlL1Ct1/IA++hsXlSnMRHDX07xVOR4bjbKdR2JO6rljvm6dDnKKtAS5OXbMHfNsBoVs00gwFMxXu
lSJuDe8nuUSl0PcwFo2ACd/4hIx/5ZXy3guwJHWJwko9C3Ie8Ot/skqPkwZwuc2fpCobfA/M/ToM
68KypOi68gaZ9dTqfjFpJwGhu3Xy4bjFHIx8xyVG3jDXiOTi4vELRLMuCekcSPq5WrCPpmdgVF8i
xogxDTrjZMV9w6UHCcp5BU31C8VX/6waja8mkmskcwonmc+aULR3FbsXkZR/JxbO7nsVP17FmyJj
m5STUQx6f/F+yr7caZyoOY9fu0uLvdGn2QWW1yeN4Iv3N16VHCW6DB5repDjca3maNdlEMghElVH
yQLYKrfnEWAfsm3sXOjs11FjL1YNSbuRCx+2AWUwDutGwJhz9N5zidWInH0l3FQpsHVl/ftYTKvP
lGYdN7VLl1W8fYI6pkwoMW39nmf0o8SmgvbnYCI64YOceveQMRKR8WgrZd3JjN4nFer5I+kWLG+c
59XENZhb9lWr7EDM980+hZ4XEwzgMNGBhJ2GXcpsfsQDT4+7/nqVu2jUNDNAe1AY/IBky8kNL83y
xuqmU7tTAN1eJxohtIJniKFxqUrdQZS3HxTtSk2hJUPThyWbQ3EF5t8F3bkLiw+cYRD1ZFyp3isF
zLquv/9cHYrtU9cIK0TOYilHFBQamWqfJgKWvF81WjkjqR9fUkrNZeD38vYsQrebIQtIAjgu1g4j
GfK6ltAu9QuL+yICJ59DvG0X5109v9B7iRe96hNln65a7HEzAdUCprAoA0nVByBNx7YQWuVfSw40
0X3paeDS7e1IlPdVEaDDGjURr9H6CxESqlkqYImiBD6v9tKQwNX/fRZf68YaoujrTuamwjBkru1K
aFfX7uhzCR3opPaTgl9z+iKZOqlQvy9hTlHVLUqgSeezWZhGA7PfKOOITzdSYqALItNowQ0i3qHR
8llwsX298uddVKMdaXf32PGs3oODYt2AtmOB8rwrS8SOYauHn6JiKHjGhPhc1y7y2UhMJajAy197
cUtrZTaAChiElztOn8Dh7+p4Zyl73IK2u2Rn2DmQf4N0fa4uDDpCPzQRkf0SgLS/MEjrLOBCr4no
WS6prq6tLW7O1NnBoAegJX0jm1mDgXDfyETQanNEgJTVAb4TWUEDscAI860AFJB3+S0bmGHh4TUt
PiWuXD+2jSU8VKO08q6AhoCZAx8Aqmxv89dx6/25jbDGgn37prZHOsSjV5NRvex2PNn1n7vNcvxV
bVi/OGp0f9q7ICoZH0ubwgTavoSz5fKfj5Qgz2GuLUzSqH1blcg01j85Z8uqJ+SlDQqlT7PvKmre
J9HC6jSONK57R2V+6RtnsuFID3YltVRKNRGCdYlZYcx1GEPJgI0sgCpDp5Ky8jjYMmpclKkfSRTf
W0wUPXhFZwP8Z1oTZ4Eydy33NyZNGNuw67PCmaGIFzknvIfxCj2n7++ih5rQtEV/550wxZjZqJ3g
1nR43b27nHfIB/SYzmhoB3ndS71IUFwiBCXW2bDmfoprVTpbOmE9G0DThuEUtfVuN2qu5m+35X0N
RbHSxNC/v30oE7fTsq1uZrMxRMyNysH/mk+K4FV3mtLrPGc4hs7vulmU69LdU2IlIHze6NYX5pJm
QOyUcgY6wLvlsVJhSw4lauhtxveHmdX70Oc7bjW/DkDRZs8nH6TDX86tffDjY+zpyguXCR0i4vD4
yLCCyhDNIQcBe2P26kBYY1OM2S62N6rJPDi9ONveILDDTOw5adHpFpVGs3WngrLXQQ2mfYi//1k1
7C0LGc5eNnfU/TRhaBIFTaQDK7kYAG6CoEQxUv4OmkLHTfuiXi8TaGs3q0ZM9e/kD9QP0rez+Ykv
a23MzKJiVXz2VOGs/uxYacvMhAotbJfPcR7I8VG01E/kOILT5FRp46Zd6IznkTePa0xtMmlX0sLL
PCYycw9qjzY2ow3XfeyZQNvvv+anTzRHvwhmgl27v8CVIdZ/J+293jahPpZAgfJlr3uVMCaLC6Yy
MbqteRl5GM80Vlwt5IFFazEoojZAYTZ0A3ccldjwZGlK17qlQZLcZScBAQbZflU+RqXsEZt+NoVP
XaXYBO7NV1ME7vGbjYQ5yY5Bvq9zb6d4GzdjN9NpQNgknBj5rbyP7rjG4dPOf654AJ7rEbne1lDX
e87+gUKn228lor4u/xsKp9sJfZMIazildEpca5d7+E87bZ2LmB5z3sDwDSPq+2hdvtxcvlfGp7LQ
9cwMxEjcJllHPijEOjUh4ueoyf9hfrLqWGYxISdfvYSdyy8JZQCH0JQoRofVTDm7S8yXNxuOyXi3
miPxOO3rRyG8AeWqlCQzx+UtqQ3ldRDxg41hWb0UzQWIpKKsSlp2cAGx10Dk3t2LOpIFddaiDOma
4jB+DuV1cqi7TetFScfMyMO/HMV7O/gN1DtO1m+1SmrVxRYtGZwM1YoZqigVTjhE0pF+Xyxs7TsM
vwgya6hrKm34EeYpwnAbB/pADfxtD+qzatRLWbHy9TSiVgzhO6A1YnrvgfcZewL4d/Jg+Aaiob2q
aL1SKw0NbIVpJUfc/zhHX6cRtW7TNxN7NlyFMrbTc4xQ4hm1VE9kMNFVq2meUUv/AOKYsoI6YOPK
H12hsHfx3r7cjbZUM3XpUPnac+2Ep9yHiF1SYaVaOSPh87ZHLReFtA/FCUc0WPHaDNmoHdN9DvBG
FaUjUNrFL21xU+ww4bfozDMwOJU1r7OdPQR+dSBvhHkbKUC56alatf28JCK+2OjDuyn20ck0zrqM
e2Y4Flzq/CMKMTsqmw8PC/MRt01qKPJ4fcNYMKj5pR8mMFAeZJ+vNrEdPc7pdMz3jJf2rR4pqKOy
Sh8s5E4fUCyAevV7npsvJpSys2DfwEivdLKnKoOFOziMgKjoIyvmuvwZFUl/QKtb/y8izYGY1dLf
8s0OJr+s4jtVvAkdywpTHOGepFpwW7wfgc1E3vhsqX+wN2sUoIQtOGeaWhT4dAtNu3G0VJHzWS/B
dnmQETfapq61AsXzPJQuQCBczmag2/DmHy5B+n8NlevVvGzplzzktfHcFhYp0J5V5DyjRMIlW3Qg
IpGT1pQ0a+ElduP+183h4oUaC+PvJgQ9MI0tRCA/5RD0jT2Tf/LX7/QsE/2UheZZQZqEmPl0rrjc
pMWdte8c/plj3+5Awv2xRfPajWOTKsv7oNj9FGU0nQV+1OyBmlhPLcqzouU43YpOcmXMzrRHaTJ6
QwRZjV6xFbZ0Pg1dMoO2eHIiipRrUCq468/na9ExqH/E6Zni+TDq2FmJpOlKrN0xEF9wvXOTAnBG
VgmWGY+Tip2XTX50nrCBbfQ49J2b+Yefff+0C5HlrUL65TVuqTdSyPdlQmXGXGE0ZV9SwOQKXkb0
s7jJIdFjjECIi6MyJ3s6EddVQ9i2mxac7xgMz9sZ+c5ZBRSgBO5i/eEFaGvBQAm2tZqrL/XdlvHi
TPKmSiSTlRlx064M8huZjhrakW8ogtnYx+XVzvQlnO4mhZbrLxYaoTPHee2/C1WI3NjeXM9cxe1U
jdpKxtKGss3KpuCp1HuVLYiHfjQfbe3LCGS8guDfJahD0R7eJJem2TtzYK5uPRosinzjxHYlVnUw
2g89JYpvXSzj09qwQEoMhuZ4bx72f3x2hHiBPvRBRQxNFzQIjoMpp7HVdjyHJ1tb2KzBthOoKZC1
ENlzZj/aZ/0R8+eP27bzdNCuMgzHz8C2d4V6cs/TDhvnDSPRM4PY6rBhyoo6rjoF92dwfjON0gPt
v4X9WDE+6dG6eFk4YAp5etFfHvOD9QaotuoLJvL0YJdRYmWVbDpNKD36xpZpeyNk5sj14ECz7FOz
yMBmQzEiwyxRYAj8PkakY1BaLWXuaCWf55nr7sHWPxDom8Ir+SSecPvyLJF7cn/g44tepSwcHqCU
JE5mDV0uOnSAd2rDPdAPZ+6iJIkM+Ni/h/A6cgmzF389QgxtFDO4PFv42jepDQmLs9Jj/YuC9Fi0
LjWtfcOFydSdjiBUQXPJu8ODifdoV0jHFd3Hec2oSVDHEyhgeRBmqflsJjoB+dD6Qti06jRRts+W
iWFvmC7mTDW2jnEp3sgmPGagysKVYW2mYV3nIK6kn5dlmKmFwV9aNidSMlM/p9b4L4W42Xbd5kiR
/2RSdrdCH1vaIWdf67fnvnuUSLYPZflwN+9yPvRK6OQBM1fpfjSXTXt0HgtD60eEBZAD0dgOh4UX
Z2hdN5HFKosjGFvWO0BQWZ5qaFFz/dZ9LtXrypxUoTTHDK83VrKM/YwqQtCL2ob1vJOfKwGcT7/F
eu1J0YyO/8/7quUNkX7ut1E/3VnYorljQ2fOk5mi9REgpKzotj6zkJWXzNMDTpLYSSukZrf7+63o
gaeVPLbhQ816EHobLFB4+3v3DUUhSNny3ALTuLpEDc8o4zSxzf9yb0dS9NVSpLF7ZMoBJKy87IhX
6GvvaTqHiZ914sxyJvPdMq2hBe62cMR1ApwyMVhlz6yBOVnZdH1eChJW51JL2uUU7fjgMhvN91Ua
tmcqXXZvv88JLSig2d5k0cLL2B8p3B7rMHUQJV1W5MbfKLtYZ0JNfHLbkoqkG+3PkHVhpg6vBKMQ
8J7Mdc8Me8NZNe3hYkJRLp0KiDiXjARMLMF/GVE/di1bym3isfvWGRWoJhvBjYepzfnqzdknlsyY
QzlkPqStxIi0P+6E5OfoA8AnUD2DO+nWdpaaypbB7ZplLJCOSRwVLD3O8nYIAq4TJfIIXUXln9p1
USp0paQzwXXO5YtXIuKKWxVRJyIsHPg7EpNEuxj+6eL8JzAoXLJCNVWKxbF+fCQfhq7UhsyGPkIo
b1v4XRItKrZ/49rTox1lC4HWtEJARnXyQhwpMNYC8r9OWRVJsPnwYUFrDSf4F6PH8ZzTNdzAuJPj
oZCUC5CEzkZ/RS8cwAi18UURtzZyPVWXnpjGmp1W1YSf7Nuy2teWBeKkS0VC9TNCVDCRMSgoE5f/
FCiytnOXLKT3pLt5BnxE2mEqHd4f/MnSQt9DihRhAsNGEBRBy5XjvLba17iyeEyTUBRU+MIa5d4F
zNkLhOIp6OLP86EAivHRbrTAY7/Nd3eiHfNxGOIKZPhGviviSDWRRYF8rzwtOHoiuF6vfpiaXR0h
OUi9qbmE2gfZ1DbAv/gO05RAtg3QOymqI9ow6A/xKwZa6RsRQn7wqD3yG55AvLBnIz6ybTVCz5Ea
nJUCdOfHSk+f7v+iznJmZbQGZzx/NwYhO6vfXvEYURDlzmWE/Q132nR1m76Mr2mJ1DBAvWW+so1r
n1ZhDz/CUbevkS+9MoEjhpVMBLafIg2Oe15+f+/p2/7PxKYQ5t44TSE6yAR8s/tJFNscbPQg0vLq
b6O+yuPhOFqOtKas6LTTFrXVn2cA+w3hbUilPmUN1fDPeW/A+K2SmmTkFXIQPw0e9YBgZPXnreO0
Mzh+3JIkoRpRKYDNTjZkvLthrEpf05b7hnu/jFl+8A0QAyysEeXyp6vMDXjZH2vsg2NZU/1IbPOl
i0pyOZn/nz4p3AWj4pXXJAbiJMfP9mJXfZnN9TBxto8M3LdmyaNVwCDJ7lauDX/IIQj112kyuKhq
YTiOtyCjxh0WN4w2fExj2TBREKltrr1iBK7s+itaQhtJjG5H3/53i4ofGx5UAXzUaimhCQGjC0IH
DOVBByWXqxl2QRpDufNNr585ixT3wl/3YeK+XeUGt3RhQEpJ2HSzWa0hmUCFc6oD85wAJ7ZJaJKD
0iiJQWE1b8JsTxfMA3tsuCoaqvkiZ8BNyM8C2Hr2xoCSk+q5W87n9gbHUplY3fWmMUSYz3cxLnun
Ec8zrfJNqMXlmjq5yrDEJe8UneuJF6oMpxpb8oq72ycfEPpZlHOrPbEbawJr5QpqMgwcVjnxo7cN
MTZzL74OCHyUoAgd1Ot/J5rpDc84VsJe8cFgThPYV8RsLTcnpm+i2PuHncHUPBPmSlxObKlhuYIk
FPy0+s5Fsq2irTMTaXZSCiuK89Ev37UzmEeBjRCT7tmbD/b1d/rCyCMtPhJYH6dbmZEWPl0hj0h3
xoFlLUYzP+qQE6acDjbCIB1neAkPH7QXQjc/XBE5L+jmNYZat77U23SDtMK5X8j27TFFWe1uECjp
XIO1S02H6yAhG/3rmHbecXJ4n9RChsF2YkvyhGkvs13bKdOJ/6+vzJ2wxbPLeyezWQF7uLsQJgOk
SC5KpetzZxDnsWoAgyt0YCiqU4yrAn4amGq7Rkc1h26nAIK8OOO9QtTkfYqqpE098Keugs+pXcRx
BeG5jDMMiDDCrsMX2yJYvaa6GmqMz87QZGMifKmmjrYskP0GcCRxI4rU0pfa9wzP0RnSnhhkwNFs
mfnfIYaC9lxpb2SdtxaSMoYH1wIFuqfJUkgrTuZlwsxIp06XVTY5ZeUjrnMvUTXYQCHoY2PGWrDA
N83p5ousIJaC7jozjZa0EH6LfXrT1oMc+S1uRrh8DPy9atuTh1mp8N5iCyHCaJXWouJwA/0Xx3Zl
qzQmvAVCaS6nVj1jD94M5aCGM6z6s1hC+rdzei5X/vBGKUrHLZa1x/ZY5NuHsP6idW/9Nb2a4LE0
MVRUSaMgrkJRQpkvUq0/3RqnSbmfyFbyJFmjK3CI3RYCXkyCPsS7RJmFUTxHx7gidOuHvpxRebck
HNvnNyz1/ReZTZmQm/qD69kA4b2+IgH7ikQ3HmzYVgjOEd66I41oHqPv0ldXZEgZRP98GAw9ldL7
xoqicU3cmC0Qnxz1rzYA4vlplJRsuCL9PBG6kxlCaonanuEfMvSFg8DF10Gay/TDYWoXmp/k5zFV
fB3ulR3eQ6YmIwDCptjBVI6cF2fd7zCYUWFAMgSW5akO8xPSnDqzJpjIjOsocNY/88HygRkOHpmJ
E4bLrFXHA4IuiTxQFZbMmEK4yidojl4psQyGHWtWzDxRtl6JQSvmrOsj5XG4amBBSUDvLE1yq2o0
o300baQrjNXjB+eTXk4a5nQskeG2kvTpf4JVaQFpsTD7ihTeuSNw1br4iFjBB5/Ph3fCDeOSwmGY
Shs44pYi+nIk1i3QH7h6B3uK1HCdCWso+7KdWbzQwFaKw/rNtu35QKjDVDqAZus7MhQHOUU61/DP
GYyFAu68kdmZgTtOIM/xJlzycf9aH6HPzrLClPKBmlzCiEwROCzO7GR86m53JNwipwkqkS6P0ygF
qNJZ51V1IRX+mY/9rnb3N+ZzcUQfw0AEBTZ/D8PDsXXkW43ESgjRqTO3GaMKTH54my5jYgGt6rcA
uggU+L0FifYR7zByQk1RMGtgbww5YFIwrzga83Sqo4cxutswXDMu8A0zQr3EC5rTt99dy27rpSrU
GJmK6bty37KSt/TsdDeHErs421ZOfxKfz40aj8XEzNZJ2BWv0ERWwTk2FG1jkTX7pYOU/XXsjkga
M8i+DFLDPfPieTLxMZrTQBQ11+vhOzf1XSopCwxE2EU7NZ2SRFZh17alcyjbAbnYcMgV/KsltOvd
Q1bob8mSo/0mtWFxZqG22kaRBVMoxapj/86fMp8LLt6IEt30EahIS5ToUuOBnZypGBYuGICM0KWN
sAUTusMxnYSYk+0e14KJDeRuEFagNNFi636Hk9O8PaQDHslQQs0Oyc1sLWzWhES1cjvVZvXaH13E
bCmIXoND7Pv7UKGAYoo49HfKA58mc3jDw72uvlh6i8968Y5UWap1af3+cnerE02+RMlxHWEmTX+W
9IihIOf28CrFYlb8Kg0se2JbpNDrtt5wzZGLT2titkuea/q2/H1pd2V+Eg26Ew7gh2hQxWkMTn4P
TL6vkXPRrp65OdXKuvf/e8jjAazcy6EYYcPNkfRYdo914fQaDqHPiHECYjbRpi4irxIxGHT0jYDg
5c6B2oCG0CUwPAOZqejOqw6hsA6U+pDhMmgmcVVh0/qwstUlqjs7siSzvNIbPN3n9JhKSuflEkGQ
F2szI0IkNjJTQ7qm0/ArDAocE1Rpb/DSBsUJVNb9mebutDA3WKeT/J6IR6qGQYjeUgiL1/t/KQ7e
/G+LKKfsehR+r0MFEr65Uk39U62guYglnVDciS9HuHMF81fTf7HL2onHbkJTXTiQigE46dEym14z
U2Y4MKxnknHG5yk0ciih8CAqPDgje5zyQ7P52E7+NVVIVat3qzHsJ6Bg4P+13jo6ja0wT/J2+ar5
FViZ3AFZbAZ0xgGv8L25NrC+8BgMD06Kc2pxZvPWrNvOi5fgToz1212L66acDHuR1oiu+q8LT1DD
croRE//PA4rNyyrMAiFoKo1brSIH/rT4KFBsHErsRMcv8pkgvap0WzaPWFK9cGBp95Xdb6kdpk1t
23kllUo1FCdxg7pvB2NdlcXzhIrdbRTFGyGeBWDA+VXQKX90b0pR2kuhUepyBKOMIl62Hbu8KVLk
d/jFIhY594Wx9dOPToNe+8NXoEc7CHg/0+onHQb/1LQFpLk6WcLVfVnf+1iWOPcwZX+vvPiVg0oN
7+iTr5KskNyfYGHxrhQVuoywB97i4ggoGLiR9kq8gI/z0MKP1vTXp5Ggxl1+tK68OO7ZyrwsKixY
tlE3bCQSt0vs1/E7avaWkTDYQk3u4H/vHaNerwwfpuwbyeVyx/X+5ImJoqvjwowCDUrvcydZJGNy
NhYfETdDibhFEitVcSMqxxKn+7oKBjK9EamkBQA9wYonR73+1xlzSZMP7/s0GzB5ZxxIeYGI+mxP
bcBcWvnJjx5JbhGMVkCKF6GQr9LzgTnBFfHMV5XHOCJiidloZCYj3kEC0s+xjkptivUPJnk5guAc
RDP82tMzvUzBdSlgO8rvNa4W0gHRYWWVnnWxfMtCHzcS4FHc98vV2mdJi4b+YpYOXEfLIqYFDIZr
4z7NXXNrQqZB4xrJYhXRXu8M5wfsQbM/nxphNWbqnd7ErK7rtc/eqG9E3rlaCjpOoQhf8Ab/7w1z
6/Laald4EQSXPgkKyzoN916UW9EzfOztV63bRG+kFYbpX93ZvJt/7LlxoIzkRmvWP2G/O94LeJ34
qBl1G91nh3YumATRZ5YTStOOIfubAN46CSek6Xjn1hrtgrHEQwS/e6RubD1PK5Mv/tdYrN2h2yme
xsZdHkV0iuZkTKWsJVtCM23WoZr2u/HV/puRMSKsh5TUkIEfGWYN9f20tcoS//vKqoPPeDyr/xFX
sZ8COq97eXO78ADYnB5m5kjsYgJUSwel5BdveYf760q3Sb4wudgTSDBtRkTBt/jLsiQiUwiJ3KrI
tZWksPWecPNDk+LlUaej6ZOVwRuZaLYc8eMyFOFuZ9+6hW+JbT9FvqsIHW8nONPw+nuSBlrBMZaa
Mx+CrR+apwJ7pSDiSRkBLc7HzYreHTEjrNTHC3La5H11OuOutRdJ26R0LxnsQ0N0+NqFhPuMx6pc
2IChGtNWsJFOrcOEdsagxJ0T/ZLKDC72fFy/JQVitt1gAmNCwiES/daHj73Ks5aUYj4ACdtUn8X8
IVNlWwh30omAd6XI381es81UDmticgf/ygPmPFw9KG4pBbu4tDP6Nffr4Fsf2hJX6/eKN5AsIjgJ
/41u8/qnAeoNAcV/Yhfh5zHYFIh7msuamJT9GsyzX6KWPQQpf5Oo+vb7MAjH7JpGSo62+vHEvqd4
wEo5Yrr1c2m+jPSyevtGW8hHUTNNCBSzNp0AiIN3h3LY6vTsoEE/IoEeGAc73GHnAhP/zuN7yNMk
vk2mSOqcSkxMglRZ7JqCioUcW1CFfK47XS2LOq5IEihgpkn6+tep5Bd0yB0PTqlz7zzIwAPuy8Rt
lxfXpkXBYlYFBkAxZ/rssDY2cllwo5xT7e59xy+R86McwF3eRX/p0HdOVGtL19pIY0KdLxhuVHYW
DeVnKMWm1z4qenAISvAImLyzRvUHq7+pqaU21XizIlZuL96o9qbRcEULNAbiacRj0BQTzngQgcbI
Y4epJI3nqKyeQygaZIMxbnjLlpjbk9O+3bEI3TeZm1eB5+c+mHjleiiaAia/2YZupvEUs7XYiXgt
lvfjn1TdjkF1EalnwYXtHslsBPOV8ad3MbKPNnd9G/IqhRLM6zcAZsEH69VMEKHpIm9mdNDkmmIH
fBJP1tSMJF2+/4eFBhFo2iZD7+PhDBP4fYTVbKq/QgsN50awfnbGn2HkSaq0P8zYTSsnElZKexjN
y0/XUDMj8ZOZgzLKEVsiG4zDaKbrYQTLIIqdQ55K+wNbwqhyzzc9xif/BirauswWaSWxgy3oPiE9
LjU+oUor1/gfj2e1ontGCpJPlByxuXhWyvlI0UFmUyWFEf9tRvtvzsrXVPouLyA2ORzpfG/AIJG+
V5WSxjoOnshCpnjDKiEwWxaUISHURKvE5JOM2ZZnadVd1X8HbekEcdH81VSMUHQPzwFu2i0cE8bf
VVwdLSrkaz2hbVkVOuHWqbC+txxt1LydJf/5+KFuHwVMPw5xjSAVPCQAfkTGkamozJJ+jEXVfixu
PsEpVU0A5RHYVT5U9thviqOReT8ZmvSzaC35EvXUxgE7uolax9MUZR7C+o8xYDO9NcPzQblZdXiK
7K8xkB02Xvg6ojKeOa2qvnixe+4BmBLcT7oH06oV9bMDGpA9on20LfdwHkUXvV6f5P1VqxAaovD/
AX2hHIYQritWFMxRLbAWxJ9cB1NkMcyNmG5VPTiu8sB1sSlosgBy7xq3VqUPwqtByqmVJR2Vv5r0
RBToOQ3CYn2QwYBz/QejbNrhyGTCw3uy0IHaZPC834C3tefG3Ozk+vTbkzrrGrsS6zoL8ystyEWh
3+qPH1AEc4+ymg1ZUSKwSt+wHHuu1mdlxCS/mwQ0tv+kjwN3RwwXYap/s7piVDPQItj7cXClHPkA
aQWRsNLhQfZVIj48SvMAJSFuktOClRcMDWgIL9TTtTgZG0rIt07yl7+MhgfayDK8BdFgbbwUO9Wo
82lUv1gzl845XeV4qTQrEUOmuLWvQsf7si+zM69fVQcqBC1p0heO3MN+q4GAH0rwvrc/yz7WWtWK
515j5GLe7rlV4fbZwUEt7jZE8BGgaTAhvjxXokYaZ04QBy2dR5ktrfsdOZOZYmjufbnYNUavs5s5
Z7tUQ05ANn7A7uZmy6q3rcdOwktkhjuuX3pl8lVU2vp14WjWDandSGvVWLD7f+nnDFCMHKZuPR58
CeXYtJs1/zh/z3kaJdn90usks/JNVjXc32fKH3l+T1yARSEcrXeNVuI1SVg4yCQ7Yb+5ZCwLug7M
xt1ahYh7pxHN2LYvLFOlwWMAspUxM0v33dS/b01lB8jKWdUlWQk99II2AZQQNQR14ater2cM0Rti
IO07uy513JDOqsZvs1gU++UKB/w8jeqLFBy6Ih2Q0xXX3fhi8X+zayaSfJ0bm/AszSpMm8q8sqbM
XAUnsfk4Zv3cL8a4+SBx0SThRhKyAUftYOcc8rITYT8vWLvXdq5itvuR9adSVP7kCZTrbRvg+y4T
eXV0KMNNIDJqikcK2DeegyJ/Vy2Hdp2cceGlCYAJd11vhzQQtTn+bHH/e0e1fAVIs7/UDDtsYFHL
ltX2jmkQGR+P3vabVyb+JdcGMI+uyuJsAx/ZjQuOjc6Dbn7ta/Biqil6i8mYdB3NA4tqRLAe/mJB
8upMH1hlRXfNPHh83ZByvQ+P9hGGiuUOgUJS5M39KXWOlLRmCJhEUwpClno9OrmqIgmUCcM5qyKh
jywqT77G6hrTvrKZkfj8l8+hSinanhv8ZS7mdU2FuQ6vNcd9c0jLfcY+AO5XxW9MGWC9IVGI2t6B
zkpukz2HfgavUZ4kOux1EFgrzLqAWsDpUurlkYn6cEBqUpyVM9v5uL5UGTmlIh/p4OkDOe45NQXI
3d/xBCMvXsM76pcUOvatZHzMV3O2OAtwm6UypzR+cR9b6lwfTuNJSVz0+dRCcfAcmNlCT532rik+
osl3QwHmd3J5WvfTBnt7jiGvv0Fgsyxnlgc3w+vJeU6DoHYFrUfybfQ637NbdOshVezgasS8aT0e
Yqe0G3k+dRg4TLiDg2Bk0FsmUdDjqSG4lVeJaA2Zf/HMCzS5PZTJInHIBbGmcllBo9afKvP13KlR
F/tNQkO6FA5/XhYsRECfbEPhVEVM/04kyr2kFQJj4S5LnSIcuSbH8NupE/qquHvxhQ6VajSUCcE5
THd76PP+Sl+c2BbY/DpZhniSUjRC2jdvxOcTcTAImufKyMB3Tyvnc4dXyqfSD+Fh1hKLJyh1Hy92
5d6vsj9SD9xzAc7wphlXNBveaV0qSey841OB6UjDuLGF/uC7/q8FzQrdAuY8309fF9q4Zw/FEpC7
BNSJ9IgYd/4dhSDXhZJyV3ASxwCWmefvKYiaXKC/rwMY+QCcxT7QFd1ISZQsiGJX2eE6yhTfB8wt
ZNhqAqawCSdFDc/xtrdDuwMALCh6m9CD9wluUxmW1lyYrYfZ2z5/FBn+ani8x0x+csBeOuz1cx5I
DTVxI8F86+6U7ugKqEyFj4RE4QQO6gDj8lNIV7HTvZmOiu4S0WmUdlz/hILJ0sqvCEX2yqwMJwAY
2SVfTwEDzuo00GqHrUaREmMdVQcRqKblBWlAowkzk9SwbYoVKoFy65Jj+Mgwaaj2VKWD2hlzMH4O
DnZTTlFDaGqzOCVzFQzyuyS0+KbIYPRqzkRPDn82fa2NHWihQ89xypmc8tgcVO2TBH9/sgH3hBHD
1GywWFu7YGWldyJwiK2NdJyiwyxGpiQlZ6axjoIQqQisPxmcPc7nCs+ESkRrnYy6jyhBAO5Po0YF
FqstBelZiw2U4EA7CDmXiJHl0LgeV2EJZXEXuo3ZJuxbETwt/okI5DOPtyaZi8dA3ZOwQHbsUBET
Ct86JmS1k9bfIY5qrrZBxHxj6YeZK1gSvCJ12vwrrVJVe/8cM0lgTV6ruNY29EEoQhh0aUA//9kF
MjVnshhmML4J3dkdMIkQfFAErPebPLyCJThqYDIulH3K0Sd4tDRtsaCGrlZV6s6z/2HIm5MLHd93
fhH7XRpLrsCkfJxrBnytG5Sc8NyMCreeNoEx9j9ZojMj4HNJq2IDByifVquIqhXf5FJnmzVMjgKC
ROgmrC6mWOpuKOVn7uX1pXnJLKCZ58nJr0SD2UNDPsT1MRdb4Aw/AHeZFDZIGuA0804hmtyL+td0
wwoALnhB1SKMEABB4XQAwf200Lkg+jI9PXKLjgToXNBjTtXrAYeJ69ra3/a8/1SbL6ydMSrkxy0C
iFcuK8VEzE4ilMQ/NK6QIFQV+yYVRWnUL9Y6BwsYMkmINYcWgjHFhn4LikdamWp5pi4JccMOQVt7
2IdRZYRZtrQv46CC8eJVkIZ2P4eD6FS/KpbsAJRGz9aOJHXpVsjBbFI+EHAscuVv0A3xt5QRQgjF
XBTGO98B27RzeSAECQo19TEoj/1282TysiCNjnt/ccJ20rdCC3c3kA+z6UTsjHb4JiWIdR1PnaW5
4DcXjNiXXm5l32Sa70/KxLu/gNr9TjTzP1a6PEh9eKEM7+4P4oJn2SZEmZjBseFdUWbKvolpD89x
cw9CWXe7YOikP8OUUAybVMD7G2KNnQvTMdM19Y+KHpNpCIvP6lmBNCX0YodsbTGT7fP+ULMeYJdV
B+WEHyczlmL2iV6EirS5W2tnoq5MUWpIl3szObkXA0xuTS1V6VFACfVao2Uil4Ek8h5b2GKvhGEC
WtCDqJpmj01ZbJyDjZ/VQgvmMSbADZLzCuyaH7XiK9b3Be8zKh6Om8J5U+YAtAH5YUeHstKdSSBM
f7/6JOen78rsjBxTD3HqZzRlY9bjEZXSZuryBdNuCqzWNtSVXNlix1coIP8yMLzxNFPk2lVTyuGv
F3E8AgYdW4MmNgvgbX2lPIWlIo+wi6npDXHphkUX7WnsplOeVZ/AFpLOeQBWw02vUnCTX+ZRGA3y
8wVtNumV6F45kGzTkmSd/vcVmBY87ONARRn4pDiHlPN/7OvNCvh1z0ww4S0QgnWCpfNIogCfEM1o
r7FCcpO68QqMVAUS17HRv6oKiJzIcLvmIuzkMi49CFgpalb8c7nzht7TmGbGtnSc1WQAGZN1yqEx
+In48v7h3DBakpMo7SgdydS+B1JnQmTjFXvMa9WRhG4N1TQaFb8MfCB36BfesECUmA59hHDqguCN
U9PSriTnJiw7wWlH3nj3EeAzLBHPN2x8OsL4i75xsDlti3GWxhnwBUuh16KylmwnJ/925Wpg0jLV
4zVv3r/wIfKAUL74nn2VjuwBNvRIiZXl3IXd/YNwik3Q6DR6/EJJf1n2AEpcgF4raU+2r7qTEqsI
x0x+doKccxtMyEErkhncrm/E1bpoWkBaPnK5HZtQtzUSuWhQ/6tXbIRgBw/KYXb2KKXnGKZV8eoH
1D9wRZsipiq6nT6+dxjsxi4RciDQ6di7vrCO0yFmKnziI9aOspH5sOOFtVgxzBUvQ01y6EbFO1v1
YtIH45T5zgvieY1E7oCvA/XTOJQss29TC2v4YR0Nzgqubk8r6WdcH1kU6eKRdItfbxPHockD4ANj
sE0PG/uFZF+CbODeRJ3uCgHlh2Ku0OWkS0xhxNh8ricfusSi6hsLUchs+knM4MKW6UA1YxylTvgd
zwm7CRw95plHdV5NsTbblY3Rdl77kpGWJqmkJLguTjtzJMLYwx3HnfnlZO0hHL3jql3bzm6CN7Qj
gTNgX1refEyksQojCsT6/aDX/7ioR3GjbLzFwZSZaVEDsey89rNV8aAr2oLok82kgOzTTn25PtDd
bvagpB0hR8F3OiSILBX7IybSMEjPkbxdfDSsoTDYWCtbH6pAmnYFW9N04jtqrmk5p25Mb8Cc3rk0
Cy1l8oDIFQKV50uPGig1qdM5/EA2CO4wIA5nNTPxJ37x3SlxC302dL5a7dXBLJLYUi3KAzYIrUQm
Pun6ogqz1Kbow3tgGaAykD25DVGIyxEcZgzr4dNRQTFafE1M5R47il9e6Z92hunAOWP1/RwwXMxB
7wMQVYHpkorpT/Ceq+nk+5Nq1GEcybSq+xcCXmqoutGfdoecNeJcTvtlvLbvOyA+aiIQZdjyN1jr
SluFFPulbiE6tVIv8MdeqaE370OQ0BKqENpc4QnktnCk6ZY4rWGbcTuGHV09WaWGzhw9Xd14ljg3
O+GaEpOWmnonLLNvkl/wLMR9DEMjpcMQcZhda3m0bqa0MaVwfLOe/GBsom+mSpaeOR05ib0HlgHo
cGu2JorRMpHhsfLFcsQggui8g22MYnWFq+LllzRaCjsHql+unCLiS3s8MHPlBMrZzbLjeM2wjbTi
bGnmzIDLz9+c8t83C1lqcITHuneqWy9S+H1vqJHN3hB2zCs1JuiVSZlzf7U3cjBBSGfbR+PtMtAZ
T4SSREx2o112estkDoVbpxOI+SlUueqFzeBPAAGMG3Ag/StqzFVpPPhpXpw8fNUWQuMhDovXLu4h
8pvHVgVB/lWPXxbkB1u8Fiqt3ymhWCJm8ASLGlFW6mR9HHTJl3bMENi3c7ZDCZ58xM4ec/egOML/
7Wh3HafkP80jA2Icr2qtGBoJaINTCmHvqhP4MWS/ryK5un5FNF1gmWcyGdH6/wbR1oO2Wjp54+LG
d5CnkBEe84+q0rXvRuPfo8VFqH5v/iDMpPEa6zSc8UMHuJpBSy4bXcaT0PC74cBYB8CCHcKNswL2
DKBieD7Zp6yPVixzYh+Wuu9D7e8QYf7THLNpvqVJS+eJ9mQh1u0iykuMBcwoP13t0JTVwSt0UEUK
VAsPzd+MTJVHTZO5YxviLaxfyxhuPisrMBt8iBP0ZN54VfOiQ4qVaOMb83SuOTRmEnsXyQOo9uoW
nuVSZ63BKTXAramLTUH3PlFacDi0wnz5N6CZM3Yxl4bPVyGD/PpzK/qNIxbAJLDFyNYUOU8hc+Hf
ALSyC4c+J6OI5Jmy6QxJbDt4YsIla6x5x4MZx7zeoNRGzDNBCspRODABWH39LF6iWcw6X36xnrGu
6rKmqcbrMirFLMHp8kaDpLvkVNu/7Gvn6a2GtoklIhdIdnSwRnNzdnZI92EszgF55ZQq7k7pdZ+b
caKmRcOSh9ax6cxmX3qolSJ/NCM3HoFb6py79IXvpXYk19azroTUSIiaFHHKNZGDwjBB7liIMhF7
3tb3SF5g3S45kYegB5CVOw1vRDj+qr8QvFyF6Dhh4UAh8P4ba/6vWuN3xPihK9tYLKRvWxdXPJs/
l7GG5FQJXOkveytur0LqtsQB3xHksMPJus4C+1HMjt064CPTAxCG6Y1ZI4heFz6Qhs0GwMwlWwaM
0Q/UZg2ZLNtj+RsJiXG3jEVShAR/iMEUMrqBvNGovH9Okq0gjLQiPa4bEA6opp4p5Ht+SnVtHB8H
+vSF0ada8PIuK8zLNVZzxa7rfP+UmnWH/znh50i0aHJULcgofNyLhPthUGAmL3NKeyNWElcUb6n1
zKJvK8uTpPaPwrzSUAslfASFUQ56uLwwsHpBAlRDFOVWoK8ApuQDcVMBw4xCYLWeoqzjI/sD+5dQ
9RU38KrW7Vjw/kWuVpzYFrMs0hbsSGLs0aNSFscjRFafq+H3lYNCMgdPq76wtaCTrM/sheYwuWNU
hO/xVg+95ewLBivXx6gzTojDbonewgkGMZTRuoqbl2v6BLxu0l0h20yuS/fPlRGmdBHw9vlYSflg
ArGKVV384BMyT3uCMHBLCqvpHQd3LPUzTXRqJUNpKsthO+VHgLX8/EpG3kquS0ujD+g6PW0Snt3k
bgwo7xgzOszp59B/j+lxENlQ0QuHee8vkvvs+Nk3NllQJrFEq0S+SxKQjUn/SZ5v59dEis2O9k6/
fzRVavF0mH3fQ3+8o/9DlRsjHy8p9GK8hfXcoyL2uvyFM853wbVBsfWyKbJk4QYO6hghcZs5Zprq
+3mPbDeImz/QQLye5pPlwWbR+KMJ8SQxg/WBYALQfSb93mn+UnhvsU5ndy1Rf0kZa+58Lk2bGfvJ
BPCDKDJJjp7XM6zto77qfHso5H5BpPT0CXCA1tAFvhm5/k2w4FEFsCInBcu/uxXz3E7ovzXmmb9w
P/Z/4le/q3XEeOs8HtRbfigVpLGnuiQFznocgbKiSknx7RGsqGpGRL29SjmZ/TuRAz/cATMlmUCx
rcz2qOwVcb4y0KEHtL8xgaRZ5LdZdKx9bnjXtJLf4U0GZjbBJYrFi30fqrMrOk9vfydfare+BepZ
VvYT58k/qdeKAAIMsMbOy6JJtB6/v+JTSrdRKR82taPqr1DrUukMnE+9rcaME8IS0DyJ/RBoi/XO
MGmF4/wW5l5Y0H3zVXWOZw+S9gwZQXmoGZJiEvy9I1Tpl3UlMQ59LluLk+L0MsWWrenZANiMV6GZ
S+GkiFVsir7aa+wfHTX3SvHj3FrvR1Rhemf/u8uU11BLYUrD9VUxPjbFOkiIeu2UVVJW8q7yTlxy
yVfI6eq8f9Aao3il9sFpDnYKBSfUcSG7K6OliJKVWOrhKvvLz33D/2zKEFYvhzjo10VBYEi1xw9t
WCy/H/pmQcm4jok+yUaDe93xr2yiMzHbEmGCf0mjrc2XDzT0NgQ+b/eR+b0mtjHUV7PCbjetQ2Gg
v71N7XlR10U4Azk6WSgluSQD8GtIoUuLG/5Mk7CLaEJNR59NuDClM2HoS/3YAXOo/uu6kL1GBuYj
e8cgBq0P33NyxYymL6AgszNklKhzhLec3tLNq3EuaFU19qb/uVQXka1VNZvnz9mLZDTIKxTliobS
NKz2nlsGFSVZ474PvrB4JCsscAtzoiszWpX70Xb64Fi/2R/IKMiNxLnuahzZXcVohjE0OxZoaYAN
pljZZBUvH/gwW+w93hZD8QYuF7iHjhuXPQ+7rPethvjVAYQnSrp56m6nksXGs22l93TmBT38mgTU
SJYMlWAdSIdL4ZW+NBq1OWtzOtEFS2haJLhgVo/80UlliG0EyONy0WN6u8jmnTQQ1QmxFAcY4vgn
ACcUs9dDBqsdEqAindW3Tnn6z2nmUZzOyaQesIeH4Qz7ctyW5K9TTTqhK7NeB89ohFCwfFBBpM02
fesRx7f9r2qpfkVuc8gp2ULu6yAi2Z3J22LQS/J6En2YJ1kmLnbv+s5ay+DT0qTggElMhZqpCeZK
mMdDCUex++khTlcK1Yg0ZQUBq6lIPcxe6KHhPXj7qCtbhMWVmcPb8v3u8yVGgGYtawMxraRlOjLF
MkV6lJ0aanjnZBBZgp3yiyXzG0ugDlTUk0ACR6X+SZbm7klgVNjY30DpfPbKLxDrWeeIMoeJrNvz
9bS887uvz11PlGpffR0+CqHE1QI55urskWs/7Ro0XKsRlwOco95PNGbmoFY9VqE1vQXQQLBarSnw
DhUXx6HvqaMZg3UML3uW+rRO/YcvVCdNrQcY1Ius8eWcgJICwcuD48hDwNHkiYXGxDTtZsJquUba
ZEyxOxXgDvZqnAUAY5vW8FuLHqdXEvgdE6iRlnYqJzPdF0K6/YpXybfWJ+VApAx9X6BSHuIbfyjF
xeRLB9FzUlrv1zaLN1ohposeGMrwPGnqqcMRaU79t7kOuV9yvY8IgP381WpdItTxHf8+Kpa+DBKk
I06cxv/b2qKHL7qoH2lS7U7mmgM62NEfNbV4m1iJBs19TaNsBj9vVhVpb1vEyjnxsIpDURwnU4eA
u7VtnYOuQDobXYp7tj/IQMRtt1frszCYc5KH+5ZKam8nA03DPXX9cy+5cGSQir4kbI+iaqVX91q0
APrmNrHKFga3Pi3hdNWfBxY7UwR27sddlK37GIEjrueTZAY4GPvx7LhE2teLff5a5gJSkh+XcRgp
/hJhT4NGxdPL4uHshxINJsVWjto5WM0W9Ky9xpxvA/6ybD0WXspvedrRJhiL4Md7RV8gim8b12UB
7b7LNdq4Zkk6fGkou0YPmqCuEvJMIGf6JAmAqv58t87tuiosUWvP14DgcdQZzDZmNaujL/Qr38jl
qEUNp1MDCta6svJVAsEUvYNbs/Bprd5UXRxmXpi8HPCEBcKefC5+f8E5y92fe10ZYe5P8zEXfwXI
uYbTMGjGg2NCpiVR+myyDYbBiurvesJIuM5sOKSeRPTU2jbYKxQ5JXWn7UsZH0R7eSPuZH5ossC7
BmG0HAN89UskoZZSAZr61wApynL3DbjtxcyJH56vS4Ovw9VcaD2okZkkZAeKXd6iPaQjpPsBhAVV
69b8CCFUQOK8ifAu4ap/Gql04vE5T9K/BESeXadN//VlsHsZ5yMCU7UCtQoASXZKaDpRkO0sVKaD
gB7x5KF5ZAft3Sfn/SNvPE0mo12Jl/u/naOZQ+f8ne3a7yEkWdHpO2utJyL10e6yXbQGLjtNrRtL
V0ldslrn32HHGocEmC6F+Y0RFsRYt/qb9tw0EFroIZoJULPTs3FlCC/spEGCvUBAD6bGJbewvOZB
Et9JY4gcNWo6n5UQPfZ23iGklSd+kcjnagtYOu0nUkHRRJJikdcCHqzuU+4geBcc4fW8H2hogUo7
sBpFe9V3+h9soosK97hn3sCscekZag/NWhNH6Fhzon3bHc+lhIhGtukxk7eEFFwURc5fzRr9VPXI
J4Jj/SzyUF1llop0i4j0O8bjZrk7CDespw4703JbaA0/Dd1X0CZz5/QartFce+8Bmjd8nz8hU2l5
M60Hi1VybKwLkC1pEmVBoSO5fHU3uGbnvLHtN+BexnCqkxvME0wPRbKgCOPPdnkuqK6xjJynJOVO
dhFrZVPxy/7dVr7JEwJIz0IAYVu6fiDP7He3ngP+LiPG4rhIO40GDSasssNrfMWF1g1ttqI7dK3k
7mnWWeUJVeM/jotGts5+smOx6gUdjTXzIep5pZ0RhkQxJSAWSPD2eXM0H3un/tysMi2W54qwMWlE
GH12uEPrVgDAAcCv3rnnG1mpt3yknRS5h8ktP63hotIVMThkUZYaGkg5tDA94mi0R0KXpRWeruDw
Xeb3hb4hpdPLlHZ5iivwt8itQfqy6hjCLc1iArNU5Y3e631s1OBik4CdA31qPrKAdDPQNgTAFvK9
wJMVBVev0zY32Jy8tmMLWHNJG/MaxEuurl3PJaNsA3YSktz+pCjIdGsbUeKA7JG9hsABnNEinNqr
7+LWMT65YMQKL6+ug4XG+rerQ+dQ7MLisNNqSmHmHGJiVkweuqD8bzZGkCbhGwBeyXuIS2rJmV0p
m8hXB2uNs1AMe71SMeN/agUXR+DY2EpVjfkmjQLNKM8dRXpAFCV63qPCDa3o/QItcxd4OnVC79+r
s+P0GiIKjnOu8GQIG8hMhQjyYZphh8Y7LMrkvQ9yDkjICXwN6fdMlI0XVehMPTitfFTt7T5jFBKL
nDWtEoM2suF2JcxYEaPlsWwa02LLF8/NfF7U0JYIKW9bysBa5uNYwnahg/TFYq133HmcY93ujCIH
6apcfXdWb4TeUBuNxCiPZsnZ53EuuG7kUhNvVcpCIh4Do3wNmVmEFObIUyEgY/SwXnMgHaZze/c8
aJj+YyuHo2YrPNy5Lapl6ic9ywpW6dba0ziKZDLcZI0X+WmUkBWG9n4fouIPJPwDwFTNSq9B11hD
jW1IGBvAGS4Xroc5aXED3j0QR1ufWIWqioFVujokU815iABVKpHheQeG6akpVVCOD7t49W+V5VJt
0FtzjJFscB5av/5+UeIdMHOzRR5xmfgYll8ENB6+LeA6BGmxes6/0uWutnBALwHbE4O3ThTSngVB
qJFeM3gjbB1mH7EQXKMiuSHWKHcP6aSHSFFL37D4uA3vNDY/0jF0KOayTcrUhtNCWe/zEXQLJvHX
39EQrMKyTUq8o6p90+N62z7EBT9Y1FoH+JsD65IvcWtuO5Gdy+FU++O7opzeOnUB2LQtx6u3kx25
gFPaA/Liok5gqv67i2y9cyMV508mxF5FiJZ0ZgsF/r8fExI/4eC5w2tSd31RVi7CwJVK5Rl1BKdC
3gC8ECRsyPUKKoFDzrq+xWKeeflzm4QnwK1lxTPd8Hn7TP8EV8viHNLOa4uNBDk/An64o0DnujyX
sajYliYd2ge/C17GdHAlduMGFmKukwbESmzgILBDMuaiGA8uwAVViCFQ9Mbb9DCAFfCbNDGdwAXw
4DNS+fSWU23gnpdgwIDRgAAUUx7YDf24dysiahrIRRQjntvbp3BUq2w2T1VTYchUcFELx/f3EHUn
9YoqZaTIQMlsFAzqoj1JuSNzI9v+fSN2vrtEjb89vjMvPnVHDn8BkoLuquW6jaM4S4Cnvx91pP4I
VEOCCDhCYuF7tftKma0q6f4tR0NR/SrORwIZP0tg9w1BKebSX3zsoONsMvf01V6pfMaxU0i8eFeH
dylkgvnt5OLlyH469fhd1w/SZNHBuFbq5wYKJIygmFzKCEY3bxpKlt5XtEz2K/aCb/hpFjlsuUXj
CGCPiGDPnnM9f+XtwQtozrR414lQAMiWFRcF9k5+4pG4n53Apq9U4wLZ1jezhzXsEr9NgaNS5o1z
fH4GZYnQn7QJAaANFJKWezO2+misbG+ia6fyhUfSvp5wsSelRKxoDzv2YAcxpbezhsssXl3FlhQP
180tR4l9IQC1ytPyNsvnvydLcs24xln6Oz+Tx1rutjEvfw+aR9vZY9lhjHGSISOLQJXuurG8mZj9
3EGs81nnv5J5uZHbfUwOMNiiSjlxrZOtbPwoKt7hx5keEVTUbET3ar9qJkJLbX8QlLWPasYowWns
WoeLpubEZJovSft16f8ls9OyTduiQP/6jQCgpO4bzCSVhXyfL4guER8xW1/S3hxWe/QJE84z+nPm
911hi74Gvsrvi5dXdQg0GxNYx6qkENGRZjSeqB6QTuotRDGp6DxViB7aUqYX8ERmk3oqcvexVTn4
f+n74Fw8qqnH1X/BGTn2mvZIWCyOaFLhouGLWR6qqOMuAiini9gDyiuKC6MxjrJLDKnl1Owb8bl+
kn4XiYqXkQxAFrXPn9xM/RXlnMg5htQC7aHhg3xEfYTKZd3aXeppA+x74TsOebitpkdqtdldLTTA
eaqXEO0Do8uwIk1V4QDXNpk2hc9x7/B8wodRHMnJtVlYY/G22DE6D4nZvDI/VxqBER2WqbShyrZ3
7oEgh/CYmrpsOGlZn3R8brgH82DljU0oSvy+0f2AeDClbn/FLnxRjCjG6BBtQuAVXqw6VTAPuQv+
8JpyQkaw4z1vsAc2Eycn4ql8DPvxxxf4hZV7ja3TI5axOQ+5ljssNBo7YwWgEEG5EopZ4hvQrNJY
twS65BU3Q/b1h1dwE9Ap6Lydy4ZmMtaZaOxaeyjjXlGy0zKr0mo+UBgcOQ3UBfTofwa9ruWLkllP
RcAySlWnpqgsPjpIuV0pzVE0KzRdbH2rN76MDnB6/56Mb4XRKWaE0Kr4Ez8bpDHXRcI4/UnC9r3b
fWGsNSn0KP9iYLWNZ8JRuoyrkS9PseRCrGS5bSjJ1kSE/zmLVZkopOI7Z6NFaejs8LbY8WZMw0WJ
bfquFlo51dnHBO5+8NVAZtenDOtlDiDvYzqIBqBHLY9JbTHA1zRw/LZulWl97Eqzv1bxvCCtpyjZ
vz52C79agXV3H51KFGeEJyNH3CsBgP6O+wBsCn77BOgmENP8+wjA0pGp/MVsUYI0nsD9hJsu2KNG
9aj9z9ejJxbbbv/rnUMlta3os+ZgAvoWsWl1AWCx9o+RoW0fZCYhvJX/LvIlgg7QPE97ZG3Af1Gw
6iPn2YxPPGoAVl1MS5psXXYYFEf8eq1EYDAgik9S0QRq1E3nR6Jg8VaKfhK+jfRDvqFWBmEptOY+
YpNE9Gvj89PIdw9q2YAPkREc5CSH0Een7XRkF9gYvQNxHqidglF1DwUrtEPFOdazcGl0rItZfeE5
tEf89yfboovB++OnRqNu2DWeWMDeeoaTAhVR55nqeq/v0xf2MP5ESbbgadiyRKFI3u/tqHU8583d
Y1vtjzIRRuXo0jWuvM+9CLoxwBZtI6JKG3+AgWit4kszfK4X82HNrbum9RnUZUMh+U3WjLb1nzZe
FWwnZhIgppdgMx6j+/UAW+8Galbh5HcWbD6EMyyCf1Oiz4rh0kJU/v/L8SX0YAIMqqLuE8sSlCo0
za37itAl75utkwmyes2HQoQj5FvpvWbQS17WxnRM/6Zp+hahYlxG/pkZtVZyPEy9lUNu0pZKQ9PX
UKurAmTvt4wj2ims4BXQIumPeWsqRxSZKIVQAIvxNXyUQnM/AYFt4Qrvm96Rv4eS67UQhWDmjpfM
RXNHUAn0rgCGqIZllcr+egCsPnyktb2fvNT4IM/KnP+VSc1T2IoR7azRPTVdhdT84w04abPPWp0R
2fW6Aj06Pkd+GglYEhRajglTL9hnWtTyPUbc+TNFTtFM+JQ37QXYjOxNKHcP/dB0sLgFoIdR7yWK
Ggw97dLtjbqBZ8AFl3O+LkxnpKNtXukxDP1jE47FQLxlJXUOX4gI8o635iLOo6euRb+Nmax3lQy/
2WHvcaqxQSrSPof+0qyTc/U9/dK3aCN8QFKJsFm7q+fv69MV724oqNpC9xJEPOwpBJv+sW9m8kFh
dYZe3bFGQQ7aYIj3Rtrg8iddRDQcAIT9bucH/mtArUN5GqHbASq15GE0k42VIniHyKtA5j6vHPyx
Zf4kcIHLyYtuxUKkUuS12IiasylSqThL3W6cpFOd0hbuEuhEEBk0P4ypNvc7PeOtVbjWU99xEHQT
8DMmOF4mfMklyhqhgWvxuRv7JTZ/bc1sS9vGgtrFtNC0XiIRdsDqis13owNYA8hegQy4urDbwI2S
dubdfVae2e3tS3tqIrUJnKcFXSVzohU3ttGlPTwJ8rWwfdqEEZnB3jshn8X00dyozM1RkhtjrMIx
xHqGMaJLzMky5GQOX7acO/H54gxvz5rDql8i+FDiRGQxVWSqzmkoOtm1Oqmx5Du1tC2ugIBHrsYP
fFy0VySUDcNOgzZJ5i4yIC4TDNSRay+qFaNuxXMN6xIIp+APef1+gkwg4xlVFgT6vi39lIR8QKIp
77UxjIOWa4tdixnFZwKuxd+jk2ysI5970gl9VsTKFCOsbwTNQ4Sh6e65TBbPy/CQPWGzR+c1xn1I
eWQXwQYAGrygpMUZgvBVH4NS94yDh1wHzEioMJaWFGPZ/Dt+Jj4LUeVVnNCNlglyqpE0HD2tHnK1
B0xkvbM85A9bgKRfCqs38sXri2FBmsGvssochj/rkdbrsyN+Ar0fpPeQXhjAWq3NUn2bdXaLP6S4
WApPWRz9+7YLVwFdQvCCATQQNgltmpLhF+0XqnqZ5WRsUTZNhlKXqMYJ17GVQNZlmPo1WIiS9mWs
PTin9wFS5E31o8aJovEAOpO4TnlnXflZkmzHmhOYukQbiOj959J7+1qAc+o4OzNYENiwTYdqHWOA
V4j1uf7MvkJB0yo87TLXsBVBofeoReJvQScXJM3HvkRjytBGB5dbB+gwpoV5odKsVXR8r8tW+8oi
xrXoiA+zBQwOwciGWq7GqlNetF9nRV81xoOz96qNWhToUNyZO1sLLn6tqsvEYI+ZYj8NMfRcfgv1
hrjqUePKflOBCzJ9hPtX/bYLRgaVw+6cGcD+7uBQWmLJbSTmpf6ad/pIaZW9YI4Db0XCneyeGmx6
hZ/8SO7WwbApWISc0z7yi0c5I27hzQSXIflWHVwjAmSDJ7+YXkY/GXSJd3J3npk6F/a66lXYeOHj
n2t/claEMI0PNFroWgkoCGcNaGvZ+wCMq+ZdT9IB0gWcPEe7BxOFm0XtftsH+9gsEr0GJdDOkk0w
W01j05jGkPtFs42y0H5xKhJNuEjM5ImdUN80TX7Olehj74V8LR281tddbhMYiPe4tA58ZxYQ4Ee4
qIuZnT7S8RA4I592z7G2tcDAlZ/SgQD54ZLqRbPQkZTK5ZbIbuXTVQUJ6NipUDciT8NOEjD8IqnG
VcLzowrdTjKNI0jLkqqyGMIb4C2VaNpC9Z2FgVEjpJpCjqy6IKM4MfHTYPhdpDLwAxr49XC8Kgyd
lVH9N6kSUmcY7h8kFHp16CjNnUYLriz2cuTDSmUJVhwV41Q4AziZ+qU+ONZYRm8tLLQo1RIagY0h
fbGjn3+2A7Lhi6e0iLJt+rAivLrTdofUe69Sar6QxkwgCprd825OljEgnkkQT72nfHB/rGty7NIT
ws07fiYD1qngAHvObpP9doEpAQy6U+vFi6oUxWXV5ZaMsO39fAbWbFxTYWoINUuUHY2WmM6lIWIh
QbdW7NVw2vEk62Ezzimtro+1oI/ip+m4y/UC/FLNVwfxgYjjzR3+kOJV3xZ9TqvycwxEJd7mTvSh
vfUcyDFwNEd6J1+Go7lZII8ZFgHG8lRD9fL0hacy6n2blA6mrozhzg8c0yBvZXwOOXAr2HKuXdeV
0Yn1bJHjxGFdQZHTXSKSz1pBFf5Y4SzoKdxZ/BzsKsjHYS5Du7dWVYlibOvrlBKlyuMDExiKfurc
lq3z0h+GZnhfGayyWD9hSffr/mh+a+7KicOUf06QWnTybj42IAYfwYjAH7rTyZfLflzBDGhG0UAy
jsO1l0o3Z97ZHN7oN7aldV/qghUxVlsc9vM3s9AMS00AxOxj6ew4ndgRpUTTLCoF2o3z81nghVR6
qB2ufRx5ugPCGBgTRKfLQ6NheUxsNXRSVSW1A37v+yGinuCus32ovVpL8vQl1Gy/IeVeBYmLAAn7
cX6pDs/ecc87BMREAczpTirC1JZDc4gu8OyGXUDczUkkunY1zrGuvuQdWF9fp2nBHNU0xIl9d77L
sUaxuYDbLKOPUjkBHmTkt7Seh72DaQoVaYhJagH3dj9MhX1vXuvspxEHNIGX1TsF0B4RXevvc8Dy
guRJCm/N1yvzSK0yTjPoNQbGNw9pwh32cVqc423emLS2b5RkkF+X1of5aBkZznxJI+c2vOpAaPhb
ESXFgxAgVQ6P6P5NgHvRBkxDz7FVQlZqQ2bWmzK/5gXJeqE43fxlS4mv4P1wgkiGd3HZnmZW3wU7
KAUMhTPyA5RQLZjSI+1InJXHcTVVoSRcPM04mLbmOyrVPFgmu5rFUWTxg3yM1d91OaJXus0SjTOK
okL1gCL0N5XmfMiYQEIdnEfZjQfUuhS5p9rlL3PQyTbMfJ/X1VKahzPHKyYAYWIW6FiUUos23Fas
Dm3egx1kVDmJiwq+t6gPyluBLZzqSe14YhpKxhfIua/EQSABGRtScYz7+lGq2UFDtC8x/M1a2s6t
iK0MQjkVRERxX196LmdvoK6VswLenEmfXI9tzd9f78HLxWiAjQuBUXMHeKWGOSD9Xpjp+ZqppApz
MRV8d6S10q1CGe6vbYZ82Lv8MJgZH0SWhKRwvbFj5rwoIfoiL+1R9sNDu7JAW5gsEff5nx4dTa8X
fWpbx2OtWwnRMPeMf1p2ruRr6W95wn5TRQkcYolMSnuznQXu+DkLQgokbGxSJSAc4jbeZlUGxOwm
pP055OGXYWmDSnE0dwsO51FDjqK/GDgpm4iGraZxXC4E//7AYmoIL7uu2znuRReu6wspifoAVflT
zEQNkh7QlKsCgIZg360wPCXd9BQzwQLpcoIdMt5frFl/lEtiuuD6u9mtYy5h1DqsW1O4PTw69HV3
jGzdoKcYzwoaa6i+geg3GxzplE6D5YLS6B+d1JSjqttNLQJ/4LbGPTLKhTfoyKOrCrhGRo+J5ouF
kjS0ypc6R0iXkM0TCrf7Xnhj5ZpsHvGZn875uOba1ixkrg/2cfxexshwOpP/d9nYz+xy/GjxbKXX
MhyBZLQxzRHiooElSOs9B4ZURVUW+iT7cR7+kmWpThBTx0Eb9bjnOYQNh1mZe/AgDZrGT6vgfSA/
UPpxYsHr2MhKYsmI+Zg2aHWHxQHIZMFF7G/NZjB6gQ7ym6AI2VHbrr7vNXmMlDhScTdwkLhNMCkl
ihZ+6w/c8nctBd+Ts2ajXfhLyZZjw1zfWYQxocYzw3jKjczWPw2gG7DsQp4QJcesJjnybngj2nhZ
fUffLapzCqxH2XXE1v9Dm371x2yKjBmKy/NrKfby/lYRp3YH31XHE/aXm3AK9NHEu66rB0Mp9Ji9
GwpNbQBBI4QAUtu2oAmi8LEG8MBhpSprXTZyYxPmzrW+hWgqddddjjaXYalV5TBeEkVzZF8J492R
qY8N27ADV2RhLJB1WEKf+B3WKbFQy9cJY4aS1N9YuoBHN4m5Pz+dY1d3ROTam8ASioW/RLgaaavn
f+NqVuDRFpEkk2LdnIivjQqiN2syldXgLE4BSWBwD45cEQO06mYRunpfOfNy1yOD6P1cmbl91IEa
pz15O6xwE6K8gkNpFq6Zc2CwH36TKK8kTK251zFD0i0lW04ZsCqLLvEOtdHCiFJnfp+Ovtut1C3/
ND2E6KsCbJYIlNKwKNzP2qYiIaG05vM0QWrGQCbYU/oL7bUg/RSEKKbY/8QChxt10QZioxnAHRQ0
ZRojcUc2OOF6944pr3lfvgPCRyWxGmFxqhLY+g+KB/gcSphICEJdd6SebHjlHZ/rSU7HGPloArcG
x6rw344rhq6/jombbimb4SqY16N8z6GtuWL24Lt9m9mCsnhuClRbvODKywl5IiiddHK9AOTOc5vg
NKFXRh6AFHjKFXOT2/ZL8aeXSPPZbIEaqIZ8ebn+suHYyBgbZd5d2YpSibV53QcdJA4fNxJ0VunS
kQVZxgQBqMtlylnpqR8zTfligjU80x6k8oSU+SUWQQfAQGanF/0NFts/JmchJ7vbu9cSTz2Vxlhx
X7ddT2mGz4maWrsTekA/vBUNLWq6+DI/+EhjuKVq2Mfof67BufklYeiL/GAduQOuup3f90dOmBG6
u1MjDRnXvhVzNQsTmXBIoeRBoiwz3oyk5Yh6rnt81TMJmk9q+tg60WsjAFRALc6jAcD+pz4Jo5bm
/ti6JGQRJHQjWCqS0atdcsWPF7V70kkefPexZKo4bdW3uffupgLcvcEpq9Uk3vef0FbfYA7Df2p1
qLa2Wgk74x+2zAPZT9lqyt05rSRlMpWqO+3CV8r/sbsOlB+2DGtLWJRAlfD/+lrqZvV6Q6uk2TVU
H7sNe5TTsIH82z70Xh04w8PUsGrZykYvClslSgcjwc1BUjvqGG7hJvR6vG1FtILzz6K8/kS0wbs9
FPMeXPswM2HTwSNHmgPkeoMfh/ia/iz6rH0SR4NU0PoI+E3qon3UFzxwnjnVW4UanIwOxiyqAHcy
DY4aOqOJ1TJQGF6qAWmdn+sGmrJEvJdKPdSH73hZH6eB3EzUITzu1RivnnA9994v7omKB3qzC9HF
Q1xiqRF7OvJEn1YxWbm7vNOZFeEF7U4krdKjP18vwNbKPc4Fuf8ez6kk21NxD7dxZ2SkKGjZi59m
8XYFSsxzw+FFajJDyEJPKSPeUa1LgC6jzA6G6lZBmre9q1bFOI0KxgbG8f+vCcnIPtqnWMG1lB93
/m9Ig96iE/C2Og9AMZoh252DUSq1+iHUJ8JCSEi349iG1Oo0u7kn23OjzOz7rWh44UsHbEKlOK7K
VDlFdLgwVY9Dx7iPPhbtnPGts06WyLxToaUbiXuhU7Op/4b7zaR+omFF4sVYRbM0dopQ2Am2n/2I
e7yCS591iIaHOBUixw9rxqlveqHi5NYfZE6FqQ9n7uEOM6IW+4rGaZ1y1KZAbdV5HqAwk4KpKa+B
7OOVFZGPdPJjaujj9ueBW5CrgrgODA5Ss5B347tlsB9I1QjXeb2zhg4XZcrpbNdc6KzZ40dy1/xk
JJPpZRASygxm8AWplOIPIvWrna+v9v8qnhx8ld6Sum/lauJm+th0F38fp55vOLEwqa1/UHpi9fDC
1eePIOiqnAcBfOBt4Yn3whzgA8oSq9vQ/4tx4YzWlB44NGFqZtj3EvP4yeIeSAoW2LrR+C4FT+FH
5N6w0tqKHjZSalN/IrDToVE5CyoksHOBoNWqCgqK0UwYZAyMRqhP2MyyIXl1cl82FJ4ck7i/VnBq
vp5TCh2bpXcW/WDoW9GoHEDsb3GMfZ/gXolIwvhMBgve81PfiASiQcZU4sPAvfv/SX0AaS0JWJSH
xzWuRGL56+JDflNvlleD+PhGfPxHq3ww6D+hINyvS6JQyea18yiX36EInsfKfxSiSAkuTfH9Jksq
0C3mY3c4s1D2VRJ7i0ThDtrrnExp5BKmgS6Cvu0Zup4fkNxModK0eLR0wIqFlTBhMJT4ocO/QtK+
5EN3VsJ4KBFP7CHkSRxgumckZxX8w8OX22GZ8c20TxR4JcHzZ9j8m+XHmYn9vy3ebEYkuaT8Q7ew
KGtQVNn0SEpiWR5sM73V9JhNcxJJ9n6D7rSU6oPDZLzeTKNnFUVTEHqwWHLLHEMi9f9cBg7OSYT0
j8PRyFACJl9au1k2yjHXHfG73uGk5X+phOnthkKR182MrHMvfqe/kpMZ3weIr2z7P4v8aRsMMmCI
nvYxN1PF7RCbBkqA35O70qzxFUqZhVeVkKJsYQQqUaCB7h4c2UJ4hSHy4uPfiK3tMXfMbTUnL5/d
4KmMZj3w0Oh6ig0vOZ7IC6CwCgrjiZKuYIx0eqWr/zdllw4e+K7MDNTi1R4fTrxSxEM04bzymudA
l+rWNThAmfaBLprajQvfOQdExkJ+e5lUkQHuNci1C84FpaJVN5duPM3DgQeCZTTH/aSHM3uVLyjC
CISCRGYiYGojgedoPBUeAzrVfBi1SG7qS4w8Ra29y4jKrPcr6giixOC9GvoXzu1HBEA5HegPyY3k
HkyVM+JawWXE5gldjQKbZ3+cnp5lbj+UXvOPZ72vxnRsUy52cAOYtixVDqHpOLGFIySP19LrLr+/
Zd8VBRlKrIkeS4bgtQ3fbUTZPuw3/PQRHO/q5EzDv1Psi66vs5z6s5K5H3FIONtG5Cr2a3eh55Ri
yLrQSuaiHq1Bx+dzZUGLuY8p1TG2a+M20HTWbrTtN0HJYZDwWxNnbgamNiAzHqmKojQFGfJmpWwR
Z6nRV8UbwKsezn9thBYuKDV1Ez42qXYY3tdENTvkJiNn8YdEWH3liE/fUOHsLctmnJKLRcBRewHf
ol8z1tyAWLMn3iWogYeKXwJ/lu1N0NOLzEoTLghOItmvcM701pZgHYq4MtCtj5cwNaLiUZyKkhCp
PU9O3OTyfdbntltNPJGiMOqgVBuSteKCR+RfrKDj06lKP0fRQCLFEJvDdsSSInYSpL7qzWocNQhH
nBbKNAf9/xsWo3Cgh0SOVe8Czm+7X0Vrs7drK5C2SoeK+11lE6x0ZdVsr6aABZ0W06GT0SkWAdXd
9NcDxoQxmX8Hjs/LB3WW8o6Ra5Vb0Uy/UJTASelbpuxg5ghtQPVip9MF7cB6N+vVaN61YzNwmPRG
gUG42O8bx550SRhmbM5QVJDYpxMzlM4aYiHQ3dwfL+xSJ0gQ9Qar4fGfIGQd1BrQ1RWuTgJxvj6B
7SrIgW/rDLw2R9JXjIXMgLJLPzwv8wmI1pUpxDIit2kC9tn4CH7+iMLG972OgXQ5aQB1nQERHL1Z
dJTKskfkfdmqQ9BW3cJAeNzQzT9MugWw2OrBQxUxU94ppNX57Gr1wnZlDRJLYyIc/kw0AM6lfyzZ
ct0D96yUqt+9p5f7knNyzK9aMXZVNvfu7K7hd1K4E/3r8/aX1eO+doDp86vV19Y9g7wChFIa4a2T
XHtNqpuF72VdXGGwW8YuoRW3swxw3gm8LlnFIpM2vkK1gvTqJDzc++MIuWvL0AUE7uLn22Ux818I
gISx3opLb86zS3Xgn4JAiVcpsEXgzCoCm6AM/2hQ5q6Mc6L3DskvYC3xGlZ+0oaLFusD2/RNrxXs
cuGem+C1+ThUKV7HiEaW68QYxvdJw/UuqAyRDGSSKhjj3pvWH2cLs9cJsCEdv11s1tqwXA+ksxXr
Y01WCvy/Accp2LQmXdY0G1xUzouPxIPOoFTip9COKwlVJes/2rI2umhIE8G/codLEDyGOmFLQxKz
ab8/maLyXIZoJ6/Og7gJQsyu/b5vDDmzgvdyn9+r31n22lVCDtNya4uGCAtpvZVaMpgwr92n+YKw
Sl8tJAoWcNJeCLjnKOSzNoJpTB2srmwu+p1OotclOHNkad5kJQrgyZ9AJH8KOq+ZuVjdx35k2Wvg
MQuqEnJtuF5J31Ir+kc/3Jk4n0y8q/mAgJ3CQZExBkwPs2T49zqn1jQ8JQ3rFnOAj9Z8iuT+cHO0
s12OYqiGiOIAPiY2gPN0EnJkHycbDPQytpePp0w+wEdVAA27erZIZsI4QyNyg6zJx2UEExyxuGuL
ehiNc2E2BQcEyPOnis1FNrzYOueW1iX3GDNu/gnbb3Tt+gjtuo0t+Bylpbm+nrCbai/o7hYSNa7+
uGayG8m93TPti427U5KM5HSVd8rlIZrP2ouRyXrmY0+kc+oNT26K5WLwUVqVVMLtLe/HJqXUA+ni
kXzgeHcguz+htV7mpQSTgZSbWkwvBoW1qhx/cwmYikraFycQjAegeSWDYmey0UISDw/ixEgbfYrf
dCTaY60GSx/5Jl3zQJ9s8+Tk63vAddUm4vLxb+HndWdjmrS6IBMMMyW+rMazWk+F2imi3cQ9d699
2Zu+TYnLp1Vuvg+f7lRJT4FhHhRlP+sdL5rGID7kkRSDqKn4dGendzzIEXuCzep8+nDDzIEqYJAf
tueSB6M8pQj1m6Mcq8LOPiP83vCLn86n9cznr83SreLO8e+2xmuW9N9aLraFxAs5wdtV/tG3T2L2
DyvTYtidA/ZG4QQ5XnUrWWx5vW83GT9F0hJmrVppSAdcfpRyyLCehCZ63rIX1+SeABUd8+zqC1kz
ZWQHBZsahR400L59dFPObkC44xGIsZokIL6esduCcKK5mJfRPEP/l3xOVD/AGIjEoepnhfslwr1g
ISQ5JN6H96j1GQiE/pVryWQV4pgCqV1zoFA00Wi1EwOybtsHGZf2Pk7iRcCx+OQsRVdo3rXH6+Px
CNAswew74SyaeraOMYpPiO6AvZoG9GKMJJK9QmL3GQfAjlQtRi6d9TbkB3sBqAwU0ffkbsgkGmdY
PMcM38s4vKP3ipNQfBVmvNh6UaXLQT9LnkJuYZW140AGScCYi2uKkXHdtWnd36d0+x9FX2UJgX6V
1MQlqcTGPwYrA/5sWET8XsW30gnDEAJUMDoRKNt1uPtjRptJmH7tJQx+0zOR7fUhBTNDD1H+Hy4S
F55CNwA5I+47kYR+2DOIi5HyWQElB2OMrrvd6SnxA0+wYAhluZAQefql3K5qEkU5MD6tXrEgHUDA
SIH0fBcgLVw0M+wYN4uTLT7SbA17iU27IRXybZqaW6MVtHlZUG6gIVM0VIWLvuky3Ojpblygje0e
1WgKdlmV5OD0mb7x59YgAtKk3/dVf1e61Kq1oSHwIK9yVAhDebT4ILdmQp91BvnE0rvPafnanh3o
25rRbN6ERIIXmLqy72ZEUwNDdrQQ7aEgxcvKHYKKumQXNaGzH1SfIjgyRtrPXhMDzuzkBCjEmWCm
u0pBWwHxY6SEWu+HZRIdfNj9HwrE9PrOosNdBwfu4f4QR2Wvx/EtbiEDrpz0vx4Rqhb1FCvjqsn8
2aUb8xIiDWqAEdc1AZYmgz5d9/fSgOiLBaAs/G2H+6BVHHJ3gsn0m9PEhJF9uTEolfFSzcIK8h16
zqxANS7mUeLxnQYZKs0flw7cP9SklPgn3xNSabWKAYkQaLZ3Lp9T8BfQ5TUlBVd+wZPtdAgjgiAW
B9DB1tWgNIc3k5++iV/1nCGaJ588PHakhTONrQs1ZA3o5OkLl5Jo2dLQ5K6U+qFiH4iFI7dfzgWK
VySOhWw1GSMLB3BJQFEYixD0nLkFVszCc1Y4LLNsbyDHJ6gZTMSDz6I4PsCeBFxcay4fX+Z0CiFT
Y+OLlvBzGFgarSxJIEi5NGoHqZgmXB64a9BmbU0QF3mM0S3rzpSWqiTLlZislJ0dkpy9AGFa8bcR
rmGgWk2y/Rg90Jfiy40g9S1LdPyfunlz1vao0/8l5o+ZsFkNZ43LgJnP07mzkMDOJ+iXEIsMYrtw
KKDDwNT4uONZce9hvQtQDnowbJwmd8y1OXWtATnjFjlaVFVtIhTbfPGkks6Y9DCsSITWKz4NPqk/
Hsnq8Zc9v4Wqt879EIAeI4OzCsnflqbHROArwZtgpEcUiy9AJ8SSYVHI3Vc3zofKyD1MyyGuyAk4
kt8EvObYRGcbMUWI9FCAYiEKFxBEkD5HFsQTfmQTJ389+sVWxiNpXwfBY+qH1LroLNg7BRHP9UU1
hKahgzotOjBnbnbElGgjZNbqI7aithzniwCFfL78QjbkOynSXVcFivUpAzXWk7dNZAW3gIMWWuOQ
VJU9d7CGGxyM9oZrC+09N/1xJExrggwgevSBUKx9fa/Aiqf974QCqXO+/Ssg/0/BavU2aXub/ld3
SIXBER9TRcSEAgA2eq4Jj13P782WCn1LTJJYPP64tnzFHaskQWcUkJbayRtPunkPzXrl9LvvVJp5
ThSw6F9cMsEm/c4qqUhuGCiOWHlWz+bxepjye3mjvpdRcXza0IlhlQFubKg2sBNiso7PqZ3nKTOs
I53+P6uihD2IXN4OmxZj64afMyk1G7+Pp8zPxq8/HvyIk78UKu5c9QQk1v9JAcUJDkIPZN/+qas9
CqRaRrLIsWPxo/a8o2EshBMDclhNr00nzNtlubokIMKMTtfnHShJmLKQV7vZhV+1J635ocCz8dwx
OLVn2xC1GTFBwWvR4cZir936YkP0w4H8hOEqen3B0lFG/IM284Q5NJ4/TvfxwthcC5FZXobvw6TG
MHpzo6lVR3IHvz3QfkXfksJUFsjq7b8woNs4L5YoCEcOMZXnC7Dikl4cBw9keSUfTuBozcWSL9V1
NjcxyTRO55v9jG1Cww9/kTziu8vOLWs33C0+wQloxiRJjccYQpL262hXCJHoN4g0+vDjMrHAQdCs
X6EMKtAvJPpPFO8CoDAVRkLfc7zDdFvVaRsx/erXDGScFPQ6c99Yt+uWg83xsmMLd7wy/WZ4yo/q
N4XAMEK+SyApn/5eCUy/KdIiSrV0BIqYzjyHgIKywMZQwwFcsTpTn0pPXwZT4YbqUWokoJkAFfEL
hCpJOmINjGIVEAMqJ0oNEFj17rJvKL4n3rcx1VYCQKyqbrarGuUsd4UAbsRvzOnTSf4ZIev4wpJM
k/AI2+pLjO0d5H5ffQk8Tl7LFBDdsu+hj/K0lq61Rbr4EnGrsEDTZ4u6pc34BKiNujlFJ/oV8lSs
/P0QNPpgC1o2Ae7TXmWZZPvKY0QxpsrfbKVNUqGxZDn5lTR3kuxHSt2f6WR+ZGSDEIEMpsRV/yEY
KAY9HNICk6ICQhsfCtrHsloIiXIMwn5oC5COHjbAHfrzDDgDV4lsn7HOSxbwCso3wPACc68Q70mJ
roOGGijZXOxqgrm21SHlKQREcDsuNB2/bFUdaDj6HZXw1+Bh+Wwy1qXFjGMcl13A6LvqUr2EFkaC
oRxpS2JO2t7LkBzWeynS2fB7DT9isE98z6DWKdxq2lUxa9Lx7THt0Xj065lQ6fwtNuYXUNEBAI8I
Yeen1EaksMf6KcetTHibnxmY644f28quhooyOVGFelGaBgdDcCV5yABHWJ8Z5C+27PZomsuPaE6o
TPf8QKnPL37cl9Jt++CI4cihTjXj94eQx8TM4SWxZ3CPHa5bSUW+rzQfLzld6KCLgBD/IctFweH0
ZOdSxU1+R8G0kq9dgm8iMTGfm34195hpxwAdWoAY7U4OdujgBDRgyefPAGhcjP3zo0o8zDWcpzyy
879gjmL7D32pS2SdBNZTpEHkLbH4xFzDcZqYs8SRcS2ARMHnp9HJEGXgZR+5cmc9xqQajHWIywSZ
6dZ1WBuWpmfxBqXjhoqlpmP0YQBG/Jh+q8i2q6ZKNJq3c7OMIt5ilWbxxTCUwr4xSjUaoijMMLFZ
3A72o2iw131Ap1QE5smOMPIjHSMv/K3r8xSQsjop/j1X2v2fiB4daZW6xM3vjWCQnZDcTXHA/oYl
8y0xUZ4F9O+ODn+L546yQKRQua3M/Zx7fjgbZ3y0xcROG5kPscIhyEMG/XX8rr2rgnqDKTC11AhL
z4OrovSnXpMqGO8QpM1Y4CZTyg7qBK9L0GrU9kW6uAWpvj9xSfNJT9VTD64ssu6g0EaIgHSFN/N9
YNUGrOTiqLFl+KfBfkc7BoUtV9KkBvMBAiu6w5z/UCkpZbsmrdLapt25FqDjNlXavmgzS18xF6Ow
Xx1WG4of11P1j7IriwuDPquuFnGV4MvE+MsXFn9+MGioWHaQ2I5H8yRreMPptd19XsJ7fuGXZIRF
IRDp+HnQ4a3ISQ433iS+sOQv/Y/E5Ku6QUT9ZrSii7b8BIQlai3M8OYYOMDvOMeSjZ4L3yTH6obK
iActR5OkDF2YqJe3uIFlqBknVf0uhKN88dUh07avD+AF0z60RYEZTCbULazvD4fmeDoE3Xrikd8U
A4XxawDi4Yu+dKBMATRtZBwqBAxe/d5Q3kH0nOeJr3qnKqFxkGOS3MCJaSFIOxcQnY1wp8CkkKZJ
TRoPLl02tNVMb0OsR161BFeyVh6scF9NCY7eQSihAb28xqZDMwMTKcwFlaQZOQ9lOgoB2+DUbiXh
79Sc1ba1+l2eleHudJ1LbKoHLq2+jHr3HPC+ySvbPPdFbD4UHMquhvefSUvox9orIjBZV0fQ1xzJ
vQhA9kXfWnxmEOQUVwwZsrfcj7/6wKtujkzDEWZr/RpYNbBo6R0QAAjQRW986/N+kZUiaNs0IyFJ
+y98M9f6CuKUqeWvksKVA/ZfPMxwQSCojUgNMdyoiM/ErGQYSbQ/JcC9rYMq/8G2+a2QaIvPq44p
9jDhzHv4BYDbqCyZFqfpGUx9bxwgD67d3bE10plO3N6n0JhjxwJYveK6AEtwBMD/YuTUln4cgwop
F8e0k63ehIUJ1RCsdj38TraVzSnuTV+zTXf+UEHzZC7TPnR4D+v0C1ii9P3lUFgznm9xH9TBe2a5
MjDc4KcFy/OzkoFoCTUfpwb0nTKNjAAfi62mHHtTf4cNRnHlNiBP+Nac42ibbNkY1mMVchKsi9P4
Z+R6HBNKqGwmC3vtHQNzcbpREEb/1CoZdayFJLkMUE0JfPQN/6V6ZaBT9gjRoqIGrOuVojytdjKs
fB2I+wyfb8PzLqt2XgKIhkw1fX1TK/ynEgrXdOrRQ8EKCOWfSvASLNNA6kGVeCi6YxgzlsewEg7r
en/4eZIF+hv8taPq9UOwToewdyh/WB6epTI6cZN/E9n22Nr12FzZeRFHeD0QYpa1TDoo0LFjqeOj
AO00M13hyAi8E3+dV/8GBKaZR3b5aFkGS0zB7Y7IsB590F2bkY6DD96uijYM1VTcBeQIUbV3cDYy
Jsh6w3lEsYfS+h5DLq8M87C57KYOrP3jjnoaIFVw8vrwgwFJcWbJ1LgYcPEm/NL5B284/6KjWdK5
ba5Ch0zS0vmGn8FmTSywfFfkRTDnvKr76dylrDcwwkS+ZkD3EEyDbkrsuUt8AaD2WQUF8UANh111
TH25Y9+ZXX9R2ijteJWRHIo8lNKs0vc2vpuEIId95uoVqqCI3Uh+aEFdQbBoSweHAOZPw1CnDTG2
6RGQ4yBRxwevKZfWeWHb43KEmOk8aeZIyAtR/YvMvnGiv4uiMuJInGM3wJ6lY7ZGKK3y3kq+m4+X
djRJuwqkxM370OtFX02aPufSUZihtQDjy+6lHe40AwHla4DuvAVjGm5NLQpwUF4rDmKPqbvprxiK
FM6PU79cUVgE1E2L2n3i08H9scKK+NM9dX0tHcPVjf7fikb6rXsjvP0Wcnx7ZO23kOT0TkvEA8Be
9VdWeGoU7XA0PQyX92Qj4zijIQjqjfiIasAcihe08g7j1iBG8QHl7o8AaC69J9Lp6YNKsurWN0zn
wxwuu/rovC7oPXuwrA0syauXEZA2IuihqlVb60NYuAWur61WoKGWe3gTJ5N9r2Qt38v13RP5ZDxQ
TkkbW2hQw77+JQOPCazLMzHil4CqbRaHy45imaMR9f/Qj3VgQNwhPer43+cFW5Nez5f+qOquWoZL
pKufeBtLlbN9nYiSG94Nv3v6foNdCi0GTl0beoxF4de30MZU9pG+s3N+x2tPR+qfJqJZYTh+tJsW
OV9jWbGPDm7dN+CERDCwHLozUHKUaXAMFhlFqVzGnKekDUIF5jVLAP+Gw1wMdr1q4ABUDHwrLRsn
IEiYwi7KF8SEwRE7+xvSu6nVEb49qiiO45tKuvdsfzG/QRf9c08fMP0nUDAWAWDl3YphYhHURhoq
jNfkjEssw9ZjK9Cx2EWGUMVR8OuNViOIbFuP5cLRqV6y8fLyiHXZn7BNasuyYruaWm8NUzoQNlMZ
etGNODjPonaaDp2T+frPGGPD1yK42bNqKz1tU4qNUsMIH3ccRwazUAWuzd8GMGMmR9SIui8tAWvw
mL+ZAFAWvnvHo9oGcH9O56ewfESmOs5HFBrNyH032Zjn6dCI+/+n/EO6Fy2KiZS47+9KjwkZYRQy
0zp9LZRZfJ9l6rRAd6TorvX0widTxG3Cw4tUBq911QXIl3Ms1X3INVhotCzdeBZfMPkxThFK5rfV
Kag/QIZcn/Ad72SRWVUJT7U5eEfiP7mBRH1RaE8oRN0X2l/05KHfKsDu34UEm0ri6RQM2RWbPySL
PJ0CWMtptN+9BYcQIUtEVoWBwrgi1Ogby6pof2MJOWszeuFMdy+xLhCj++KUdiiOW7OhMvI82tv0
zDrOHB1WiJtGC05vZm+qR4blbA0ZBXPlxzMsG3EQ6TVSEywOPXlL9ItnuTZJ7F2rwUl6fQT/Ue6S
q6Xyo0bQZfH/be6z+HUnwnasfgM77yACpeBzqtLsOtwm2N8mzXCMke+GYsURzggMKzeUU30TIdL/
1D58lw5ED4OaMnkbFvFgb5u4wz5hOjs1m1IF1CiDRBql7d9ilAdgD0Q5w0vZIsXZPsm7mbRCDg52
dDXyVQyLydlP4og5se41XxU7pR2X5vhEcdjDFVAUJJcFRouEMBbf2aunfTBZklBNhT0423VRsFEa
Xeb2Ba0NHoZizDVQkM8JaJrIFbOy4qfHeFDcMmLOQzUz/+jyb7v8WtxXJtnKsdsjj1kc8Mi0ImVN
zsiPPMSb6r6l/L9wh+ZoFveSgZ5fHWD0qQpVaaYFAYvZ7eQslq58VybdvrIMDUx/9xEngJudU3iD
RWglhzGijrL3aFxcNIyWQJaA9APuLtanu/jiBmc/MrPgOHqKDKup6Ep1d6vrbwGwrJLk7swLLe/Q
sF6VCLQvwHMB5wsLzfZRySTJt3jvI3TwZXYM6C7yIpZam4B9d1FR8bz9pGSusVLQM0+EitbsTe6N
JG6OFAT04J2xF4tnV8S7QsOEPURYrUk1qxNLdBt6/MA+1zYgQtqgYWQJbnvoJb5WH9IPyhR8BTy+
EjqSvmRgxbU+QRW4fuckX2g3gf/pI2bsFeufFy5h0HNPPYK17W17crOqRLcwrR2zN4nArAO/FXpz
d/A8U3I/Qny43UZPEFSjQtaeAk7DHApQKceK8qBCzbuiP9FE+XC+o87U2u/KY0rk3/j1v3wNNZNY
JWcl4+gvJbL88WpcRdfVOIITbxkDvJLFSOt1dFcT7Bm5e9T9I8KD7aub1qVyDadPnw7alD5czh/N
fxgD6HCmJeLS3ub+IBQci2Ke/PvY5B616ra4k0Ufmf07gr8z8djWUEMPoxAedJYt+MjrRLHtikXC
a4YM0i3lqEQsGkcFl2BQGVFr4HLBrQqRktIeda/M59bRLvKcIuvqIkhp79MVZdlfh+Q7qYbgB1Sa
uHskNet1FQWwLA8JXk129PfAqIFcYqDwuOxkFtD07v0mIvmWmZWkaugPvj51s2rE5UKLHs1J2X79
9Nmg+GmmUmwJXVzhVk2MXWSRcL42FrTdZlsOnnIZlDcHPWRrgoxV/UkR+tRUO6GzLvdKkGsPnSV6
a22TTrzWfoL0lyCb2Iwv8LA9QCJ2lv41FqoFqNDaOdRN72YdXq12oEpM4NPMpaBK1jCmPFDrSoj8
KPMA7qWSN8rMu9Mn4Nc4s0OBrTQAHoBJpjDDeokuJizXANHhMJF+iDFEVuuKgBLbIguDmRv9s0bX
jGC6Nh36MI8TVDdWBODlH68kRYRtTnscD7eBZIY2Tv3Ye3p1Yk8oDX+qJviKjKZngurbIbwf1a93
evH4X85isI+OuQ/1f2S9QA+R4JJvpxvEtE0FoWk5vdp7QZp+VoMq0BVneVdJv7T4zOh65GBm9SDS
Ho4XscW2mLG+AsudTe/iV4BwvDftll6amt1+KIGLoyJ3TM07g95rDSyrI7oeQ3s8aZWsX2HVoWa7
1cxyrmm9jxnRUi1waRieK9h9x6xOSbYCfhUXT3TZCk++X/JEGpOHj48k88rS8VZBeB8mzzRJuTyT
g8jcUzd0AMTfvic6sTQjOMjZkgbXMJJyalVF4mB8OTDsCEpTBoGDerWqM8z3YaxnVNq4EoDFuRWm
YKGyIakckL79e6iArBicWaITm+XgYSNK9c9evqJTDnUpaapCky07ep0sXw8LYmUo8T8GQNOzh/On
QrPfGe7GOg43RNSODr6tAI+58Wp2Gjf7lsq997tWQckaXnfvrt6PqAMNvR0HfsxkyQvs4VYahKXr
+tNBA2BinRrL7ITAXgBHArBkXzH5TKpb7FaL77PGYnkWZ7FQTt8clAdOGFnazc1yQdGQ3s8ZHS2c
h2csj8ncctNeLSPwc/9K6WJxg9eJDy0B4vRQkzJ03vklPMg+Kro3uhauWRUbH+To/u0uBClT7zgi
BNPH82F8MdsKaIjc0sB/tODlATnaU/osYVNxxdo+MJxfxwgHSnuNxI3GyqxwlYMf0piUrvF4khtS
jBAMqfw7umtbNQV/kcoEngRk7XureoR6SStN9G+s15poasZEoWoH0PL/jx3PkicprgBS5R5XRvYN
UjgkWEALSHARoSvtn7TZ55/g2GTJTcJstthb2Wyw6XjeeaNK021UiBb+lSTxZIlHFzPqmE0b4Q6X
OI0PQN6ylgd6bKF76gzoPc4BVQCJ43XSrsNqy4Yr0Z9jwbb64kDqEPBc/yw5KNnRR5v2ZBj+RIsU
EboUIriuvCCHFK1d5EDQbu70ntlDb7YZL6Rquez26bl7qvpLy8P59tjl8FLmcOnEh112s72QG3Ok
mD7lYPb1yPqcIkm9Y++8QQxl0H+8uhYUpSof3aPgtqL0Rvi390SLViwNLCuhlv5baUYFONUNZqVv
1dun9NSpdPsNrsy1TtTXtPVKrzHP0zjOOGrqAroY/c16I57Hyq6JRpVpw83EtTKgZ405d1x9LAfc
nFDO2ok9QjuSwBkFNJKwtZVRx8oreFA0a/dAVjr/bcFSVQcA3/YhYfs07NtvZM/nUFW3CBqfOQbT
C7OSxGfl/psphd1QaPG4/iut9IVMfLnBEIyFESyGJ4OVDS+ALKy5Tw1F9eE3e0qFUOPx5IiakSZd
h7y5K6TkXgRJbI34E2pQhWNkZElNIx4nMW1vVBQ5Yw2D3Ycg1O5p3IX8SmmB3va+pK8IKHyAOb+F
eK/dliIeaKYvsiYDczfokJ21da1Nhx2Q1t6AvJQR7Bc0rIoGAWYtgv4N5yKX2gfOpjFWlr5pu+SZ
wc8QH66IzsAgK03Wn3Vj1GMDhSI1clBQ7zkAO6tjs5/jcGFGVq54jIIqGYQb6VZb0rSE+mcuyMqx
quN+i36tN4VqErE+isUQljt0FSspWMDU7Z9FZBw/TxPKv5NZCdMF57Po6RLYYlD3GiLBXx0gHA2q
nlyCaUrlAqwnbHecSDo+R5xZcsV3qLY2HvHzhFa/0Kiqwb4gPDH/4TF/u9LKiGr6RyKiksyCsmpu
JXs7WxLGsh+7o3rf9VYwCKcbgcYNi/loudAuL3zBUu9z9J/Flj5e/Km8IKI1zKf511LIUl0DBhSM
WA4iiG5cS5Dgb6dtpf0LQOwag0+v5y5TIarAKUCVudmtx3D/FA/iCbVAtaJJj/f1n2/gdBRarDAl
hlO2BO9PrqF5kEABdGtvc9NvW3Hhc1bWbBQ5GpM1zTISOxs3fHHQt5Cu3ezDqyUN3THaQT3sGnB8
yNF9PiXVT67jvuXnxnv03qAq80xJKPM0eYng1CvmeubVxmM05bK1Kc3+Bh2pphp/56OZliM4+TdP
6CIKneGUyciUL/t0j5fx1DYFgFQjOkPB3jlFmYtD//QsWeg9GyspMztn2BzOVPp5vvSXHnjb0sjc
pB3LmDlVi8Qwkap9f/hNdZw7MgOOgnc1y9Np3XLNNwmCrjFTK15Q+V/iABoQkuKBblsxbwW7zafW
/89kJ9pd3lt+4mxwpN+zF4IPhvAvuygryIvtOKwOGx0Ix4cgt6bDS3Tylcl9rcSWTaIm6PuPFQyV
I24TDsVPgUCnWKGY5sFnHj5Xt8Boadu4PFbTGJe9bm5nXs879LfaanSzVRR8GBPr+6EEzNbdH+Od
ESsRd//+UF1w1iYlmZbttBjt9sPWroaQqsvOriPiHC4tpKvTKL2GPGWbOw/bVEyKVCtkARnNP9M5
lMrYihOGKAotWyWqDFS7jiliQbqqGsoihOJx5pBZv0B2O8LrXoXaQ7DgJ/0ftKV+iv7BXTu4N5Ql
td5+/dfSuzS4qPswTdmSdjNyUViQsyeMbp81HdSKxOLNhgxyNeAXQgbqm+aAwxTOAq6cMTQBBSOw
qbWq0AOSpk/7TnFMpMHIT9wYJ4ny0HXxfMym5/bWJp+kcCHIAXJ9874XhSCxdcfIhTM/+z+wnL5k
BskNVV7IQ7XSxXrAPb8bRb+1CZay/5Hjy4jmE4kfkBxWonGf6mxpfhoQ0i+3tICs6Rf3v8h8EHkF
j4VJTvJE5YqqrunwpS8m64XYxWAHvgCvz0xDqLmz+5a8XHkcp4Skyer2LGLwNT56RUeuF4qnq2NC
Yrqq15r1Lbgnx4CMUpyqioTD9gHfu/O326AlBM9Icj+ZE8QQaUeUYQ/XeSmfhnn5Lkwj3Z+NXt5W
TR5kOAIwYeqzCTcpZN7p0uOhq6k5aimtV5BhMOu2utQ1jA/O3O+1rTizLHv+WQdqlx35p4e4gOd4
PneFMApvBMgMZUjI+1mTRronbO15RQwa4fOA+DmQ5J2tiiXlJn+uLD4FciDrdyz2bKMDOTbCrssi
2F7/y9m/mRmN9UKF1vI7TGqx/zvD8EaTm/MotrfWW09pady4TZZ44fYOgjx04j7USJoLRNR6rXo9
EmYXJw79VEdUOo1w/QcMnAvsYQDr/AlrWWu8Yu2Jnqapive5v11vSY2X34GH5QSlo3+fpNYb0S1Y
lwCMi2FkSsrGVNSE9tFwCtwRDo3jENsfCuoFiEfLEChdmcsT0/EbiP99lAI8AT7lIqx6d1LbLQQK
1jcM5SDR41WjzRJKGetBRi7B5wbffwKNzCLdfYrLDiU1Fx3oDWA62j/zZlaJ60vd9C8rmDOPGKHB
WdVat6wLlekCCtMY7m32DtZ4YEGJc91zuvEDcwUahYIobu98QLolESxOKPKpMyhCFc18pQ4CnERQ
zQHaHgdLu/p3AD01GgJ2fAapbrPiDoyZPumw84ogZ+4LxRgzzPKRgDoopboCYrc7ad0cSeE/Vu7X
QGL1zGgyBjKNjJU4J4ezGjvJ7JST3dd85SIuLw/TZlPgAwAfESyVShliWmTJbJy6XYaCoxjJtm7l
6bHsR7uNfCcUJ+INAPCpLLY+8znS5iQqDGH8leRQKUcgUqGkXvwoCqEA/J4zdFQVo8uaEWGLIo5r
jWwx/sDYlYTqDtF7798e7nOaG5Mj4wgZvZ+WzlGe/nFqp4q1BM35/eYOYB5Fy5GtyGAnKbdt+z2T
sTbIlvr0LazQ5wKAnMK/EwF8PBKR4v5DeyLcUdc8iy8NcZ/H+999MNqWZzyGUzpdSYaedORoz0KP
XB6OUVbPaFlhGNGVdJ03JRX8L+vi6+EKidteRS71UvnA28mjK3cQzFBBM7FkwajbglMR2WWlVhof
cuNoTY5Cqdda9Y+oOYePlaS9EIut0niw5GWzgBwun9ij1hK9zRrCusP2SCBBzBdUTcsubbu/OOBn
MFSjtYMLFIX7V2ghY6Wo14VpWV9TWlcx/sdvUb/JP1YSHVbPQNOmP5+8HbdXIjh7YeyaGK99FKIF
FeEXeXx8ebVmHN9i2xbm+A2ahVQoWkUnyWqF8chiVpBRjE7IkgJViS1pTjAnb7/mVZ948zvioMIP
sRm8lnIRSCejOQ+B+AMcqW8HB5hcfTrVo6FoWZHoMtlj4B/9yehBeImyP3k0A2/QvOzOTIMfaKx0
taVMNJKjpFHW2vvDwKhF0eBO/PPgZQL7B7q5z4UlUVmQhEpEA1f5vrv+YHDWkK7orS3J92Pv9Tz4
W3jJUc4+cIVw1wb4b5CXCETi+sJ/WFxOz5KqgaKSYgrCUfXtkq1ksIM/vRo7da1ubiA7VqdCe6DS
BlezRh5l7Owf3OrKrKX+vUZAKkYiesIeWH0nZ17MdvbICFsCnuQmMlPR1ixzALTdB8IOTFv8XGKZ
iZiCeCuNiFzfSdTmxoMVGH6Q5GhCbyoUdwEIU8/ICrobf0fPsEYOmdieUIVT3nMK2Lk0FWir2Y49
j+V8q5J6u4s1pqb8IuPCm34UM6/Lfn5VRQNPgI+7GU1ruogo+4SAYBIabJk14iG1nQf6GPayLel7
c0NgWrfaUJvvAdzq+Bba1x+3ETLOqDHB3bSVEwENNsLYFM4l6k7NJN/oUd9ltI7b8EGte/1YmIPB
JM7MZ+8N2Sy5FK+aVYxZ4Jwrjpnaf5F/ovKaYtmn3MMFNNQfhSAXf9xdY9X71ULzVwzpiTALa3/d
6NUxGsj2SqjylbsmrJQs+KdlMSq45Q0rlInFdcZPz4mEp8ER0/aD2rIp8bQr7n9QTT2sBRCFAnF4
Tc0ek0lw9OhNN7WdmxhimhxTAxhXRieHpUbDguKyuJnbxVycmhaOLSjEeI75c8Y10jT3wNcuNqJF
ingAO39LtvuS8U0WslBTt+sR0ObaNWzYbMiZQBme7FNBOn8xVE7l9xilRDxXq9eFx04rsIROoN82
yqiN8uBUo74ESQyEuY+tW+oKz0/ipjQU8FRa+e2d7kAjUMPfER4j11Qr0AcRPaoozB0niRRB6vlZ
+o+hUg+S6T9oYAqmN+y4V9gaq0T7uAOnwHWRpffN+s6kR3F4T28EN8UfADvW2HQbBLJr/zEPKvtd
iVQirNo4ly68EhbR1v+WvvAPIlE1ovn/nUQ2nfo6hB0v45/YTsLNM2+QpU/KtUHizsha2wY8IPrc
PecxzepyoN9akpCMPi8H5z8C0YL/aVrFHRTkJ2hGMJFBBO9jTMM+2sc5n187zs9xlfbMkwqQlc/P
xqVgRwlB12uSCl3Sr8ZHh8xWsvzs/G18NPaiifvRDcnjHCYVqRaqMA7il//0+TD5DX5vZasGSKTG
Gz7o31DcMRBeJ4JuLg5QkvK1doFyJqaYpR1atkY7ivDwitqJzoCPeUnjH0Laut2BtLLyzDpFBhws
x0y17o4/kwJfmT86qiMPqa11GLX3tWjEV0vGz8n21j1dKA0dzd6FT/iH203KZdBL6q8xbgIAM053
xWHQWmrpu3jvdpXSC5lPhqMLgZlgKXjden/KYsHobiIGbSSed9+vi/QaGuJq01psD0oPQVJrtpx7
rCaVXJIzHKAj76DRx2xDQGrS5pJ0FmCbcXzA2vPOGgjVMR2w++eG52UaqufpinmAALLw06wV5wfx
ewvCGtOsndT/WBACHAw7Tifxh9JwkuElTnEfXZKfGZSyCa+uD1X0oG7EsAlnhlNY1zXv17kTpLng
ewKuLRubA/3zv7Qp8CUE/qjwOcxIltavlIBTf28PgJ4j3nZmX2OBLCV7xV3AvMrQQJPIk/bFbw82
rDqtm/9i0zfMLqhvuK6OiLHb8NX0qaotWXIq49ElV6QiD/pGvYV46mIeLXFrYSJyc4wjV/V/Kuqm
VyQ+m2GLYVP9ImxU2okZV5YEVOCNSPntl1Y8QCDhoDzP0OnN+1gTVitf0u8rAhkznv4SPqqaGOOW
tzSES72uK4dzg+nh5rk4q+9x8f+GrHit9QpFBKxulEJQK9Br5nRxDi4c570EnPP4RuAfz6WZ/oWV
cY0CHzrn1B5W2GRDFTaiwihFfBJjaGfww0h3D7amFu25R0B34DoAQfylPBYwOO13Qn2dogcvjicZ
75bLLugT7KCRkucIItBkMLOnvzNdgwsfpwcdCtHYdV13dMWvalxYlp2jcMoqPdS8Gg0OKLwqXfjO
uAXgMRWznQE7OKc5yqmwLJe0ejRfBAqY7x1WNeaetMzm1lj5zAkbS2BcFR6qMWciaMvrf6gTItf3
GNtmZKQVJ4UzgZBsy0uWG3MS8YSjggyahV6rXGn6SMI6+NcNt8OdtuS0yr4uWtbfvBO+HfA5xpej
V5JDs0kUXSLJQ0vTWAlpbybkHhH140/jCWcsJAffiXvhoi5zfVcPoFHZzMOh3a7dL43LJf9tCQkW
E61AsBNYc+WzCLMq1nOyQ3/3NIg2Eus6mknd4vgJQWlNYfHX70WcltulcwQuhwV+GEZajFnt+DYm
O3kCutKDagi4QkAXlFO7WFk96kaoJWwTjMqt1efBHfyO5eD9/xMEbsbm2h9A/y4lv+0ZOaqVcSBO
H31V5CUyTrivgU/ambRXfn5npLQ71mv3kVvZSEKsOtKfiH6rUMTZZLQ8j5dP+sGcTibLSVHf/run
49Fk0cZzwMqx4NrYlyzXyVUbt18UP6RBihP/fuKpganR4GdxYVMP3MlO2KialSYK3QjlyQf3G1Rj
EC1i3iax0lV0wxpT4mPJOD0VmDMwGQBB4dS4dgp57stEnGcc8IJvkNOQV+AWEHQP7yPuANjcsLWS
bHSMnafIefaROn6DhltsR5U3adEqJ/KYpeYlvZZjTvwjbXva/JCqAj4rnZFz7bYjxiHEy4I1wmec
7g9W1zO9rFzuyrl2s0nOYWXybK897jURJFd15iFNWr9uar7C9LaiNFl4D6eC7H5tdItg5FevjS9q
fTJkuBYQJx/1BW1jaj9JLcWO/BieHKGUpsKtafp1mN307XfNImKbN9BeaJPztj74CZOUrRud8/Mp
VTFqKNTC18Zu+mAS3whe3rbCpKqoQCk8QVMmcGr3rHsN5S5ikLdX8+H9mNfGT1GrDtMAVeufiP61
QaNgSBkrOy0JJB0Kd1nfTZ+HHZG8D3s7R7sSwGau6NXr7xkeK1SpTTc9BvUr0PmHO8K0LivnCivL
h0nY6OT3vjRl5uVpMeTS2SWgRpVx1oDqnBbA0UXi61ang+iorDrkIW8HbtX6n19JxtXy80MVKIzs
448Adqc2bMuEKGfGDl7ren/dE05+BYeon9yohfaVwtADE04utyNwmFvU1RFZYCZk6tgsM0/wMPEz
WwsYIfz2jXdJwiewzQ2tcmaBqOahhMbLdXCpviUmJNQRe12zsGXyxH93GwtT2U6Yzd6JtE40fWk3
3hnGOu/YBi9TA9b9U1eLCK8rYNbpd4446SI/S4sYYFItqOzIM2mmusa7M/5rvV2eo2Cc/FmOf8Ge
wjxOLy44pMOw3Tc0uLw3bXGESDXpjQXTrQ6VsOrGpQMR/fBNRjTg/QfCSe81UIdntvWMUx+rRQ1q
4ORRTBU3T1dNunZJJgI9t3Douj64H06tgxiRLcmxeZVMkFXwovqQzTGESWnGZsex4r2nXksfMzo3
gPotNfXqwb37+IXkWMxSRROlKvAYOdn2yYaFs4PAO7hUfU2VbJcM4HHwcklCpj7mdI8nnI9ElpBq
V5AefP7XgGdipDKR36IwuheEWx9rouJekNASdk85hMn8jM22ifysHdnPuTF8nE2cI10ANBOklslv
qNSnn/6kBaa7kmqKol1DQbCqTTUrXv6zTto9pelQedwXpq01S5G8udRPLArje4Q12nBWmc0mZR7a
EBkO/jvaasC3DsCwDRK9d4A1molZsxUx4/i/SOl2xWBUXbpKF4652AS7dw6LIFYh4ldv7NJ/oFdv
I96RbR0X8pghmcQWK0EpA+BG7o+6n8H3slDGOy0Zv6F46m8ZEVFwKO9iBwPDwyax0/RzRi49PxUj
uU3lgN3Pi4Oh09Kp11qeahP0sMX4i8rsq3dYkBqIapxguRkL0nYPfYTDdKJgUdRc/0C8JTu354ke
if8IjmAJ3U+H4OIP3K0VAzr54vKdkVA/09kf7F8WrRKnd2WLJlBvi06yg4vrZ7qqydYGBtIJOg1N
ZkyfuGvIoUIk09z1w00r9gfD0e7Xp3jiDuHmfliVfKFUIgwm0cFVoolJKG+XEGfMAbOIPiiF9bBO
D7YrAveVVO2pLjEz5l87T8l5S12Drg4bxV4RoNq26KsJst/O/ewcltrLM7vXVVzCtEHYoTXQrt93
x+k6Y2cV4VKAMiB7N1x90RoeoXljBJ4cvDfgqFqf7Ifjl0klMkAYgg9OVHH8dnUcXh0eun6JeWny
oGbUkZxtqSSExOQydm9xm4WhwwOhwNYDNkMKrW/69aQY4zUdYyVaKlq6CRvgHhzIYUSvQixwjzIc
5w7MICcpcGRq9Pyn9PIteyXNeHZGURvQUwu0uBZ7MbMtpBHCSNSzI2O0SYzTzUaWGKi7rPy1wMfX
dudEQf7bGJrL2YjwaLfFm1ahoYUNo6lYAkj9uI+nP8D7oZJKwIFfNhrtaqmI41OqyaPudexp1ctd
/Sqfb8gG4OKlsAXkVj466+6yn3d+fBv1IDNzPwlV7uFgq1wixrzP0KyvrJODIvBLN4oo4bIbu4+w
9OqrssBunS7KH+uiTyKGbSlRRfiTiTW2+338RsRyLYupDefYKILOF6wBHgM1gzheQuTVbIW9Ka41
+LyrgOBxvKEGQNrRzj3hwAenxRET/eO5E6P2qnjkND0p9vHp1o9dCERqfDR1oip9g4VAbLrYUsCI
BRNir3Q9zuasrju+2yN2NaUO+Z2hMLeSigull7BBQ53y5wt+hipM6NF7PkonAFqn9LNrs1Gl71il
Gmw/j5+nmPh5kiCz98wohAL9DDF7v2m+Ndr73u9Baxf7KXd1KfkGZH6sFvu42vltigABtvx4rpnW
wjKf0hlBxG0CbFTfqD7UNnOz3rwx5BnxMGMyDM0zuDtJMFS3jfHVD7BcNfUMoVVAdEchh29y4jSU
+/02ZZ8mHLcDrTX1rz1z1jO6qdk90nuymLrkMWxHGASGRH4hXixlsO55F4AAak1nv/ZOO7OXQqfy
hteqYmSCc7hM2WAIYi8Jv4XBEGh7enbwc/J+B74la/5+Fw29pi5SgA906PUZsbGPHjUpJRxPd8Nm
169Yjq5yHJAYrJPcjWILPlVuq3gqGTwlohPYjBPNZ5h2DIBAv3UKrTboEB3K2AEFHvE4gEAc3Dhf
TF+5gJ+ywmqcVGtc/FvwSOkelBm9uPPCSYR/SHZhaGBLetDudoQ80QsieC8o8d2lWj0W2bLLgULC
5uB1xrHgSs7eB+taykyvhtkOh33+UeZTbdqxit71+2C36jCDfLY2l7Jl1nHRBLGIQRJ5iAhQvY+V
nUzlVvD3fXtWl/hfMWybYvVt8XmjHnFNCQolst5ErdMWbBcOacMP0Fo0+gMfgBKuRa/ixPBU9aJO
yMQ/FrerLolvf8ctzCrapIEaBH6Su819EwAV7vbIboARBghoZQytY11MCzDVVto3SgQ6+YXYMS6Q
ZPj/DHantU0HOFGQep2vbGZJLeZTkKUN/pit1VgO8mKXo779niW9V0bp1O9tjbDHDKSspfTLwO3m
kpmEjuJEJCU4em0m1ed64Hyc/UjIHjVu+uF3EEygdrcOeNfzxjl8+4faHCLpM0KEZ7Cyz49QrpWz
69wbd+vUmfTrhMj9yPu0skUtwhPy8c6qOvrQJh3N4Sh+3hlTj/lppaBwIx3yibSRnskh2BFujNx1
ERIQdKnTErqNngRLJSotpCPTzZO9QURyaGCDNY2zC9Rfvx6bP6EzzKCTZIY8hsOweWy9FmYuO2Ih
xuA5XJttVq1Whml6CbDkHLX6OGcMLkKgJxRHx1cs6sSLG83hSJf6Ftzx2W46uFIEalB/2/m7wOTA
9mGzrlSHqzUl8zYQ0hN01CCmTPh43FTOE+rwGEZLQp9JaTd5Yleh4Mtxm+Cs8D88pFzV/4EAz/qa
t9Kz3NUa4hV5sLDuE0fq2RQ2vL5OXmgqm6ePclxbOcLxzAzCRA3CG7yjVfwBfZaoZexkqq0/eSr/
IuDpVpnyGtioNQwE09Yuz7guGwLSTy769qQaga9zCqLs/pPtQ/SNW59lPzv4hZzbpONda+1/t9EE
kXE0bzmPOjs0SKeA027r6r3uYHYiGJkoMqRKRSqAYGsH1EIN/CW+nPoeNn4ae0GmZuGhmaU4+nba
xmx8JQ9VKP1GLqkI7c4BuUUfRfghK2cWU5dKs9UP6wu7vi81TCeEInJlh61JMKlMtH0acBPNppT9
PSc4xXwp5BQZK+65yr90ZaXEshWhMvanZwxhVLKE8fDQ4Q7xwSOXrt1uEH6zhrKn/LbnKjkmxKCO
goTlzk7weyIFWd/Ccxminw/AA8inFpO3QUFMLtYRTVR4z18ppaDFDKKEojtvGOHcDe4/zZCdnGtf
65/VHj/uROEZt9VjoUKKEeV2WGt3JVScMmze65R7IQcMDFyqcV6WTB/Se3+7JOYL1YqXtjI1AuL5
CdLULZrQeCOFTNnDROYuZpnmkrXGAH5JHxo5V1HvapjvLm2WtipmoXV3VAPODjEYwj4d5Aj7vJbi
CQEW3occESTzsr5nCnN8VHeIT4DVXKBiGvHzeJdQSmnnuLqSsC+IMgf7yamI5nEZB60d9Fv3fVj3
n14Q/5TLYUY2ys//1kHI8Oyau1wfOLdb8C3AGtY8+zi/a2+TETcnVNeaF1ha92dHVCmg5L9YcwDd
UAenfb/Ajp/fzd8q5l9dJfm/rg31inNV2ZO1KcMXq6D7bhzD3LEDB9nMS7jm9d6aF7NRTHoKJSw/
LtCcpgeE8zfzmwThIKRMipDlZ3sE5IWgHUsz/O+Ofr0Va79CZGdF+imY0oxtPN0FhzjMMOSxMcg4
EiezFmPpqVUuTWgQRRoFao7EGUi3meDTUQWlY/JZhmrg1yZ3uq9XsudrydFI/DBvm3qhPiC+wdmu
PzqKYnz7suF/dFZ/OR8OYGL1EwVZXwwTbHQgO0VDMOE2sEP2uf4eLwoBK/zhLaSwIn0IK1dZWHps
+ehr/VpD4WWM9L9kOtoBvOZnCl7jDYGXu4QGK5BmR1Cl7z/NQzj7sk1cVBNZ++S5KCaNJq6He9OK
/dlne2aGiJM5SxC1gL4vVKR9BLWAiTyNbRhy6gY9x0nRbQOSJsP+EfthvHDVpUXFb0xTPhOPqsL5
Q9hHf7RvSmAhUbMZWZOrnD6Rl4T4x9kjsCrglsa1TmORSOble6I9bNb7RWqP4RLi5SmBCepTXkty
ruQOge1K5jxzcNIb9zX7zcNZzk51111DB7uIWvT9myzMdAeNDFGNEFEtySzx4XqODKRduBoBZdEY
7uUSMpEItpWo9QQ2I5+sP58g4WZw1jR7YY7TkqHXNyXPOEfFeJwuiurQCFzrObIruJ5k01t6wnbV
Sl73gOg5Yg9MxcwVgShNoEGk/hJ4xf7Y6FOdYwW8zj6amwdju4GvEC7UOeAw7YPNYBL5qRukkfWN
Rp1JNpPP3AY0Xl3D6BXEghCHSDSQjry1AIcj7wGFUSiWxGYT64VUXCekpWrLlrG/U2GEgx2Nb8Gy
DffRrw3N8WZbR4S0+hJCM37PSB4N/qiHMaXK1lQou44y5ElhjhVzqrS3H9n6hPqE1pmwKbuAh//5
MBpDYMVzqwXA4hOjOCJgDxL/0DxcBd/G0fSUMjeDcvRag2B1oc3sTAegLo8BUpHJmT86JnLeIwHe
luL0APzrviEhCi9b6ic/b3fGBECq3D3keqsRMvwfgHkFIkaNVhQqVGydtiIm7Q5Rn+RPRTmrCkYW
7D22rNmR0dnROKONyWzKSbBltyvbc9yKsE/BvU3X3gCW0uUcvRnHwEeNOuczPW1dA661sJZPJmDS
fE+Q8pMfD8h8K7moDzPr3ur9H/Qaun9nyDFQ2W8nTyPBbOVfndDuIRm3ecOQ9L9f2e+mLg//3cKz
Y0P/Dd3m3G8aSd34wQSGW1CO1w44gNGPvJKur8hqm4pxLliMIdx5TQYRGcZ1vg9OyjGR1ziKmb5m
GVe4iFmH55UxmtHuUEl4xCjSSwAyZpUPbksZLhFm7RBuxCFUWoFc8J4quipSx8ltpsfGgy0Fm80l
2R7Fd5V4dOkJx6qzKbOIo2s4gSfthfyRxJpArYT54l46vQOM92QiRtTAlR9Px/zdWDPZXrZLpDTB
cYIcgfyspGDAwpiN7OWNyc2OondnoaPRVhknBgwBVKk3dCLXJxlY2hwUMkDziO0GE2iUh8D2htCd
4nsyM+CSDxd9qf0FpUkd5NL8sr7nwBenQcOdthIPniQvF+vRaUB2kpi9LxfuMaEEahcvGPaoWnHM
NW7LmG8OqmRmpVU3icloXpksDy6mfOE/FoHlJZsLQk9PU6mRbTRRXApRKOg89B39UA6ux4mRuovV
pUjYXFdfMJ8z2WnHoTP++F0XSJrjgqbrKnFwrotbl5N1PhDNV3PLeBGZhu73yuKWw/KX0roIuNR3
PIn7bqHxm8AK0+WpC2Otf7JaH0N+CiIpBBligix+FDjX5Ex2T50+em+uTHvI7NBv5mYX82AJ3EV2
LA+xPyDFv+LAI/Y6yadBCAZuWzzXD6V6/J2Rb+b1Sd9sAOkuFvXfnrs+EBVHDG4xNyMbut9icpbQ
V/SfpiTQovwecuTUM3meSOF9Br7eFQcv1QLil1gzttkuvlvzpA/GNiB1B5Fa5es4xZFzSDE9Y8nU
bsZltrvMXPB7l3N2HgqIduC8E/R/3kK5UoHpmtejCP1HToWPw6JWsJWEVVM2kss3vxV4SjhzmURP
w+AdlTv54ZYwL8qcDyB+QpMGN069H1SipN5xQ7zVPmnCcpr+mk2K/jNJEwtMcXEZXDepYP3werIb
Xgv9LDf++HtcP3W+VQHlo5SU65nmhBM1lZ3F1CiunGLhkxTZ0I5ycmycx9vAk5gE1TgRzkQHn/6Q
wcsWcxdNmLm3jLIRZFOosRkyN5RqWjjoB52iaqe2ytg91iNVHTbJPKMGbfIUdnXhjsTgIIr60ShF
JsxUufiBsaG13894oCY4+EoooukjQFD5Z1tns6ZaYlkxZHop8CbrS0/sw1A+Vyb9zzkrMvQ9bUvw
X4GSh+jf/84Hv2eNyrdE4EouBx3Ujv54iyWHIrgdG8PGq/GWvBHOcHC5TdOGikf3UATB5bcE95zp
GppQV9VNOHpVT3YBM7n6bM14zoQSinobUz4F8GcoT8gIvC955HSBn8kM+cmDOGyC+Z9pqBNr0Had
/+Zlk/PBEBZeWH3YRa+PdGT0x65z+F9exrJTzERMpoItHsqAfj/1aNcSfIxNEVsNuDzGwKtVXg9y
GzBx4DhyGtDKEyt99H6nSZbPZLillMtOHZuks085jLKRHHdCO7ZskGsma3weiypJR43bazKAit6O
pIaV9PwV24bqg0JSQi/DJfUcNmK/AMYMS91eSUxd0CGGrUfVY/mYdubTpWcbZiBo+BcoFMmrKeVj
F/SUaVHslXnCalUA9rxWIcShqLSb7uDJZCzfr2zDmLdHGEGGk0D+fnTPjAxZhliOIeK1E91oJIR+
8tDsps3Gv/mAAVfEAdHXeykB+hQWNr/nFpzESAnIIA0Bx2p3cInzBboA0nXQZ2mTtioH7Nc3vAx1
Vt3wwztwHXjVvrZ0t+cEB+IOkLSS0sxsXBdh9j+shXjMGX2zDG2/OiF0sd6eJ0Z7t25h+/3YJ9f/
0qr4h8v11SRfLT2ypKUpmx+ChoR4osZ+TE8Edv7m1qeajBYC1Ckyw2ASJC4S5+8Tpym/vdPSpcrU
YB7z+G/veJCqTagssO/GWkQ+DWzd06CoNM2XsgDPPrdsfFIV9LQi9Cxa4fihmfU9vfNFsFc4eHaz
WdBLxwVOxEG6XHYgPr4TLp6k7ed6Ouk73W+SsWB5vyU16VZ8YFGbAGydiyLNOwIGWPBBcprT+hFl
OON4KoD41++Vr5XfL85IcIdwwtu1ZIh8Dnp8Por+NdwvpvKJAuK49xJ2WxHonUsKMfofj92aUl9d
tD67KGWSyc8CbP25UQTl7y3DxJT1OFwD0D0EMgUpPgdkbZuea9gZzzG66VOoD1MicFdwTHd2XUa3
T/AgEAgkT6W6ChzX8OmhS8VfXJuhFZMftisS7ewdpEwPfljMf350oYrI2X45wi3WfjYZtzHSpYea
Z5IHK0XzndS5VidElWb4PgI+qhBuDylQrLCJEOmLX46V9/lnBmRLbpjEnwTssxCuW+yc2mh+NvV4
IOvtVYF9nbf+P8J/JMiGnn1i2XxYEP9Vy5nxqCRZ2ihuC07kH4hfzqA5ETDZ1fF1PWOHzDAKwok1
XiWMgHxFdBX+xklwcGBSJ7Olf5q6GY0BXCX2TptqX2PoRl4BPxmvrS7mIu6pk3shboJ91Nd9V6cJ
8rNMH7tm3T3QvBA9x9W0CgChdSIgDV7j5AcbEWBTkK0dz1AZTO2FkTwNB/s1duygZwtkwdS0vaLO
FcQV72emUIgZeYE8FNaUmZpoVh0Qk3iQmlAXC9vgLaR7KDOizJvfCNPwD+Q8gekjqNAK7G64HBU4
sh9nLDiF0Ojzer0vd4fRaU6De1gyN1lq//jmJpUf18LKz+VPBqyJNk3u8HS1ZzP+/fRCmrIBZSHN
znyMUvbXqd+RUCBZY5BA82lWdY2/bogos5gW4QuPF5Pyof7SWQz+1jYjMSuFHzIX+tdDaskNzGg+
ayJGubE0VmW7Et+9uScxZ/Tc1hqFrY/7HSsttg3MrCz1LJ7Acn6SWv7HjpTV/X+zvL3MC1lhuTJn
ROdOSsAkVN9UTCALomslAo1Fx+TXVAtMrwlReTr6k5RsvDxMlqDgAGmVx79tWAHOrzIzUIXvwe+K
LFbQR25eBi0hVST+tOHZb8LcgdXzuCZmvxiklgrr8xUUrwOiocV3bjnniuMoNoHzINovW+qBvrrg
EqDd4L8azhQX6Bqve+TK9WV5dc3Ww/8nFkvs9TzcbPPUrNTHpnxETGiPuyIqi1QmsHzKAKGEEGiW
ZkIZWb3ghJsiF16zejbUy4H5xlUHV2jIVKyYnNVVBpm4O1ODjCfN1QcpJmVOlZvBVEC4m2q++8N8
vqCy1zURVyMFL7Eyq7I38dLoIbvFN088eXQ1cQUPJvECsE8d8WWLBaB92S4hLvLzPoI75jqt4Ews
H7PVdw2Z5yYDqWHZRrN55pNnrtkVP1pr3acKKUzL6FhyLQI3ZHCV5VJJmAwCEeh24blylwYk33j6
/zWJwyD+LCKxahxc5Y8hRt15miQBJHr1kK/2ogof4TL2X3GE0cU48T3WlYFEhmN6yms/Senp6Dd7
e7Lhu2xcyvoZUvYb8SvNAhG06JIvCk+qX8PKtAoILgs4cdpNEfFozeAVkH/PirCNL8l64tJIPGDF
UVWSHNqlBwmMUUB8m/2YgbritNWvWUCMyYVTw5CmWYtq0fW/SO/DFIzTMvdN09mCfCYVpFdTJInz
U81m+Ioz6X2GUKRuR7VGZvq5SbtzNotg3Mh86JxnsCs6DS08iHA3bAe99/IdiTSOWSiTdls2Vh3y
UZMv/ewNSP2aaMSdC2GB6i+DPJaBPb9gt/Y8yINX95aNzSMQ+vCZG+N5kNpXqNyZVlUUqU0BO4My
jAOgx7bKO4wdkDey+8yZNVxSGFmqrps0LbwaTpf9MX6Rp5c0Ys6+TO5T4vSudVQsBuA1XpKbCoyd
y+3xkYE39Q2EjYEvxLqM9P3zqn6m6WDsYLMN414S26umAkJb4pgOnfBqf7Q5EgRlk+u9k5q+UI5O
Wijtxlqr2EB0bEFtbylc9k7OSwc7UacJ59FGhKEvVmPJtbxox+MxH1Cpp8wU10YJHc9As+6HNQ3/
5EZ/V7tL51+JLRKJiM88eeLc/hPJOh7nRw/vt6fT8t1HLggMdA7lFee1KW06+LXUhQrA172LnX9N
GwWg7lIUDt2CPCcJv5kn76l2F6LOTrE9gp5M75XpRsyXQE+iXx8cQOipqx4fggMte/ip64VojkKn
qoky2R6bpYWC5qqm+yG4p6I6LOSYDBBo6XRKT7xpW+UnektRS2yH616JTqg42oeexlVxta/UPfJD
ukqmAXpIQOLGAf4EWZR6IMS+FYMXNLbn83naKs9u6b6uM3dWrg44UNecum8OfBMUWL3HyO/fOqxK
hKA32p9zCyVeTlckvhBeh/kQAxQt0hZxeQ4RAe7zXYN10LOzDy214fMUT8dWkXt0Eqhe1ZEb7SCI
/Qo9C/KLHhUMabaUynuc1D5q+bx3yRTRTiM7k5wVrdKzM2gebOvx0yDa5cQix2VVElSlqUB/k7nS
5lqKRB4uozx9z5HeZ4Uw/i1VVlUOfP72W788iwY0+sU/kgixfqBwIqB2FWEl3e1h6dsONZEo6DVG
+V9l/LjkhPN4Z1QHUc2hwwtbF7viUZmWtpZEPU1yOGl6fcXcN22BgZ9VuqzfTqW1UDYcNV5UbpYn
spbYgPdYl40vIQuAadge8ZADJ/vLI8ZnqDJVHKfbcvN7dvcatsjBaCao2E23gt9f6QQm34Kt8KJU
KTiaDxeBJ/uQm87fIoYZJKCWCaSl3HEpFi2D9+YaL/ltcOoPE5c0QUki4TOpf25pC+WjuhnHStnj
Kk4DwhhGcf8u/LWN9u4vqv5vnpkn9SZlRjam94xVTti/OB5LiCaW9hS2i8PvOQ2ortj+8bdxPpGa
BQD8Qm8Oglw82sKfRGtz6wueu2FiC++x+qOULyqKUittpq1T0XZJZqqlMjcWuR2dU1wldczJcMLh
8WfJIjrUcxN0JpGycSaimAQQtz29vdnqxeDEgLBaZh13bx5rc5uJUDHFfAhp/6MXF+BA15WUHd8B
P7pgjvUiOT2v09SYUCBbCqvt7T9MHfoIZo2Yn0eb0987O3xgfzFs67u6DDNQLbEFFOHXfSZn7izy
z1ieAvY+smp5o66T4GtnX5cdtWHK9i2HnRcRh/R+eQldml+htArtpsUrR+vSnr5NsqtJ4PSccKw1
9paxDmRt6vOMjRIc5KfCTYBm95rQeTTVLO617iqH4IHCuRfi+SII53wosFkmVkwimX5+NWdRYwrO
1Baf/udFVTrQ9lcq/Mf1Bz0K7jw2xIoPNhp8ppYA2QxP8oatpDKtRtX3GPKTEMgmG96qJqlnSPX5
EXOcOFclXqxiaL98zy+s3dYw3sfaU1ctP6xqbVu0dwh/vQlmc4Dvd2tuY5O01Z3mMMmdtfIy+k7L
hFsgDpzo11lH5SL7fpJPsvAbpT+SsoUeOPftdT4fR4rSp/nWpAUYwbKZsdfyJy8wJi21u8FHSSXX
k519lrl7iU3XF8d1fo0oMdZVWmBFjGBTW3va7jeRt02iMIz15I2G6KEGaP/ubWYPem3uCK4RrELm
un3v7eECWQw/oti9DbcsQGkkCV3QMvM3T3sgh/uXk3K+707AKc7Q3sfLCkSMxC5eOSZb8arGcnl4
AXWoCuzv7BgQrt/AbMXw66Zmbb6yc33EBXyDPaptE65jFwCOepsDMbTxFpufdbuFyPAoNSOpbsQt
t4HgsEM8MqjPj1qHBEcItuDQlaxC2n2EKCMOD6625oUt3am+FMWvo9y1VVsvSTGuBtbumK7I8JW+
ZfsCIX/GOO6495igQYHViYZUiAUxVWbMdRJveB1enc3Ur9LedsE6exa5wVHxH0Dotsfme2zyApmZ
s/ku+z1ncfcEWpcP4TL8rOYXhvAMr/XQ25WuiybQWwlIrwsrf6uGZnZME5Wym6uZ9Dah0V6GcfWG
efNRs0Nn9weM9O9BfXWzG8BvccBx0H8IgZ5M8Vn7A92bBwUFlnOcYBB/iZydkhLpOE3rPgbN6eJu
ckMs/f0KFG/2NyPwz0+vVtIdEpQ7fsy6yjV73ZhOKnlO/cbJpAA5f3hYPvDAJ53BnKViCeEP7iin
o5UuyRkpTS1IVqyAvqHnsm4jaH+quKwXtUVndNF7ZqFjCOlwmYqlVUdsRLvLFeaXX+DWQOnYAMEK
Rvw0AmUKA4vimI4HOSpKn5ebHTAkGePWguvJ/arj1i0czrmOI4LjCQqffWySNTsoxed35IV0pxVU
34ciDQvQBxBPmGj+r3prvQuVAii8KWOMiOCvg1nDH59kcgLPdgWVJUyIR0SyIjeB8YaJnnP1UXWY
oPT+o/mRI3WWnOYODunPNGYH7aUzI6zMFvJHze/EehtbgRfgcWJ8FnSuvQtnJYx9Bk60/tIuk/G/
p+OAtsr8mneFD53kzMU9v06Aw9RWmoACRHQSNiOH1iF8lmyp3t4mUY916n1UI9IcB+r5/3g+ql4S
aPjO1D5mvWLn90Q29ODXx3HE3TxxelRzxdRPk9efWiaFUtmW19ZUSIBPoRroZ2YGBz6ToKbMh9tL
RI7L+4hEwfRCbry2A1JY6bUBhseLaEIcrwz794y7ob38FtjwkF0KqFfXjA5uN0HUq73+y7/ClK+A
24Whb5JeAbVFyuEGvZsapDvOY/N/pJwqzXvEKNTDleBKK78xjgbWlyhD6kXuMLC0sWU+kKHOXXxK
3Imf9xG4AnF4S9VSHbKyMTGhEW/u7ktgEN+oT50m9v3rPLBYDaIqKFYnrP5r5oaWxgpCAvTjQA6m
gsLjRhHzWWKx/qvVCyoKcmew3xvMqL1hGcPnT9aHvt/JphtdHdyISZ4IfONFdBJcjOZzO6ieX1H6
geU1ChkVvvTBw5jsGxDsJvnKh6zCBNgtM4sf4dAiUY/b7ZDdP/zfWJxWYP8xWUetFnHIW4cFTVgX
LKRzW/KxBJNvFosnvkbg3BcDiKdLzrmQDV3OFNULVAVym0jT2OlYNQFTymVbmUm1y2sFSjweW0wV
4Yz0kLMAxjuKZlsCbU5ZhTi2gjf548LPlyvCKfJsaxdkrMjcwpU7ra4j8+9l6J4Nfozz3zhPZYWu
DPuno4vsHu56WghKrcRjIApOEarpuBA8XA6PO17PtYgDP5G+1QTfOpuXCjS5gD6H77ZmDEqxEf9g
mODlmrYXFe2l/kmRkEtyiaR8j33kJtqUm4trFVM2t6/dyRcWkNyGfPCDkcIBd3DV7Xbxlyx4oNxi
qQTfBmBDONOK5zkYvrV4TZ+/IZx+jAPZR29WyYGdIUs56GrYkIV8hyZtWU2Jw4/nkNoXTBmg1oC9
6ehA3X/3wKG2xuumE4BXgJeNTG4Zq2b1oSD/tSGgwMkY7ddGklyH4guMpRWYABDs0wXEF8caBwYX
z7ngFt5IH3Ay+lK7ycRLjUSt0+VNqGpiuMmongXrS5CqyfkJLPn+KAeDP/Jce7yr4W0IZBeISjjo
+igK0N0YrdgIFhUS835bdGR+zp8Qqi6cNnlTVaaL3uqmEVCnBmZ+E0yJon+tcokA5U/hXPZt8/6G
PdPW/hpUhEUe4r+CoUvrrSt8hYp4cp1a5d/GHuhOeqadflzisu/x9LgOj/jZZuKbatECUqMOQvu5
qdaE/p1gFADfDY0sfsWx3dzLp538T3SLmWbwQcjV/+kemGwvcC0Vg6q+wjPik3uH0ciQQ0QlvOc/
4lYY6b3Maujqdvz4S6WkUy9GOEurXBYHkE2VQvTJhGdrqBdtyxU71LFGsH7fuLCJagGxHCiJYCuD
B5qIJEC+tUHS1HJq+R97mZE9J50aH1ZJrYZFsmSjDvmSTRK2k5hzgFazHkPVJPQejyg0iOjXqNqO
Xv7yJ5Sb6r6mAn770GN8Qto5EC1lOlJiPM0XDFWTxndN8ksdyF6/aAbjSNXzqUx++csgMsdCQ4uo
6oXiO34ayG6RXEAYAaxZc/f2IORPzoXi4ld1cVtXrw8PR8MaxLZax3omexUP7kMvZnMymTdCxsW7
BhG+F7LJTkwy2IpzaK0K/Wfm2/wuIn2La4xr70rWE0O3SEs/xxumMcfXhqQrtNwShL96gcA91Djb
WYJs/eL8YJ3HfrIn9/e0jkcsWV+IpmABXviVWgJMcNo9g5R5Oo18+7kAV3Q3ixFzNNrZBJrJpMiQ
hR8QvWiDElzjn1LSzhyHjzjaAebgWseQgPrh1LYuQ1m5kp9zkact8cL8smH1fkdOU9IRIUo/T63G
UPnBAaKyig5xaibpFx+rlSwy9GzwpsluatZ4ib+r9zObKN3ye6Zy4mg9zN3vWnkZu2k/V2YSp1IZ
2nTwOAi5FqiaYmuT7VNvj5gk+6P3V7/JlufGmfpjUVfUqRfxgmtv+AiyqUnbukOq/bSDMdJMPzEO
14ShC9Q5DKPivTn2H4HKHYhgE6rI8OJMOus9eIRM/WXs09Qie6K0rQqX77nlttCLLy69QIavcKWA
1rOCRcmkdA+L6zEu7nqdz/DH9nbVKJPjZJXZ8X+vgH3aawvrhxMAIeO5sW7QYE7W3LQn13BDfnpM
8uWlbz20EI6yZBJFqF1/s0PM518hYpRuqeLK+jfHBQG1yPiHdCsZJYns0dT7yz3ezMUqdz8LTB8Z
sRq2TpRJa9uGyhNpwzZjG258jHt50/SsdGQ+ZiUDR8MEsgxE3okNWiMXOD2Zpq5WyIaJAM1pFI/T
wAC/c58DtcooORMe1t7cMkuNPQgeneG9lOxrF+Ro6lEgbe81fMOyUzUY7XkOZo2EcSepkPa96W82
bh5Proii+ndSbaJN3eM+Iah/735uLSBq8ZzKrJZv18B6jqcXJfLGW44kTgXdvhQSrqohE9TmjjMG
GrTyI4v0VvR1sE7hN8+ECosHzliTJk1zdez1pdQeoZFQcAelyCk/TWo6P2uWwYN+h63NI1pcKCUA
HV+slaHxm+GlEUHuy4HhKJwwCi/6ovRwOYvGT8qOiCstBy7ix7fj1/GMYWhGYa//AfyDCe5PvRxQ
5pY4fTH6ciLod8XQte2h0bc1RuqXMr0rqJCXU7d42uGUkq+YxoEMXJBVACNcAVysh8Ho5QE7CozB
EdXZU47VVM1yeezWy1Vg6SWkllzMCseu2pNalojRhuWUh6d6Gchl15KWoFJYiUq1e4Xuems48Msk
ZkLfO265Lh1Ek8V8zHl+pa28jAzec3YIc5yEu65OEDGaO1xrUCYDkxDA+iBU9aMXVw7izgF/Mfwn
dEZ47fweYcL2PqULG1xHSp/d8VzEjDKkht8zyPvw6L0VZt4QUtx7cfrgNGyF/PtWeFUzEsO/YwWO
OXds2BScqu+PuJ1Xbigssjc+e47w77NjeF/ndqtdmE0iYmlR9UUBDjdHyBTtCtxZRZVie/NQ5pDr
XedWNlx2hVp5iDKx0BVoKGWXmDRjvXDXbKnGdsjjZU8pJEMemR29HMvH6Pez3yDgWBFfy992yZwb
uRY3Ua7XZDRZVa02TkgMwmzAzHA/K48TJUmRlz4xhbGFZQwSLAm3VTvWPpqwlDIXOTKFbD7Vpgx1
IL4GwC12a8P7NaYt4cyqSqz0d73ZTMx50sLbu+osDBqEbfkGg5u1Sc6uG1IJxrxg5TvUR0rLZ6s8
Hu234/H/v05b1M9auujZ9bU3Ik7ldDBJ1IFExMN8sBdfHHaF9iOXWOYfbBp3mdNAS8ml7IACPWx2
45HFRGdyJByIX52F9+dCUa1seqq0w/tUTmrxs5TzSYEKfgmVtWOq3fk0BDO7mv2RloLoOAWTqIki
JXdIEXBSKDLgEAAT9kmT0zkRynqKcMpoZyhCMpqHHj0iPKgfw9izqeC1yz39crL083ogAawj0VSq
ywbyOknYXxrEdCwehkpeuykCl6XFhMzTaDl4aZECBGZRZOYYWYY6DDO5+N0HxSJ5hf3/QQj4fx6A
vLcdJhL2cW6i3v6ESS5Ba7HyoqiutJG2pDvrsHqpOMWz9yVzeyUbhooUJndLJpomLpKg+zP+Cz3Y
r1cXh2yk9o7ZNnw+zZ5Fx0gY28zAYJwJtJmB6XUEPVqY2BjYEnWzkq1GDilhOU4sy0xlZyFLu1sr
lEZBy9I8A/i767kpiA1KPu4N66j6jRW7ItgmfjHe72RAGHoE11Yw70k+RbHmP/bGzXHQjqaePXHY
9zrq/Sxc9dOoGftv2qHt3G21GjbMZ2ngTKv4g3gob4+7n7/xmuM836+bzaOzrhzl6KCWq2rNpI3w
5da/wx8LyhPtyX9MWqlekeIfHhfkERZpn2I8CPTPT97wPgEMnUg0Ac+7/8jp/ifJAn5cc1WXbyhO
521TQX6VjAQair4Zb6IduYcqQoOgKqwitSrLCYWMfpmLYZaOD22JdmvMnl1/Di1esZJErCDvpR5v
ymXv4/Xj1S5UOoY1q+ROhwVweRNko/4SZWLUfuytPlM7avx5Fy6X3oXHqUCSk5BBW1oZgMLWX+be
uQ1indXgyDWa+DyX0JCSj0w7cXgbydex3gsOI05pMWpLgQYIWUGgIQjQakvS/lTcOlpWIvoEGqjF
x/0i/mKl5d5THXBK6cA+TTXobNFZANTsDCtTQLcpEMUXDy1BfNrOuYIUxDZ02DBiPFqzoebIYj9G
QVe67IvR/lEM4CtnSB+8lQsLylfmB20/4Iqvv/+GzrAhkkOCXrhxjzp1TQ1RuHCNNjBlJYlQ5MZb
N+Y0pGRmh3KKRIDQW6Wgf+tc3Q+7gZKmDDZr5KyDMu0jGvzOWQQ4fUQjGPa5VfAZn9B+0pYN8Jci
deBM32gKGPpFQxIdIKaYdtdClJzYEr9igYnLWowXI/Yb+vr6ntNgJoFiKcK3Lwm58KY5Gzza4Tsm
ATev3zIlU0/nN4bmjkauWEsGs5QPq88AIUcAkJQdoYo3tOFzbzu7+M+2IVa+L0BUHU3rMYxjj3tt
qiog7c1/9g2dpc/K3MDK/BSeZhwtkwLCoLsdRsdCQfdwomWliDVNeO0P2VjaJJeNwioPK/l2vVXu
FpYmM/jhqZOXz1TWx47gywFHqElzXn1WmGZFDYLgB91ixaSWWPsM60VBk+0pkSIcRO79rJaAZ+eB
qJkGDtDrrrDyWyi+z4Ppgm7hDggH0zpSR3CXnicwA0jYKaCIFO+mr/GubQAXNtbMrK4alTmYn9nU
pefz26F0iAxijezJQ1YujPK2PSo4+TvLzEVMa6BPTP25VpBfxNDuuPMNoNtG74Q8Fi9pDsngDfs8
YwTGIbd4UpX/at02i/gGyoW0K1osB+y0MV9RLjOJ56klWLqhtkwahiCjWVCdIBjN6eBk+tyxbmfe
AIA/g4mOBU7dzbrnFrRM/UxtYMsnUii5ezJwWmTCK3WDP6INhm+CvfyqXNaLcHl6LxW5cO1gTpLl
OY+uuPuRhqf5t7d+XBR4eC1rzmTdj+i8FE+0iIQL2s3Q9CLSu1KeMgCzfJfZj5yqgmFeI5f84FvG
8xCq7ixzX4plwF3HLeBNdMD9xU87SSm847EPnTyrfo5HBMU5UEQ5jzTKKocpjdp5iy9wdwq9ZxDm
91qRSdjwNIWnTq7ckBw+FMn4VPhqUJslAGcn33sah3X+WZ+q2QMcuDnBfTWYVjFKLoD2+nysnAXk
9NErbFVjT/3ClRpnh+EFM/ZT8xNcJGkXGmTMWSlRSqXOiwUugVic+CyOlnCARvvS2N/sYXxGzsBB
mwiZHHQ8A+uFf1NeSDvVkghOZuEDyTrTrFonuC6/OStbZth1ZS4V0ay3VULUSJsBqASyT3f7oMzs
GykTCxN7nTJxayQhAB54Ydg57jmXInMwLIfRO8L3EiThb09djLWoldsYdfcpYWuVB7JLZEu3DxUR
kEjDNwCBs4XlUIhCv6SLkXok0Via23/38dB3enKX0VMVn70mA73Y3p7xUpUzIcseOaREl4Jdaqb2
yg/FhwnHBUmXiLHe2E/0OHv0X3OETaNB0KBRTBL9V2n2e979fNN/lF+Hq+bKUWiflaB59hIkfqkJ
mX9ByaqMmIuGnxlzp2PUswk0YuAbzG6bkzssPUtepCvaQWCrXGUSrhEhN+HCEYuErCjqA6edDujo
ZzutMqnCj8M0xc2dWfW0GMyvWDEDxlE9p8He1MtfNF40dK4W6K41RrwQHhGKaBt6L6/7PPt3hzjP
fJxN0XFJlkr19nIe2uwTFOwR+IHafBOz0XOeIhZNanJ9gr2H961CcMPsZbmAhGCFAGYK4XpSZHgg
eTQ7sBw/bdswH7nKlSjPkoIbNU7pq3PT8rCIvvLolViiKD2wRV9aZ7NX3nl7d9hrG3dQBBJdUKpp
5xXtGFbA49WdIxvQW6NfeWevpfjRJZHNT6esXxdxi9bZP9wnICNf3Gl1GhfIj9XNJmKqQ7xvlhOP
hJcD5nGu8J++izDsyOlb2HVoEgyiLeHtv9/GqxNZ31HS4D6+SWH7xEQQlhNCqeDfJR8gnV7BqRR4
H/yDKqcuYOfbYp3h5bhig0iseccm9KVWWPE4ojunDo2joNJtTHehLEQwEVzRxSECZoN+OSvm149o
iVGZ4emBfn6uH7JKm27ZT/mgHq+HtO2wdK4CYGruFLuNEbUQn6meyS722WdL4rljfmr5ZdsVyfmy
Q/TskhSS4LOu5GF8Z8EFyYLg3zn3DvbqUeIVqmSih2fTdbbiq+eJsXu+Nbu/t7YFQ76f2UMNaeCg
IfJDwOZhiLg27rzvws/8LN15AGeiNx59MT5VN3kVDSB6+BPZZ7qEnMQQZ5bUO7d1IVL+o5bdm1Z1
CPleSJ88kv64lQvBwTJJdrvR+I9puphFcB4iHuWIZ5+f502ribLyfB1f7ErBpKFySIO2A7/LTMeW
1r9SPIZ9k2+i2nC8Rt/e16i4rsPiVuG85MGj6fgeG8MEwLOKEEQRSG+HugvczKH9cHI/z7QyZ2oP
BAbmr7++wNGM1unEUo4D0Sdm+mM2JXDNJkPLF3xGsHPHvLmdA8u7Bt/k+Fn1t9NtM0X11iuzGIB9
q6ld8Py++y+uf+F5H2SFcRcEy3dO0tVpozhWZp9QDJ+k3e7/qXTkx83kaj9BF0rlcexO39TkhR6i
zK7EZXJ0otoNZ95tt3ZPM1BYiDG/fy91dQJabe55AkN1kD54RYnqBpv+URSpLQMmz8SSfFWU7Lw5
QuaxVN7vkj5nOamiLSDwz4yVDlR75ILV8Rr9L6os6bLOq0JOlyS8n3m5rqnt70ybfN/HDgavjaDg
FPbQhQUpdMYHSC3JUUUV4oim+/dlKs9hcDwg6iuXhUHdXtsQr1mwyHyWUuGpLKH3jtF3NBqkoFLj
ooR9i2Vm5FtuZU/GGxjFUU4yKB91uLDr/bcmIhw9TkWHp32f57HjGOdO9Fm1aivDXwbUZePrtXwF
qzaj4JXNYxKIXVxqhkNZo8cB1/AfeMT0ubSa0JQZD9wwNiwOsDhGdSrQqik59XjMj/h0qV/wdwHj
eFVFaQ+ePpzKYFgvkbWU7l9lvIpBMFJtREkEW7/C99To9q9Lgz7Org2GwGoEw8Y/nh48UkBz2OYn
bzdFP6yxsEVbun4ERXyHiEoOsSrEnl3X5T4eNfktfcMpsnwc+yf6diaQwZfuelO3NEzNF/UX07A1
uUzMCBDRcKjxC0X/yRQsYfxcyUCYDOuKw98hVEpxlXr54ZDcCLL0fYaLozaEKXrKINDWJIiCMqzn
u7fiz1K6nKenV3POfQSE5kvGVLAMmXbkBZcIAC0HJF5dY5KzjWAwCmzy0vQX7qILcb2fxYlOkWVy
JoFc3UssWRaZhRQB7YinqxpeH9TSeIyf8KP/1NeaZscuxgvAbvdRbgx4z+LhmsErxPg8jppNN14S
nC3Wxj3hIzblsm/vRGiU2x4ubJGlWCkRPtIOS+aVtJsqZHBxlz7nM55TRfc4xTHZDjjJSjjR5xqC
lIVKUmyrUcwCCD2UyICVYWwWTXVimfZLJUCL9NDs1jLEA+zdZz7ClB+0aif7gKd+Xlf1nB7DXLze
L/Iu9Oo86aydLf4zovKVT7ipFRc3Lpo9I5wIcdyyUnnlUDuq9IlnA6hs1Rizpj/yr3QZNVa4Pe2/
imyjHeWiaWZcER1uXlqykRz7iYrcUoP/q9orFByqbchSaQ7M16KXFzs+cDfBJzJPnh9a9kc877yR
2aXNxAvbrWk8Q/SLwsVBWUTvJxlnbWs4yeZ7kn8h4IEExR9RmJsHvRm9Avo8SD5RPoOjCBeHtQTg
SwOlZehAvDKmCXjdYdEO6QNfWBjkbeRFI5LmbgbiGiNO5VA2tjWYgT3LVmmwyqhjQL6QV137RRFn
hbaNk9vY6ZJmE8QYZEUL7hoAjg7MxgyiuO7EDxeJVFZ4k9Pr6g7ECMFDwU0Cv5igVNpXj7lzFxgq
D3H9dQZyl+3k0FvZ4N1uEid/rGtaF0cR+2d2WYyMWNIGvtuUF2uwaKtg1ieIwoazYSDDdY7jnYAL
/tFrcUZk6eX5UiGZWc+WE3gEBlMMObjHGsJuUwBnT9VfctYgdk/0jE+uZ9n98JvLyw3ExGzMaWoY
sghm1guE7t+lvzIJ5jEqbxTzmcc5iPTRCg9peWGtoYhZc7vrnCwtQARlWoubVvrH1pRuyVito87M
RsvH32B+5Uyn8Wi7inzApQyLXt8Csh9pjPCfIbZVllwZFFjIMzRY06/KsbsuZb5EWXbD6cnxY1pL
cjwGNq2PYb2Jc1tc0ijrC8I4OAE/Kue2OEErkdiK+otA+6L3gasSMVGmgfMXTTaZ0AQlcMS+LHru
1PpCUPe17vpAIe6ybgSwXqUCevIEKAme8Ph66AvF59aQr5egQ5fRrWALUy1haOY3Rv77lVdzryOy
aErP8BKUbSSv/go604LnQtSxSWW4mDfxVQuXp2lm/gAzuecrb0pWporNAWvVHQBP8ruiC1V3LSpS
Q8kAQ+bXAJOdG94rNQHROCEB1Vm8E1qiPSuptbnxZnztm6n6bXt2t76qYUgrbJPkxU7yZGuqHA11
j7NIBBZC+A5Lkr18sYzP0QjHygOA9LI4FB7hRKeuNHCv2X7qBRjvpzbo3CgvAxcPZjjQsKJ1umkr
uSXvwLawbBWkGpb0rNxPYwRoODpqEAxlzrngJz46/s1D4HECaJ+/nI5p754Hm4fkB5BV90qixbqA
0fDpilzI/SUqskEe72jIvIKsKXyQ111qqljwGOh6vXyglnCLn/fhfF2vWku4v2GsxdCi/TuIMnHW
bIvRdZuFs3VtHXqovV9BLvz6NlBXOQORQvFK4eE/QQY6EHo4f4bQB+ERklWbFDzNi6S3eD2ZSlHd
rkx7ZmcfgQPuIKORQMoOwmuLHrUe7Hn4ZNz15hVkl9I8QY8SQjMW5MF5GElFZkgTDuBs76KzAg7W
LZfNViJ+eAVL88ELVM8BEzxw+v3NieVgPEVwVYvTa72kNAqUMqhFL6P3DdL0qL74yD5G16uEv2Rb
r8Z7BZr1LEEMOuJeYvLtCtVWS6PrlV1DfbhQGvllSw18RZCXXU6wZ05OMDYy64S4B+fGHNybMDqp
8EWaPm1Jj0A8poMjcyuoigwjZi4e4ATfBKFRYK9l6sVnv8P+TvHip1wgAYlUx+yfq70j5HQ100iB
qpBttHTgaLtLkIiK8NHNYXaQln6fP6gdy2lVQpgQqWuqokLpFoVQUTGH0wCKSueJ+O1PZhJp/SBu
lrY7SPM7NrV3E3cEftwhIDbLvrRWKBbLEL0jHTc0xr9dTouyeCPuqA79A+7Wx7aje4rvq9BT5MqN
WP7rmBOF4Mq+TJs9oZEeWIDfzji09g7dLfDAjyMeMfTQLMR1fOL4ALiCUwth8usOBSdAwqqh4fXI
vjhBZ1uj+fhXV96NGiQjXO1b3peeEyN/ZCQLcbseNmmq8ecZ663uKWoxg/kQZVgBIBYfvh2afkF1
LOuTYOCKS+i/l+GvpQU0o4H+9DgO5zWgnif8U8vZe7PeIXQDUWSEbgtI0g5q+pio0rJOPZuA2Qg0
okOkLgT98ZuIE3lwV1fcrBoOrzqvPv/gOASKPGSIFPFRFxwOOaEpHZJnl8kT6ieiyPboEXvMcjyF
f9+6viIPC0jJG9YYi0mDxx8t+OxsQ050V4u369oo5PMkj4gOOHjt2xlAP1ARl9qAhvQs8sieRG/F
/NDsc7lrOVPzkpUiaDBKx749uxesPOL1IEzv0azFcEP185P/Af9mMus2YKtfMOMNBWNzY/ehkX8d
9NoU5legdId7V25SP3acaysJbBmLPJ2DtYuXoSTqNs31XGhpOsXn2DOaPqRkM6Ky38DDCis28oic
4g3x2jRD1egP96aVCTEa2DBZLWD/QyMaqKP74NJn0ND5qlFCWDUadC1NI22q90nVYZCS+85IwRuG
1tnh1ntJSlfnkdeSp6LECkTSclyIRgqO6pmybosAMLseCgEb4wEUWvNp6BkUT6bk0u65ECZ6nQN2
jtCB+SJJdIRmNWtpYl0bdKIZcc6TpvYzFr3aSdpNrZtmR7JyBhp0DXshMnsEsyHv/uzTUv7iGVaR
cOzJj8KHAdbDzl3bfpowDJQ1N5bn1bH7m1N3zxGNhQxwlqIW0+p25rYYMnI/1VDV68sJf0nZEEP4
FezxsSBhGKoFPohzTMMoKeTrfEs36kpA1hfgt4V+3CZbk8xBewPXNrOKIjYoKyYEa3OUadcG2luZ
AUo4VHaHDW0eo6juq9O1FR5S1kQtnNUDYQGGYTQW+bWrKgaSO5YwJqamY+7Ph6hejPT4CESdsH6c
BmhjRJLqUD9wZ2aiXCR1iqdiQXLrowbqnsqfbY9/eJntiWogdY+lrxpyMsfRvOG8E/shODmRstTR
/ZioumkpaOY13lfBUs7cYIKbCzGOFI498uM4Ee0oEJMJOQA6nAGSoBT46pNqrtLgvFRyBmX0SgAh
4YEjdCBP5C1Au/CB408e/0bY7DZINzusqjWovspJ6WIdoZ9Xkg/JWWfKsomuao+5h0jIqHcSYGy2
qyFSJ0Jb/Wg+7TZlvhju2HiG9/Wj19yHEtJHYa/6ZBXn+G0Ykf7Ya2QAvg+RtJYHmixj3VQ8VHJj
Gj1DNUUf0z5YUGqZNnJJQ2dLfSgppSADi9yydcD6oxRHynkfNd0+P/Z6BmeTC1UGQa4kvgdzG+nr
gTWwCbeI9vjM0IzUP/0BvNIRaVY22mLwmHEIAnhhjAUzjV4LvfV3OtSfJYqv8rh02G9N5WreHkeF
GuP1L2RGE5dg+Rh0sNZIao6Q0eVE71yG8IeFlxSyQYaWCWI3NMJ0g8JlAfkCqFbjNq1UXDdUJp+7
0S5lYiC8cbibyJeSRB1CgHw70AQ0HJavMjg90AAQ/QYBDHn3g2f68e1CMpnrAhvtKGQg98v9AfwF
CkkILaw/g0e4W8Uiewpgv3vWO9iNSn1tNZjko0jDxgXOkV4akN4JFOnpKJGcsWvj2CxEVrWMQwXf
WM191GUfz5opaB/3Jr7VMpS7J1mTO3MTG7kodGRKc6Fo9ZL2DwkwmXgJaCjDIQaoXCTPhHupFmzx
aNVTQeTocTT8NKHU3rkAZt/sts+jnEZNazFEMNgq4tTBjLdwmmbR5TMhT9x7mOScWlS578OYmN8T
A6DjQ3BMX3kxR66pIxd98wgP8ZQGKNyJtbru5Wi6VzbJBn/y2zrvu2+SlwjJWitkgjLOzQZQ9770
SysWN+52T1eB7mSCQNMaGkUtNb8IzgX0kib6qUekNl7c/aHW7/WXDZg4nMlBFwlbD9FR1gRwGDYT
Pyy90ZQhnD0cUZ4Dau4Q4iKylhnrR+BmmcadmSV+TvWNrvEaS+18KPhbcgoBONfyqi3zVG7Qlo+H
Bu1xavj27BePcE+nCNh0s+/CaSlEVE0mzVgOViwHEcseq2LXpRRXZMjfg5zkyI45AIPTmfp3X1s1
WX2sdh60dZpjPumr2p9Dv6Sj5MRoJ1EUPjxu2SWalx1Qx+G+uNf4LxN67ju5mycvZvFW9jtzWEBs
qkGu96eXpEZx1cb9G+E4KZ8toSpQ4OQjMhTnrxfKTil8avNvm/w7Wft3OdJi/QZBNnOJ8u4r6gNr
NHL2vFEoozmJFvdmYAl/IQ7nP5UFmo9BgG6styAtW9QQpI8BA+1Gt1IewyJwCwwUT4bTSnbuA+j4
xWAEuSqxNYN09Kjx+FjJ9km8JWMKAzNdHMcGHcZSVIf0ZGdwn2vOCRe8yDiMjv4UtFKYUm9rav0P
viTVAuwYtv1CzojuXG6YqldTSdX3fEqk/4HwY6S9/cSPbdi7Z3+kxaw51qQVGHq05h8wAYluzmxg
H6Wtv/fwH6dspaoEHIkYt/kqXd7S3B4/yQijDm6GiAE47rNWayIMv2sMbJicfjNfWCcpa+bEh/kR
G8yH4XG0hC3fzNHjUEEffKD8kiB+ccxfobskERq++zOTSQub/fmdS+F4Z0gCB/f7mcsb/94HlBik
6h/gr2PXzHjOLOzX6wFlGby5EXkthSGT2v75Rg9K6Bl4rySoP8EGFRR2Y+qSyFpEPAu0Tz7u0LCa
+l8prq6moPnFF9K5gsnb9OVi7LJhPhEz0mxnzlxcNWxBdVFhi0TZlW0oDLsY2MatFPgIORYS5QVb
Y4WSbynofirbUKhWr1ox8OTx3to+kASD2i2jBjhRsN5XjwpuEfHCaOKor/hluKjYpbhDWw02r0RL
WbJLJOGXJ4/b+/oHKR5O/n8U1v0/B3Im+NvJOdy+B10LTfn0EP/7fueloQ9mm6HfQMX7pBYbq4Jw
OBiC0qD0fJcR0ucap/ght8Sg0E599wpWE/Za8KOjNS2I0vzgv2c66PlpPFV6g+zMslHHeu71OZIM
HMiG6txpH55mXlNXe2gYQR76HoRLJ6BDR26gvYMwJCrdQq7wnP9h9W82GEFykCu3bav+59onCr/W
KWM7MqmKlIkoI27SIr4L3Ds1/9EZxbSdh6GDS/3K4s4rMvf4o8m7ndAPMzHKmYndVwmEqbWDAVce
w4GGRpxDRT4vHU1hO3UjZRNFcCNIT65IEA1Tiigwlo3f4Nx5Z5IRapx2AczvKWQFsKyNKaYSvt0X
Rr4kRsM0kvIoVeYt82eUx5vbcOuA8gIWiLRqZL/zPfmHFyPVGDGwhMmIiFg/NILqy655TymqTv5L
RdhK1xy/ATTVRPYl7pawSi2qiG8bj7Aux5s9gJb+QCiJXdu+rJUXw2oNqHBEUQSHER9Ukj5FUgoY
mv5q/K1CCJ079G6WAhawI/SmpZm12ijP4deah37qIOc6sAxobxnDKYuaor1XyRRvUdQch8j+YOmK
uXO+BddS6mT4aoWUjGrtL4rES2t8OS7zPBVPncIMZDq6DLyQGm6BKm+2kGYT3RfgRPzU1T/Ct66C
gSVzLut0SOrRZVFV/IuYucOMavcRV+PaCh5+h1KlV7xTs2t2BIfVdTzcrO1NFto4alLibScWW1x8
fk86u0x0lZFYVSYQ3LQb/nb1qhdXC++kS0VsRFpmbXYxtDST9irN5pRlwXUbqjZ+W63IE4qgTMZ1
VnrHBrCq9lXweoS0mHeg2wpWf9gVtWIyo4spg7148+K+VyksaBFnWz03EhBb+2XsRWtpdrnYtgBl
4iQeKo2BElyZXA01zoGY6CnSzZAylZQ/YjFA0XHiEuAfTV+36vhzxZgHdrDovQZsihICP88Ajbed
PGOHmPP7IjHpenFrsWQ4NG0lL8lFaNJhlsABA2gAUXZx0BNdH8WaetkWd8211tTyxrOoAIYUo3xQ
k29C5ERFclZt4N/9CDlGur8xKX7Th0Pzu8If4VeMoHLKpKAQbJX5UNod7wyUZHwBucOyfycc4RxC
KWX3ru1ug/51c3V2n5zZwK49j7/OTR/tKhy0i5eXIJfzw2kcquMtCv9aUC/prwYeV5IUd3qx8dsH
dDQaTxQj7Wqj+AkbCxHUspktmppyn3kMgOyChWN+bM3ab5c1k7910vSD2Y+Z131/5ARTqzXSPPa1
MWXWAXtRl9soh/dOf828y4rXkZwFpSQNg6Qw74UE8sPsMhDa/H+eAqo5OEjtn3TvxRpVQa4T+0Yp
d+MiqbF7E/p0YkBpAhdcKSVjFO4GTHZRPGr6P2BTpbPW1tbNY7jPBWCtbtCsf1F2ZyIACIodQDKe
96eORVuQ9QhW/rWrL8SncHiSxlGouSlSvlGe901ekMSkMNhduHn8QuaqBAAofEYWqObWyuIu4BMW
imOAUok+So5jfQECqfAhNv7+Al9+551BWMqHuv4ffnXAXen3smsCmLjr22TKWMkQFUi9zQdPak8n
6/qbAVy8cLMPY0eNC/opp14RlYOuh6ZKgDNYVzr6D+HMYyGN1y6DDCAo4LQ8zO2PXXRTXBCaKUOt
hj4c9dyKN72UC+Enn/oR7O9V7W4wt03Q8dZgUpm2EBZlVcfx5c6GAsIQTNtIT+ubNaCZBsEs8+7+
TyW9XrWBsXaV8RRsRs3oHDjrl47qdV9ez4LcJd0oN4yOn9HKnW8F5F8vaJyY9HlM258HNL9WPk0p
zzHW91ozfeLgm2Rnn5BvMACArXBWuAujDBtTvBPTG98CSAoqm7uPL1kE0j2skV96j49jkTP0TO46
WfeV5ogLq5L98Ncw63BPeVl9eCihDYadiKF+SNm9CpnQy1CqNcidMYvP0DGez9Ap/7NHs3gYMVM/
nmceGo+GLyW+dSaCqeQvvEhiROGbP3pgRlV0SNQ6VHJ14w5zWGSN9vqVTHsX4jSd61DI6Z8BG1wD
23K8uF1ZBRlXtx167nVVfqDeqH91WwWlaTbTjLeq/yqbRs03hKFvq6LCVMqn95fTN1i/C6hV/rEQ
JXhnJ9+r+apcgcX0dLiuEGADxrFJ3xyarW2u6NlpvkoDX+jICysIv9OJsftYCk25PdOqhHOvSxLz
CuhScLA5y1X/lWMy5yMbNOp9zc2DroapFNlJVxuZkhwtynzyiOw+8qxXbtu4WZONSBvxqvG2Y1Kx
UZ3O4S6QW2MN2w91D+3J+aYKyHV+qUU7KBozGM2DMpiW1ZIZbvw6qJrGlnKe5G+rGdeIZVZcjG7B
TXypKbZus6yOtRWrZ6GdyT5gRX/+XrSIzaNNhsb16LRJq/zDtgDAK7y3PSy1DoJFLYgVAhu3ig7Y
hLdGtqpbCneblZvH19KbVpiNyrMbmfCrVYG5igefsJEVKyEre4xGVwDK697zqHbi7vrZkrmHUNOY
hsKwa5zacxhRfNvaqsL4/3fBBhG9wuaGR8jwnO3+xlI5qkBUy3Wr5MLo4zdDQKegYAq0WXprHMnD
+r2HZ63i+2Z0WKvcDfkdZXlIO20OHUNABfHXjXbnJHzecyMLJ7FGgN0JI83CRb7mHIFwyR9KVPvF
XKXJvbhp+s8yBghaWna2ncavFbZnXvdM0T377Lc4i2yR6OgGOco5tOAxOLnBMxu/dYrRU/NtqEQO
Msx6tm4xjzy11rjgfe5GRv97tHfQ8s+c+OfMdXxGBbWT+Nv8q3GGVfqREc7Ch0GtBpEUqWts0U+M
+F0qx197S/c9nMFcAyvrY/ZzPiMsnISfa62aZ/2xtAW7gxPUBsnL3uACzkr8dgoFTbO4oeojYKn2
/RNLbZvQdNSmusOVNuz/b8gecemV56wFDZ8d4k64yWg4thS6SsCvZ06tenmyUjBSoHsbyWFr0vcc
mqtGhIJhW5UyZDkTlP9IvhKV90XM+C4v/dYQ6/KkSzsX2y9BGiq5/1w2Ry4a188YlmrqB5BrjLar
Ex3uENiZMenpmquEzM9QeE7Sf65ibv5x+NGDjFWB0MwIDM+sA3gJt7n8SufNFGyaMFahaf4w1IfV
Tv0GXWSDxQW6VWk2yLhqUNtI5+oZ5mvXb7o8q5sUfVL9XhCkDTO6yL0Bor0rT8xPD/6BJKB3UEW1
jF9EV7FDv/YoBx8ib6uKFV/9KN5LZSICnODm0xjrvKOGPVOk9GPhwZHQ0ByXzJf1CMMM7vb38lh0
ekt+npBVscRY45GlWqm3rUPQ+ryi8n2xOOJmjzpdmnHck0wRIOx2Hd78lq56KavamlL/x5YSRRuI
iME1t6hW7dmDA3YI0shSrNHce9GpjR7AN7++WIMBhjPYfcDqlscH8OpNAGsIGET2W2/ANrw0JEFJ
F65E6abu5wgm+A6OBoEKBzvy8MuOUe0gEWI0ypcYhz/1asHjuw09B0y0D2uP4a7ebyTEIZBiLaIM
Ocpq8YAFd/+bhdQDlSWbG2gJ+gjYkajdusPNFwxcfADI4a7PQcs+lVeBSEEnlhjR8FdvUNuMAcFy
T4Xlri3jBZ+A83AfkQH4wX6ab6vEwk1bTeDpfxPhPo8HiTA57+9VCSTFmUUBt7vw0GmTLUpLElK2
efVlLuofXC/nqBYeQXv9zYI6stPFMDi8Mlu3BgDVtG3tyyMupbbZQg+0qv3vtx4Zdr45QACvdZWD
hJE+eWIpudd9OWiLJlDLX91xDo6aStWTUFF4N5vd+U2X0n8TB3TdlQFCgwitFc2zPKtjompkvnYt
fqiBlDMPiSSqTovi9OeLWGuUpxdljleZFI6gGRvBA3ZeQQFHPGxUieTpt8WsSqZA4aMWbFpcsvo/
zmjA/VMOjXgrgt5VMTIAmZYtckqC3IlLw7mb79gtfuXtEgaX3JjaXw2XNdGeuUtvxFOR554gpMKk
S8q9fB08JWLzicKm25CpVjBPMZT3LxinM2EZEvmb/BNHYNd+tFMUCghUvanOdcEw2MM0U0QSB/5Z
YLfQwurUhKgc09etfILEiGJkSWUOgMG7HpVBl59nsM9e8aF1/cv7c2CyqdqLQvMwr5/ceMBPlzcN
xJqGba8vzc4rOh8SwwYqtFrerieZkFs4KM6LROE/AUOpg1A7gSroNCj1ekFw1jft8yXkPx28M4QT
Z8S97YYI4jaowlt6MiRPNAN/nVYIHugFou4f3I4jj0xD/bsCS1vmEcZhbPk6F5LOZh781HfQs9WY
+nGYXPfq7NhYOnHuz4RnNKu/Dsi5CotvGZ7Ang4Od2e56VFPeA+VDXcI908zRTWYWiaEUZiFqIX5
/gyp2M+5IxU9ySPXdAt3uNK0LNDHPhiiGCe9/dGDEB1ReXqoj7RZq7tbpM9abders4npYKyPpEKB
1VRpJ03Hj1Qpekbxkof+ByijmDS3ac7y3tvWNSqdHdWVqs1s/JgThfscUomKJ9jMXsdl1p7yxPD3
4osHpgpHWFlrFDmGZ8UN16c3IjzQ6+i09r+Lk68C0fSLk2McGEk7KcMZLLvzS/wliIPVEK60Iaho
DDFEcS00pNbI7MXA9cCSovfVCmay8cCu3h2xr5jumpGnzxXzQZcJ3Vt1ZbPxOjLCRjEqRmKxZPlv
9FRi2sJwM5fU+bEwmJmihDGUpO4loH8E7gYR4HyGCDY9k+YLXB8xmmJm/2SMzJvMTkIUM/AYIiJ2
vUdwngY0PdC+oMRIly7sOEYQ7oBuV+BvuOib8SZf2nJvdUkoADZmKNqKgvb31qtaFkwTw/ZV/tSy
7gdvQwqBVXbn6Nwd4r8TVcoMpv70LKtA6oIyJYNxpfQ0jApxX5jWWlbyafKk/oS1g4MRlaYvRCgw
T1BKMwE8Z2Gv4RL+6MLvyS9fxXAde4+WuCRK4HHy5BxRsC0OKDBfQ7QmbY6hLoCNHmzL0yg0oorO
H+viy9pI75vzp01AyEX1mnus/93WABbCb+pqDU8b3qTh/EwIfYLVZWzNkMgEySuzrahI89FwnaZr
PyiSdpif/4x2wCHYrpoDLUME5YqNeXCGgLV6UVZ7saNuM0hZOBgCtpWlsN2GLAT/f8Y+L0WNEkJ2
ktKEoJLJ8kd84xnJYLIbnqpHI+5pE4CJQNqXPwKKF01UdsSsuoEFswAqiBJAYMsUE2XCmZCxAwGz
9Oeo3nHDa/UsO0aGj4+gDUgYieEVb/j+g2GAXJZRquT3yDCD1URH6cJgibjqih4FsFaIQIPGUIWB
Y8qIjc5Vjl/qxBTh9zq8DjjveUsMFTtXhhJZn3f+5jE5zQT+GptWjLlxFoekD8iZsc7BA6oVK8pO
fHX41PJIaWUFTzZly5027866b6D7qvTnr7xGUzLZr2hLnwz+mYDSRY9MUm4gPBLPEFnV3wbm9/iO
pp9o5/OhTZOwtuWz3dq0mxXNA9y/304Ntpex04h/tYbn2t7YdEhcuaRIvYVFGBgZ5OHAfCH+9QRh
47KYVlUu8V/j2C4Gr7WzDinLBTynQnbWP0UYJcJJJEgvYqn7ObZCmk7u0kldKlhXWXgsVra0ecqP
lYDo6pLkoExDUNO1lHVfrriBoo4/si1PT2OtNTszQ0l0dEN2+SUqkkrJ0X8gfx1bj2/qi3KllRm+
UZY2wFkEJwYW4A01N1f7/XTrESK/wvcb5ZlblhQyOlt7LqJvYqtUFdIqx5N45K2tnSdMZd9siqRV
L2u1wiEYBx1gC+UVEQQB2k9UWv7eSIw/IObP15GNvY7hM8f1jZbfiFPBwIh3mijFe2qQFcdtOo+i
iRrjxbj9YkqGi6QLMFhkFAUdoxzBZnvYZiytGopCmEZpYhMlzK2I/tz7OmTMdBXWskB2jz/SX4kj
PmIsF1xhl3KY8i7+8xdj15p34Unxdux+rAmW0GmidyjvP7SMmHILhV8ds0cBorxhPai/lm9Q/jlr
zuZfZ8cWPfT7Nwnnt2QZqjb5ies4ig8XjUXYhou/b5EAUv3IDgMaS85QuECpv9SGnnRp2xdE3nzy
QG62R3hbziV4FJlFNdFtnVCiyVpVg1q33pB77Dmn0cxmomb4LpDMd4nYAQA6Qnh0PlN4maXP+Pzh
mEmxwbjkO8nAK5/GLT3T8BM27NmHxLPOINvHdf8CslYNnR1eECNJ5cHepjbojttPBoXrfi9JRPNn
gBOORzXVGjG2JQKDdpWEkvf6c6B8J8yHd42/Zcbl9raV03C9xUvb0ELLr0CBlhdUIPLegxcLNmfG
6AX/pIRVmK1kJe2dQoT/O1Cj/EnAisBS7ufPvcYLLscCMAXst1RGZzAVzPAyX+UueDTvCbpXJfjO
yZrcoyEljD1kBzFncuG7tmgmqX0xvfEqpwD2r6B8mSERDfYYuIEwb2d4G56xFdIso+yARyb9ESsy
J3+dlJcN35INXMrAYtpQQ4qpzp+oDNpuFY9F0IlLZlRMdVwvXkDAouOlqND9F954MBLtPLG9LORr
OxcG0FOzcWgYZhpR0h/W1DK5zly5dQ94zsJ7cGHrYE5DJ3r/aPbnE08c/W7kqVYdX9A1NYEl1pJV
HJysmEc1u7cLJkbYttYbfb1kgm9VRmDg2QiKeoQ65AHGz8si4HCkVXZd/Y8TQpV15CbYRXLDz7QK
pdNbPHJNyWgyET/4QdkAXYbxwl4jCE4Q2/8X/TOa8aPW0Lqr65zuMrudRJcnL9dyxxqsxxXwbESw
gliU6L0S3PpytP8ygMrYqOZq0wvsY1U2FsNle7rEu3avHZsunKNH2j3hZCBUp4k8te4/1aZg6nh/
3ZoQ1ZpDu2C77i3mrjhyyrXj4oEdI75Xo/TsD19AEudaNQnjuP0g3AvuX+MBzWcNFtD2de/jvFfv
YVUY+DbLUABGaQN8xRy9uGI840KiwEfBvZ6QBjVUvPzXG6zWZzW2j0dXznuWsmdc57jp4+oci6pN
6G+KbgMX/00es4cXQfR+VNb9zSculFDEV2/L28IcNukR79PsT/p1kb6VltxvM59Rf5LD495VZObw
ingbNvv4rZIuVcF0Aj0gkfQ3q5Z0ZkXEaEbuTXlJuUWONMetF2tqOFcb12Ki0Lg52dPsJGfGSHF9
7Lh02t67T7RkFoAbHyOljMMIZmiuzHfZTouyVsuqznrBn/gTdMPosbMBSj6YtlbL51mdSl/1wVIg
W5fXtvyf3/Q6Xl+9Z5linS7Fiv1/PLUU+G1YEQCM4l5WfEGIpjtCwH7ultKjGM/7tC4yM51yfDnd
JX1mlwhPtug2NpDgg5a7iLKHKLENMRz+oswPZJXDexuGF5ljBw9SKolHl8EQdk9fBYoQXwrReUgI
ATimeuECd4sp037e2qlNJS4iA7KmvIvB9Aj2P4/DbOw+hJ3D2YtOuHg4KFAajZd8imZqVM23CZfi
++fPfi4DGV0YYPXOQ1/HgDY3Z3jEbgV80ekpshyZXhionjMGdu4gEmL2rIAL4KVpGFBz6bBEK1A1
hycDSpr6dbhKO7utH9nivwClWUZHoR3H5T9ZiryAQZWnHdrsNUU4HhUdGlNRYePK61dB4P2d8KN9
RWaVqNaO7RF1oVPLIyDDeFj+PvpFZs5HyjPSwMPJYf8r9leqPyu+a59KGUEK2b0cZIICfrHvvS0s
jAKEmhMlGXb+JvcTjTv6C7HsDMAK+EfPNH4ew7H9vbp2D5A60ycUkrNqZYLmNs2rGAlFFhuqS+rb
77HqBcfPI/Mv57AHSWom4R++o9orwdLQdUe4io24DaP0HU1IesuuFfJXiOc5QIZ9IXcD3U2h0PaI
qxOhFCzFwSpum8werK69t4NRL9xITgWg97+MlA7Iqptn5JuDvv3tYs6Lfq1DYEW0VsV/ePhyv1fI
50v4CqWjyHhNDtTja1qIJoaTz5MgDJSelata0eRciDz8NMf4du5Ir439JADskQ6id/2O7KyFVnHv
ZRZMNnZsb0V4H91qKrYog5vwXFRu/yWUV6NLhdK77HKyfbpKb87PlNMjWzK83PBXfxFMiw1BfIAX
+SwVMDEOVeVQpgRMIv27K3Zcb0q5N0cJ01V2NIHbQA4JID98S1cVBV9h5EabkQojL/hi33GCilFE
jAmJv4qZcdu9tKkyi5DmtOxLmG/VCbqknhduUmQ8YfBOrhs4UUASgBAGoedRWXpklyhJ3kVwpAvz
dZiueLKogjPEw5bwOKjg7q0D/6bSJlXsNcT6cesVL07Be2j1jTlIOJiZRz2ueJItMc0ndH/JjV6s
Wlhiw8sCXO8k7UGeS1z1n/48Sj/r++WXhINE5+aKCasscYQxpl/4DB7nBuTzFRcEj46WZkRUWMWY
Lc8TbHN8lmJgY0aBcY2YShLcX56v4oWRT6jytnuriEQDXX7p4fylLXX32Z2qhapaLQdyI5US2uhj
x7PapszNcdaXCZa+zK7R/R8D8BPv2lRBBQEfHwGbeTvfOp/VoDdhtLP1jGjrAICKom1Om7ywe/W9
lMNYq7nlAxhli/jEmk/59BMSla/M0xJWP6X1X9LNu2ahWcnUYhbPkgdWzccZ5xC9WdybO2/K9qlI
50PzzlKsuPpAXoMUtUZlcIgTl4WWNWi6HhA+y0CxEeGvJ07fjRJ7hLTBkYQgN8TrIInguWDQrVJf
FTLteY8U8E+Kj2O5YjXO7xoerr4eNGg+nSvEVGba1/W1VOVV+JkisM7+HLZkKNmgR5wNIim6RzUT
lCxWinJoUB8OCyaohFMG4wHxb76V7mTpZvKA5AbC3xemNe0LdF86McglmIb6nWcMlxPXufcH0dSu
6czuJ42nuID1MGRdkbpsoRZl89dLKA+/yIZo2eTOoGrCFIY613JSrApIAtQtG5KLmdSHOhtZ1Z5z
tezg84/CxEnfloE5aJUdv74kHZTQdCvNqoO2jI40FaFSlPNEHVKVeP42yqDxB3rITYo/7HsSz7T3
CwEYtKrI1oPj8x/MolIOjFlADl30g3UNK7T1UkihlI/QJrJPyZqwUsi9EDIPc6QZR7sZv5tk9mzW
5rTvD+5FxOP4sPuJ5tHMY9fMjBmd7xWbNfK2fVUe+IuLFUhYFgEalpIcOTBsxP9megGxpuc1zWlW
oQhWWYG5gRYnPrB0KilWBZdfxy/QUpJOu+ZathSUyR4Nten0AQmNcyEu8hEfM7LafFvB25TE9sm9
s7s2x6zkq3MKvgOeMmkUXd68BwvXKTsrgldjq5VbJiQAAGHivvlArLGemh+cYTiDMdU4kxnKMWuS
/pi68m/Gj3HL0E1iv9/0fE6PDzyfGReA2SNLD+Q7p9BlYrTlvmgpI0JbcDZhYxNUoyDGPu94bCih
Jtp0jeTnuZ5R4+W7+7tsMAJw07N6KQ+av8hcYbvhTqRnjXPgwogdT6p4YTLesA2hV9BsJOrUEpil
vKFIFidhI+9KlG/mwW5Gtw4vh/m4QBUEqbv+HZq52TYI1zGXSFMERPCBOQAuHaAoCVURyLojKkWS
Ffz3PTJfUIAE0I09NNX4tVPJNZNbKR83ANAcArA/hasfAZhtdEUj2kHakFz++eUi845pdU2JPYJJ
WcR4YD2J9TZIcsg512INydf9gpvBcW/KLuDCAQ9CZNvh5aDkTNJcjntpGSPrcBfoReRB2t0A3et9
Poi9QTrqFe6EgFBQGLh2Dkzl+c3eMddcpihVG5n5/CPCl7en0qPpkaeYgHR8llAnlKtFDZHTmwT0
KTHavravnE9H0SNgYt/eqJNwAtWU2UtQ1uCltUxb3qNgk8RkiXAya/g1EzaFobLMhWutmdKV/8y9
lYgO8WxQNbynS8uK7MF/SJG5OOHKC3D+VpVPs392BdW0aRE/yDStAiPiaLfmgdh+fHS6Ju2ud3y0
KMskMJ9Tqsh+oQrL4Nm36bMw++igSD+1IRrIonm8WRYNPSVhg6/UQrdvDsdYFJV3ifhb8PXg912K
utCD85unXUIyakfXkENRla9oujsj+i9JMebke6fRUdMvMIXuDPT3kx4ae1OA3O6Zwo7MI/whQDyW
NEPIttM23pQ3cNVTlgLHWn06fY7jyPCAlP+PBJTUchmiV6c0pz2BASNk0vzK5OIRSLuqjpn4iNrG
U7zWuOiSlDJXKv6oqZ3mkG08YVAqeeY3sv0NGA9zAOzRJgtr3GVCooE8s6jQMPxpXGXuy8ocMpN6
yu8qTwuqSgdNRBn5NKfOZV3xj8rut19yC/TSd9LvDiuWA9I7dKLRUAChT38u7VrWa0nH1bgtX7+L
PYczRXWECCarQBYt5FvQP0d3IazvpdtEr9t7fpfF6ricnOhS9HdcbrW5Ry2RclKEy5PFTR6y96bc
jDRndKUGDy2aVs65TmRpmuDEYCG0cSFSn6JUfZWdOmnkAsHnaJY3pBwCZWyBHF0gqcT5OmucZjJS
1NIInsRLhcT11oKSlPRjd5sh534jX89MX7giI2nBRg3YcvFAHSZLrt/9WMbHH4BOzeQ/adi+ec/u
1gbHRlC/vDlECWFzOwiXryHWoXsJHx4vXsAEhuic7JALHwSepPlUujEv908VC5v62oYya9nrRjfH
GsyD2ssR/i9WN+1F7Z7cvQVsuP3oPhZOiqVyrE3QqRtIQ3EXqhd3wxurzkwqTp+uqblnRepeJELs
zsjCo8E5P1pdZ44x5yM3OLvXL91Bv0bWiXHC1BLArUB0ZD1zKVK+yibP0+jUHrhvcTLrFZDvJiHa
aBDXdFUzMzr/uemGfAJm7+HIPXOTTz22B/mbrP2oavMmuWY+Q765oXhqACkcwJH1wGTyxg1InEJq
lFOd5PUCRRzkm3+FDOMHkVdA6EBYh4HRDb0YavWXWzaX0IgduvtLPDevG/i7Aoh2Jz7KpAeCPBn1
DVSBZBHFCrhnG22122ChUAuTbepooJoTf0vM6lgis0qiEmC0mT6255BWy4/U7i2thEnJCl/2klA/
GMCj95PAYP3voyBXG8lRnJzODbj+jWchWCHmjn4lGJd8nDpW0eXcm6sMWIdB8L4IdXaWfGEreTUK
NmcXC6TCuJiUGNyJypkmWTm54/yL+LSOjMdpLqHkJLq/oE1M1UIvCSX9VnJIrAZbUH3WmHawRRij
iLEcs65sawZWV1dYtpSFuYjXR15/sDp6Ef7GcMVoerAsEvBWZvZEX+L6vblxkAj8AW18rJy66Ins
NskxNwYKVF70A2+zL8MrBcXMgr3/Y67GykGIBMHGSuRm2HZwXJeJXNuKLX7IyaA36ZWdKk5x8OQY
G/2/Lih/KhRrt6D395bKmoP879KfuwgJE7iK7h3bk4tMXv1qJFcPW+tGRtr2KAGd9MRK/gNhQ3vL
A+OH/pv5iRV15oEr93kbwISGSA8L+ZNYS7PCrMAUSlghcYxyJnfKERgWAKpY2G4khHOLFEuSdogT
ImmC2c/sRMtaJ6/YPoPPBHeHe5bcpqITKZ+5IEqoOg1iFkarTZqliiQxeRgOgjYx8UkIsbiUNTAr
3//Ic21FNToRCQJ9U1VzCffJGtlh+wcWt82aGxDK3VhlbtSi7GQM0OHEFbrQ6HZtqufUQ5F3ojy1
odB2oTdhc8nEVKgOE9keMB9Rpf/Q50ZN4x9IH350KCKBV78AwcSXogDLJpRAcMPReSMKiUDlu6sh
HfYe52881bPyss05CTOj3FqWj2/wjMICCM5tM1TrxD2ftQKGWXXtAiv8v5+3s9fBpII9m6HX1qGJ
++T+9fTxN8b1wwe97D0S8nAT38tZLgStOKVk6bTY98oxZG7jlRBviAwqN1B4PGx3uOozTA0JvKgb
yXElj5iNjLhwv3qWeN2vGUNVLEixGH7NhJkeue+TSQjWirgICJPcCsaSTffeE1ri873/iCZ9DAlP
6NRIjS+/MZ9ToimQO5PzlSTQCUs7izvLnFkUQt3vR5cY3TeUvezgQ5IxcQ3tnODaVl6rvJZraIAd
ablJa53S5n5RsvOIeUauM1FhEZnvY0AgZ8l7EONJBXZUfu7+LpS3X5fWCqlpWbqcq+o0VeHdoVgU
x3jfRWX+QsAEHFzvb1azeMQZ8wMl3j1vH6SIC9itH5qDFhrVzu3H7yseUVhbZGQ+kICojzxmSF4A
CPquhH3RLQUhXQoGaxNKNYrnrMmJIHTqzLvvQViy+1QVTM0xPMOvSKRhTnm/Bh/Q3BcmgWl93Cxz
kPsU9YBx9g5149oXk6usUL1psFH/Q3bj7VZId25012hqZxRJ8NfrsscvLz4sEqHb5X5vpBb7a24g
jvaBlI2TL8OeQEjBKtM3bYeSyNXE5RKyUOAAvFIyh5Rt1QGEClmpRRfeM3ocEphDAagR0xb8O0QR
yVsDQFNqBqYbgHWc1v0gQQrOSIUkAAVpOD2dZFvPLhrmdEk5LJiND4jFF/onA7NOoWJKzw0TryJA
br1sIGAh8cDaqRcmCuw7XeAz3tXGATwFZxd8N2E8dyVcgnpFIw/lrpoRH1UV4cJZW7JgrjBHBn0G
jqBgUnQ3O2n6txP3bbChcEuryVJmZP3gGZa630xhHNnKQtG1Kz/Te9i+GjeijD1+ZEhcuwv+JNr8
/lMcqxvV8DnE+UiVUIf/1MVIX5AXpUGV8wMEzlDe6pGfTQhnLA3gO8BnAs4YWOXJSwqe8OlatV3D
Nc7ts9k+kfEpWFCSukKOgx1TW1MeoIMIwFzBE7q+EsIuuE8e2/T/0C++Ah0ObCD8nPb2qzJ0vWqf
d7WHEJ1kGNVCIPSa6esHp7OfMHpsRMZw554gScYxz1YKl4uMaLhIvrM4q2vPCFFzyy6wdoTF00j9
nV/up/9QivSft59MLCZdD8wX0SH+fwyHe8Z1gkEsKMU+r8nFsUOUAmAk7vZSjb8g/qiR6zyCVxaR
vXf9ixOgmlUiA1htHD90TRqxqSLblZVteAgmgFKkhiJ77cKkIBL9y9JG6zKghJ7wWWKYBoBzSCoK
l2yNnj5XWsCWj2tYbaH8azHysOuYLbcTkKCYBRV8ljhkbJJprGpgpr7/XbE+oAKRy5D8ewslITNv
xAyyUP3H1kebiUv9tXMq2eUMlgteG5adDyupSYZxNbrsA+pvlJyp6S8h2uMobSyB7vCxJAO/Xpid
rmpLi8c1C/0NnAp32Mgf+QmwMQT1MuQauLaYdsQwFTcQO14X8Zv6kPCMvqAgIjlAOnS2aee68DJv
oq3z6Cpp/b52cwi8SUKLl24xJIij9NTL52DPPVByT/NMIBO78U0azaJ0LMFeYRqUUPxgWXVWWOwz
Mk9H+ZOxw/fnSpkwcz7wdq93nm9e95S612uHe+O/emdysTxjRC2ZCeAeDGunzFq+o7irreU0uYA5
umvbXCJOTRzyLHhQs/9fraEQfzfjQCCI3W10BRaikU5D7CGcpmqq6hE0xuF6a6wbWcF5LH+qVaDl
A6JAITaQ7qln0tqeOgUuHAYmqggvNigitkmjeorMOQi44GJbKjaOsNmrYBPqWETfk75gkA5gmBYa
qHZOMtpL19y4w5nDMOrHfjFC5aqk3O/W2vifKVmYapHvU8INxHcRNWXD/UaDi+Mr+TFSKeT9ZKjM
htIkB4BFENQEGywLGk/R6vmO98VoWdvgGxFN6fCVjL1NYTBxRwTh5hkb6RLDWEW8KZDNHYQruBVi
Z147MXTIx6YanrvtP/lgENWTqSFJeiUz8QyQDKM/DdQdngYDiFZAN/y4k0sj/eOpWDOZJ7emlrqr
dNTXQf/0RwBoxntwzQi1uySsPdk16MbilvB73PSn57LvjTp6CfmECzxu/RY2SZbRyxN9d8Uc+f0y
/CSCcLqCsyIpupq/cvmxj8nOlue4VoMate3QR9ajgE5CH0oCijZxInJbeuUGO42tfQ1Vrx6F4I6r
xZIHoYIbUvyVoRz4Da73+y2r31Q2RxsI4giRlyR39gpo4KNloR542R7BDhcyTYzkRnQzW/ZibR8O
uXleRs+JkWluC4BViMKbTjayiPWzZlvvKEtAM+IgD0ZC77n26hIWIXudrxtJxY15d+geK+tcGB50
j40n7dUNY4Q0wXCJYyrFWqYPKUcuSYoKEih3o9bz8tUu1hTSPBw8AV4TBT6KlvpjpJcl2e+UsZge
xK70WxTLnVzWRj5Y5CtJMFqYP6Entd5794A15to0g6tk8ASn7KArGTMvcIRxsVpRzLuj25Tjjc85
pqfPpeTBKT2aOggk0t4abrIIXW5jQeL0TgYNHfE5v18K8e38w6LvUSHbtztlFj8G25Elv/Ldr5+/
CGHO2151QCF+NpWiYNvKUG1Aby7AHSyc6RVP/Rz6xotODx/KS0gQixSE2ysKemt7HwgMNK8PArmX
snd263n4c0zoK3YqMM/KBDopMCNlEaaqrgPqVoA+lmV89xwV9nFBTFJF/hzX99OaiU0dnydiP9ZK
dCM5PikGKOp1MYaWT0QGQHxHFly3iYv8TeBHQRQg5JdJh7mrmGmZIswF14xQdvmRIN5GeAr1XF3F
DWJsBS136MYCuCjvyv5uNgN0d7pjo1w4s2mp4fjCQT/HtB/RnnL5c+JZ13AyTm5w58EMBWvgtQ9s
nAfIOToYX2P3Sc8N1Ytn3+4Og4274sDwvOScavnauqUc+HkVXiOsV3FNiH+p8+SYVfgd0L8RsLuR
nkAf9QQwisiylnayMUE7anC6MDNqngatQK2p+J3wKUUP2AGDWsSdr6uDRaf54rANud5/5kXbX/pa
ssj06tr8foJKBXBFkgCMNzz1+Cf5YRTgQO4njoaf7dJoDLHG98Iz6yzVuLRz7KjtBU5je6ukwaSt
B9i1ZHDs4wHXascyp2LxF0nTDOKtZ9JFnwTR9kzrhXZ0ekKi3o315MobGdtWeE7+liLetrpdu4z4
CoSdgGuPMcMR8OG0bkyM6fny7x8cvPtdXMLLycoK2SJvxxZixSn/WK3WziVs+5VG7tj+Cs23HrV8
rmkEVVDgpXhlNBQiMhO3txsuMP1Rz0Mu/d/5GaXA56S33KqW6ho6vkZe62UGrbGSwBLbfu71GyMS
LwmgXR5p2qLX7bslipQP/E33pVffcObFTqMBI3tFOzUOXenTr46qnqa+ke7tbRcm77oOzjy0DhPl
wwbC30s5cf2YCAX6NwoIvuEi8K+uBH9jcLrgb6Mhk0dXClZ5W+nhbNG3aZxZQiiobFNua3V48Swa
5w8jZs2ZpSuctOF4JMoxp+Sa1ZreSgKTDReOtbpf/eAjaj23Llx548bcl3aScK644qgjrhL7JKAz
7bdBzXDIE1pGfZG0arNnI6g+Bd7/LBwd2Zxl4hNrV5M7PByKFKwKt7YXmb9Lhz/BVdxHHFzNdbfI
L83XPuO1lWFnOuFLCX+uS7hoEREOM0GfpVLoSoYv88sbLDVKqmzzO5QA35GF5AaPfyTTpQ5DSBxm
KbrXLGGavRm0sGrpnh99j7EmDeLXkGxtY6IKQWOpo0xhxPLabLrfp3EE01u5XK+/UUQ1aGFlp7Zr
ktacSQRcrR2U5Xwv1porBpxoK2GcBlXMlMeBUly2jc+30QJJNb+ff0aIvq6krtyitTbnm58lErRx
0SaV2EejOrhcv7cPu1G2Hdrmcv9thOODQMTYeBckHeZXrNEA8jB/zmb5+yqWM9RaB2x6xb9C+kMb
BdgpdNZYuZqBSdHUB3jkm8gxlsE5oD/quGEYUobu6dGwB9AJOhaMBMijG2xW0jOqsJd/7wsmk6LR
sdSo+zLWZMn+cO7t/wv4OBBF1j4W/Wcx0Q6Wk4bPQSRSnR+HJFPZCtFD0DO52eeGvMi7J4ESfqDD
w1gUK6tF7DgWLsAnjR0XrrBTdqdyUg0ODtNgIrergTztQoJnvsLV2sUFZxHct8vLqDZVckUc3Crc
pqUTDr/r9NkpoZNCg7P86nBm99be35rFgaJI+GXzd2sXoD2h10EE+rAWTYvE1pL7OpJzlhl4c6D3
S1/1ohF7VgPKMz9CLRVtk4GNJxz5z/6DhnkzUvzeMaB0vwp2iprQ7vD6WdjuiAvd/eN5DO0JvE7Z
XvoZAnWmaTO2hMlwzFwjNRCr+He+/uEwPVmNX+YErgkovYLdgSwloSIk2PXg8NrDBQqqPDxA1+Ns
pNRCtepUw8CSXuXHicMDC3hpB0fJY+bsyMS6V+GLlBHW5Gbbm9MLvKmj23jHqErojUjVc9j7eLiH
yX0r25ChW7+YaqXCIgTbhYwkrV76f3GyfTTK5CNUwTEDXSJLQHYKn6+ke5Sxb6LONSndDuQPnsGX
FX77E7AcO90s1HFy3vfmJIJ17S4GhX4BtgwvqGtKlZUJNzHVOgkWJ2moZT39wF+TT5S67sOzoCJ5
hiUFafkBwYyUHn74SyA3LmsyaHSGnzXiL9BXUc1X57nLHnD6AzV964HGI09i23DQaOHGpX7uoIFI
EIczDqOe7DPUsIjZXFs6jjyPyM7RGFQZotu+3mbQPWW6Oig8VAsbTmwbJOG9CjuTOdUJCyYEtGxk
Je9bp27tGOBoRrF/1GkJw13s1qkEWPYz3N6H+/0G6/SmHizPmj9aITyuxBrn96luRvORxAYzVtVb
yzIp4/eXaxuqxvNKk5lgZgqBbk54/p1G0D61PWWKGsjylnaJ4NWak1B+reS9WYilzdDa/QbUdrYj
fSuBzhNkn/HjOggHMpATZbfVu8xpyBJDAZfM8ovtCydBeWDUUlhRrCX0IQxd4SssSsCHW0as2B7s
LNfDIFlSgf15yDDQwEOb5eocRJav4UX9hQpIYZspGdRBYlzwj8OZt8pb1V0QhqLCpKHRDcZj9H5b
RufBYG82p2fdPme2zP+epTk3GVhcYIvzQuSgS1qsoFLiULQREU9gB2Sig7/ibO9ELK4VsOxQNFrE
sL6AkyYRQ951AzXfJfrbFswQfYHUJpub9fROBZpt1DJytQm3ZYuaLGnsY08gqboIXS0/Fn55s7Dh
PAFkcDYR09vhVKaGsSWTSUlEnq49HLg6wtAwrrivFtVe9cTfgIn3PYTNDdHNQZ6zdRYmFg0Xnh6h
g1C8AoXxBuaOQvoDslBdycpHkgbK26CqCEs+MKlucmhIPvGoiI4RLFkLAozdpdXqF36BLItAvGXj
gtLyeRQQyhjJcxS1YmaRqLX7hLdBNVSYo2Z6JOnQt6GXG8H6EyK1ZZr02hSf0JAFFFns//tz0DTi
ANGymDg2LejATYbn87UGvLOUWCFlo00bA9VYVfh3QwuRGAxFKqdO1eeTqexouzJsbuwbqCc/0HDG
9tgZ7oNgu+MYg4ZBd2Vzk0qLD07hYWqMe1p3mO3zZJFU9VN9/tS6amTHI9SNb62PgRi6eJMW7Hvv
FglF+cPtS9ggQv6adIXz11gmsFhSVn/GbR27oHxGnBCDkQTO+xU6FOZTzAkPh6F30I5bnGJT1v5M
5Hf/2QVlutOb0+/GnoZJdN5AN4quMB30XcXchQRPzNAzxMxtXjz69PVJMGkQRZHHd90JTUWHBbF5
SRuuRViw9AL09nfhdnqegFd2QLGxXZ2I8GWMQ9el4BdHABaly4aE9XIdApQNGrqKLkcuc92pL0M6
ZIL67ubJ6mpczF9z/bP+q16Cjlm5m9tHR2myYX/QeSIWbNzcIUhUgxgonhQucKek0fHYqsiy1vxc
17cfkMawxWu5CmpxvQuvvK4k9EuV5r9J5lQPMMfUQZgzmgcXTeXdyWyqDyBApDR6R3wSG3HBYYNS
J19Ii4cqjBTtO0MdI6QWggMokGs+68UI5FPgeVSgQCzJvMym5HsY4sasn7Xh40zWCcGAmEYCcrmi
Mtka6dAHF+gmU2ElZIX9onysJImFzd5E4JSjH2bcDUo+yYAB055HWO322TZRYI/ikdrg4drX2P78
YAtU9qO3Qz/2yPeXnBW4T2hF60sYxBf4+CpLg98Gn0CoLx/4P+R4yn9mN5o/LqYzEAdpDTAjP7IQ
1BslFvDu2akpfbFtEwU1qixu5uYzwbKeem+tgrGjO0qMsc685Hhb/7/2nrNqQi/N2mKG9llxJ/Ra
rntuImYdX/32a5zYgQvyLVrPiqurhETt4FqyM7uL2gJ8vW2KK5MAHtzcKCNdaOacqi/doHO4LZfl
H5OA9zy54U/jsMx64ekGYSAQdJU3txsWHBd3wKyTXp41il/7FAcKC8DuoLP10K64KfTdC+cBssjT
kzn1YugdIiSh/Pfm+GpY63MvkZjNANt5Ic6ZNMhXz3fStZEASRIPod+T2dEo8uGmyAYeQEbqDmaO
iPhnesfJeNkAJH7eG4i8l2eAAw0426EYKFg29AfbBgb+jTBa6C1/OFoV0u90tQ3qXSWbIBsTjiPX
BoCl2mefWwrtqUv6/ep3iE34eYNMPa1aWJj/kIBo6YjAwH25XWhfGIy+IKrjd806O9udgopP6CQa
NrGhJJtpaX7kOocALXrmjoTCxxqUb51UZQwRWG8au8prS65cp0BJfmMriqxgY9lC+dX1AGYHUuTL
uTIvqBLzlQZkN8e2l3TKHX8UCodtY/CyxDAR6McrwH+yNTQipSNSiimOE/Co7XwAFg5Ka/AmiOvG
QkV2BTP8opuR9yEXyJqyXHcumP9cwJYf19Vw8qFlo4aLoqhfKnR9xoAb2yiVWrZ+hvOVvI/+u1pu
aU39dCLmoBddYG7dXZRSW0oXibXB2tpD9Z1CHk7VJpC1pMYQIkEtgwdlJSd0g6S/uT1JpqlvGG/a
KI2Hjqmsc0yCfz67QTPBMejv0KvKdHDe8qcjuZQ+4KePVsw+VlHenz+WQHrrMyYHLD1TQnBtzKiu
5qO6FXAGOZUmK7vhOJ12h5jrT2vLRMRQAvlozSmL4LQYCDmqKEU9F2f7bJTFWbIqkCBPFO85aJd/
U9Y7ZCtRQ1TpUaaCMyMwbkpyJy5A9rVi0cY7WtNoiqaemuCih6ggKcuGNLjG0VwQWrWuCjQLqcyS
IV9gG03zGJLAs1wR/H9Fp0NqFFruhh0R5aI6Ag4dOGPdN2jKcelDlX/CNn7qda9zjIuiZ5yrrriv
zRYmveYlrQGwVLGPYuy+cZbxhx0r/kS3E8IxW99eR9vkh8vtePQECjtQ9Rbruv533dpWE9BWWXKU
HBLJI6AMdR3v527HxfzdE7y9n7OZcNcnoGmXyUDYGe9y3uDzXto2A3l9PMwNifD1dPYqdvaTHhdf
FAuMXckwJ8BaDqWVjI3wIv7MfRIKc0EV+YDe8npBXTU9bvAQcRkyV4UJkCXZEnN+7yNqikBgPHPn
RqfXKeA8rI/Z5gAsV2c4hu5Ax6mijDN0AsoQc3zX8lQ19geJYXz4DEUpNqih1Vy+glQBqltsoum4
9zKFiEXzMNFDJZlCLxHn9dG6nkIwr+xkmBZUDmIioiYrOzIFTKUNK2s6uNWInEhv4KyKxWU8+U8m
zKaZ1JCnweM6u2l1D9HtBwsyaBd/I0T3bEjowxaKN5MYvt7uZIIQMrmiTUR1rGtU5YSNmij0BB94
Lej0zgVDrQ2frv8qoexqF2tfZj54JmUu44a+fUD/+NITJgW//GPx5u/o3xVx2usDU6Ghb8L/geAy
jSiF8rN5R7tiw+z3/MnbUHMhSU2Z66SCQNxJIJy8ZeyO5Dja7VMPTIrOYycR6uuvHKuYReiE+eFu
VNtS9l73uj35uAnXWlxZwuWrp2RgmO8fzbl388YMYSFp8YyQmFc34MQhiCrcWX7JNI9tznVlvw3v
bngMbBUO0HA00mivdBi/qetL2tnWZSWqdvOlEroSmf5btSR0I48H4UEVaBXHPsBI1SQAFnxe+FMq
gpyVtWxODAi1j73IRiq0ItDcwu9DXnAo9OMB1UXja29fdwLcfL9Z4QGkH56oRjAXbXLoDvzlre7g
MQAwSlI0jO33yOjRiBjtz/odOuF2b0vYOdJxvd5m0t53aAAwjZ3+99F5JU3X6uRUdsSn1+1ciadm
aDR+AcdD+cLEmPJfohEsrGQUVmrUfLZtKH2QHu/4AvayWTAhaILPI7UVvKxhu1onogwP7uYC89Vy
XeXdk0tdqD/Sfq3Y19N0UNnkJxSP5cBReT5WN0TAyo0lk8BfxfyfDcZAcws6xESI1BYrjJOO7Nen
8RfUNIVzg4zaj8ncESmZ9WCWgoeW3s/SnQ9+Ql+IFVNezvb07OINhP4MpmLTwYanEVw1PKSPiDO+
Cqnx2n3kFwD9leEan4+0eAgosnW2G0/IyxkW7cGFZs7go3uqLwOuAnCut1diyYAA1zuNzzHFBq4y
Q8B01t8kAqxyQESFaed3KyzwPsMIHcshSHqluTjTfEDAl3hhhigqrgEkZ5sQQFNmZ4HXQnhZRfGD
zb5xR/vDQHSEiMuC9Pe1G0kZcqxbGVWnH9JV4qWGc7OdR41dEiqS+nrNkpcKUM4Wm561F9gYJ3LZ
D0tcIdyao/uQNM87FX/V1XEM4ovP6xxq/izk6UJHHLqHFvCc5kI64OOyR3B3dW9sd+7SjygvIwmd
00ZXUjjzbmTwCDXdpYSEiYbeWW/tEBMM84gCq2f5wsdb0ebOCB9NAvTy5YqTcYJhrp+HVY4uKPPU
A9DZHnEG24+ZnlYDwlrqb0A90/mrZCJ1ouTgeTyH0BXRNTArt23LwIINCXhuQIeXqxbuEobi9oyO
iam6XMdHhiZ+T4M7cfKgpMw8RLttLUbB3eQG9JgAEHT4r9hDoDSnUEBAzyWMmUVB1yroV6YJaI7g
oGLL5P/vZ4IsAvCgvHcVoNqJz80P1aR1SRG+AF0d7XuwgEXO009oMl5VE0hHwcovbsOViioiHrb+
tX9F7iyG12ZvdNDo0X9BQKtElhIn5gR9M0T884kvv3JM50RJBO/GXLMspbj7PVc6xSNKlxcledOn
vzbyQKKScnJI8T64fFpVw2/1FZz/VIvyiXtAtCayBMmYJhSeU9KbYd2upX95Cl/IwEZ7sw66bluo
0ZF8dip5etKNLtZOHRsrpGW48/wyTruei30iKdp1YTzLEkV3znI7bXApyofM9B08CfzhL7aTV6rL
zmxiwx5VbJ8SeaRvPxIXx8IpQdLlz9Uso+XkLX/KT108Tqs61hCgMFVgCG/OcvYzVNXRDcCsdPew
HiRUklRcvuGBw0IbUkQWRj6CM2lXu3MrFG51DPdRHgaMLhX+FwsLI2FdVE8lzCOSquTUKhcyUvzc
YAruvkzE6sDI9xnxo04qV4PUwCNfMdd6fsfPW5vFTzg9Xx5b8d1mhJ8oCEmq2ggn91KAErhPCebE
TRuSusHc8CVq2+jw4iEa/RsGEOGIOym16vUA2AnnkKXbR8G0BAgy07EicN27Um+849bVGNLvV/Q0
cRTMGIB7FpVbFpdGsM2Y+q4cXIo4vCW52wYhD7yhN/SbRzeCV8NEdTzdoXKFvve97L0Zw5DF2PN6
UdEjSHBp+4LLae2wzkETw4eADqn6diHGUngJSQNORpiWYCX1kVwpNxIlYqmQ2WS1kIOhA6Pf6Lqy
06H1mV8+LVLjX/HwddWhXTSJs0+njilo1X7SP5pLARl+3PEXl6vC3WgfwSVNT8XQyMZ79WmvPp6w
3niUH9ighRbtAeQ3hY649+fqJiG/rbjYj+RlDZgWiT8P2NGJjffq8xtZk84xiEF7dOjhRxxIdRG/
2ukUUdvBdQYAdxLIJnZWeXUCArS7J3d8SX4bS96AWyRUezdltpMb1xlsJeHBp9Begx4ds9f0dW8n
cyGqqwlRUpxFY/vG5dTUADrQhkOnBL1AYVW7KDAYx0is8zgCcP87tZ5DBW1VyH9dTlN+qsV8t9zv
ZGaFox2zxNuNe7RfME0au/z7OdeVPiomH6YJ4KJJ1DvWbGMek3QCTEFoI0BucrwPJdB/sw15/dXS
Ivb5dUcGrbOXVNHpa7L+cdS05v95nv+nhG8VRjHXBwNtarur7e7NEzZ1R8C1ZBDcRUUMSoKU4SPG
AtKmsB1mgvU2kWiiVd+HzC0gDy/hgu6yE7zhv1kfJlFJCbMzUyLs9Imsa70g/E9f5hjhNDr9z2kc
6VRwOEuy3W5rWO9L5Vm5JMMO+kmrQPjWXu6nhuCHCI02HK2JjE/2hDD0tK2zkZUKE+sDjhDqlncl
Z244y8yrE9Ya3Y41eP0YBQMdyraqkkumrwStqpgdOWlCmtRUh8ygSc+wdEEYE5/wsT/7JxRjLF8H
uweNhhV2lgQS6kcsP6bGyN0s3nazJaHW/XZpuQRtUkhrKfbcdO2FMQylw9cBL0yf5qazQX3ucxYI
5xbg8oeEipYjV0dYWQvP6H/bUGQlh8BZdEwNQaOuLZ3GkP9ZbP/dKcQ40Ra5uX78Xcgf5UaXGlr+
E0e63odThYT8ljHuc4lyq+g49VgHtoRWM+C9rnmb2sO0Fl7fNLlanaLXtG51K/ufYxQ8hm30Qnsl
3Iq+BiiJBwpmk63joduWnh3Jeurx4EIx7tXN8wpAaT1p+b0lZTYuM/01X/cmV8I1O+visynrWHbL
sXBoBUI3eXn/Jvb/RYbG8ROmmy1b9vVLpHQk8yIdebIVnzIkVbS/8wQ+/Nm3bV3dZ+VdVdlbkJ9T
xvudbwq4QcXA9stmHHOHnbNR3Gq1MoWQgbGFDFDQJGtz5jlu4EkAllQuL0GTbVONKJtkXS9xtb0X
7AUjFo9XjsqmkKYzaQJXMMMueMiNh3gwLgqWXbo9sX5nhsLq654eKYFWaIeVjy7AVWL+Q9decu4B
MIIdAfoofAx4bep4w4zRvY8OK7I5KZdotaPkhRGhY95xI+BaHFGZ8iR39XNG+rk2EgMVRmgY7ZCP
7cSDLBlxyELaEL4PXoF4kp2V4T0SAlyN0D+8SrcOanbIIY/M4Uo5qLvk+ExT+LQzFbfkAZ/ox9B6
JUaG3LfGd8r4xt2njegm3+PlU1EK3oSI7GAV2V/CQ0ocr289yhTD86jZnOh4FW0qE8p+38f/ksKV
76rbBQ1TgF2p12RANBZPquZM6cQdTREbBzN1yRL2SkS0BNuQgYIneQBRz6TW61wuVYo9RHCqwR5m
pQZd43WrcLIBK8r2BizACZGDzVXCMX30Vc66UGGtSTME4Kx+IHBak7xaDYCIaAtJLs0qsHsjLPAt
yvHkCmdXHW0S06KzhzX8QTugPymtdVaqARH+sOMADDAdwt3pdOEx9rcjpIoS7jwUs9Ik/7Mm9ZLR
Hy45GAEH0bHVsIN3H0bjoYyKM0XKkqZcAI6z9E/aKF/gXTC+57/3qWHciHY9eCzr2SsXYJPOhpqk
/pqQ6ZjDzRYsp2lstQL5+OxF+DmDkqwXYDH+ROcfmqNEoLnQLMYHLRqNTx6zVPJwRSK6pDQ+L/H0
HeZyd3e2MhTicDJuZDXp/LOZ7BO7627WdpWPx+mGMnduL6YUN4x2K5IHO9iOMcydkiywZnzOk968
HIVWGUNkEBwjO13v8IRNCIuPjR+wTPeGEcd5+UwQj5JDPV6uR1ViQjSkXEak3hvvTMV4ZDKuaxbD
HW2vsJw5j4oW4847d3/JVSlkywfexVOn3oi8G83xGcgaXPwJxY/f396sStdzyrGaZv9YQv9UmsMB
R1RzinglBJvYiojFgsOb/qqAcprcl+c4RxIh/NTazOYu1wjUFDPyjlQgruvq5hrFPupdJPWcRfNq
soXjOXpHfsEt4/A1cdozUbUsbZwtS/Lbmez1+Dr7gJZRPafG5y6IvoqXur9PaciPO2oTNZOmhPNm
NzI8Ed8YaKWsQrL8GwpMrEGIrAHxYdSeg9wWmIWUqWtpit4h4VLkSWaB74JPw/JlLv5co6Q/q4DD
v2IEQZnc9IvYDwmEZfxCEUax/bq0Wbfjua80oo8BEz5P/END75oC9BpMdpDO0g5/Esk70/+gCIGj
RaokjNEIgy0HseRbQp3P4P2duxe+6cqRARM0qqxiDmdmo/0f/cUbat2Raztb0SdhldkqRe3iStls
Lav4W6Dq3z22f1FLjWB+ZH5ip/nvXuXqhm0mthmR4OKI3dTKRweDqjhDbprnJo03kQKXQ57cFwSy
fjzwt9dw5HvYXyYRFBB2C+eFtay6NXnoddnW1qw1lQcCjprVIPcjrYISTMgczcyHxGVDej20/E/Z
JDyzD7Ogpm47gV34EL7AXuRB2uRV2Mq8hYu9AQrzKlT3HcCW2LXnWKsw170+LJrV7UK2ptQpAHhq
UXGShpETmXytaqmgxZ3pSczHAk9bpb1xk19+tlo7DyCEGyt4TBbPdpnAsFBdepjgl617mmOcVTet
CxUY1bwPVtjoOHTGyeRZuZ4vt0dQjoNvMnsXiZLo0reXHj62S9r9MB5+sUErkRcM4BQ2oEjF6+JP
Gub6LuPi4zX/GcliQAHZkMZ95MUfRnsbJu2el0YZxNLCG4LiJoTVBrSkVQNVqV62UufndnrlLv7V
F5lILR7o4oTARP6SYa1ABfNw/XzOITxe0lv7liHWEPvc2Fx76dbSdQ7FlXM9a09qShRsWuPs4qMn
8Sf2nyM3uisy/bDW7hXtWj+3plmxQljjh/aKDMm++OYQ6p8usbjEKKhkFII5ynnZ3BTSNGv7uxBw
nwYvnyMnPMJNutp8Yt93up2XURpxwv7PtRcVk4RptoqvBp1N58IJ/vXM/TZqayTSENcw51osSPWT
QXF/tshdvw7/+0Ee7meCVaVAFdjzZiYbWVU9kQEGQKZXfJ+sLcsF8KVxWHoEbGgVsdLo0LRC6qOZ
Ks4GY14t+DbizaIW6ZVPuBlSwvCt0SZhI1lhXaMSmIMuWVdKcSwYUO3jH8aXgFHeN5evvoHWO/ut
DbHXuBYfN21i41dDwiMNw1VPTcZ9+H5ncbY92i4XDZXGUiIlRpebLFWJYbylGySnsLxkkplrHOk3
EpM+Mm2vuUNddfICFG3uj3JhqUPfu/VN3uut2yi0NxxQh/ttBfotXzXfx/9I06NyrruBMQ+63kyA
FXeNl+yuw0Ccuauy+UcRVub7Zb126n07l1xS3uzoChhuL4c79ud1gkxXEPAE9kIJhoPcg57sI0JA
ZP+KA93+98EMViQFsJ8jBdyJbGJE+RwKrdXXZqWloFTzffrKilWUDL+vNfeMmS3Y9ej+RCAG9aVo
ELPv48CuE/WRZHDkrRJhB5gHfqjIy2oVC9BauBQZu2TdaBzDOotZn8zoNaTvkj0w33zZgA29K+rA
NMFrpjjsHtUIvxIrEMmcLPbn0vaPlFW5aEDLi5eVVhcXsZAJmWeHXfjOM/Fut3j75/Gczxz0mVLG
aJSuz/xvYW0iQCczqXqOUdZCWLQGY8Q/TxbmDLWNMpm/DMwkfdNILeL9W5EXOcJBgrFELnzoKU57
wXKOKARE7GpfsgoN3Otp0NVmlyhQzj+SaNxjJOm+9fPFH2Ak0q/SUCysSrKQnuhr/pzY4Q9zdch/
dlqEI+ZxE8QaHUdTJThRdWm5+Tk0y4BIxvWH3Uj+DyV18yyyiMaFu/lZA7pBzH37fF91KlHGj6As
xhyGPOU5SEP3Udg3dk2LXgWs5AVJkYIjFW1UCmci62B8R80PfoBnHtm68u5fo1LlbovDVQbIeqZs
i5g3jtf/cEIZMZ0P5YyAfBba0C2vQN9j+OvetcrqAmKlbGwMD48Kr9c9aKdERt66QuOtX5tL7tIk
U8s59x7im/i6z/KNkzytmBQkHuBQp0BzkOgC1cESKqhaiKMUPIbD7p4tiuw8LYYACIsUHNFyYiRq
pN59PEOzRbLlAoFMXl4v/WeRdweGwndFh69jt7hgqdeTnrpf47JZwsw31BuWnwj0+Es39izfkmz0
qduRYOAWZXmuumj2ZKSjLHw369//s+zcGWhMich/lgwir5jGAax23XfrieSciq9KbPnwZF9BQNCf
y81Ha/hofn3ID7MXzCCo2t27OolQFWGb8YagXsQ/NGbZ7XIt08bH93h8r+KOv9Z3u6vo+8V64gMO
vfYmqeHml7n6EMk+qTBeHL4lPibSKkru2IrUub4cZaynyK9XokyZnwoOGfWIUlgOE9Mxn9OoRQsV
K8XE95rhDPyxYg8e7p5Ahk83+4rScMPp3eJmkHsacKzRsRA3pL3M3l+YCpfK+oSpX3yT4WxfNp4R
ZNSKJcIva7USpB9NW8QGx+ALq62uZTU0S8wSFldFVCb6FPQRoQRlAw5Qwx/hTLlNVE1h+e38I5FX
sec0n2NhYKhpV78jCm6TCIYTpqgKomV8QDUz+aetIDswR7Mo+Vcmq1pv2zYqev66lvqkmsvEISnt
uOf0ob2uvXLN6VweS2y8v7iqwRAycw1GvwsfS4TO8zMLc2b6ZI84EKokApfB6OukHpRCVmKETsJP
EbnzS+YIeGz2WTc51QVG7GvyDpBgm7zz3TWFTsryl5cKIfEEpqssoaoWUgwDUxy0sAIuZlGEL5Rs
nZFoL32dj613td41SUQV1ndN3Ij1de0nejadoz/t4jzf4HqzQ2BB5sWzsSH/mNEzrGVNYev9osf4
YM6BMOaBNy7VmaCmyJPjyJLj0vAvC37jaHmHOdaZjw826ATO5G7ckMkdj9lii9yHbYD+YKyRr6Gh
/k6p4Q2Xd9YoJCxvEsCyIIYZDNQcfcYwHn9nhDSP301BJIqt4eSpBjE9FG84a2GSCrz/UGissBdO
uPPyWykUPNj4rQ8L4Js+WpSXSTmsfmWYNzkMiQw07cDjXihrOVx/CgapXlHibzC/B97ry36MzOUE
q3UE+yKoG5szUc+KoKRfA7RLfZjr2e+66Za9OCJJJ8T69CKadiBWnqBE3ujGe7pkoPIzo7aK/Wz2
0QELy+s6pd+leCajDuYoZ+zz3a2qRSAbkXql5EOe8F5vzTMNVcEwJcgFUerBM0qEuB/dF5u1kxKV
swaDXfa8Kn1h/VuvI6viouI4gcnoC2ckpz1qA0li+1wMTBZuINGvcKADZJL1sPO+ZfapXyhWZq/U
ejqx/6F6OGuDL+AXsUKaqrhD8Yfgizzer/YrCrA9WIufxVZS0Ha15BL9ghmfg57wKQ+GcERm/pEk
jEdvivwsEBxuS0W87Z45Rm7jD2x9fPG1aRENK+pGi/fmYADUyTFfI7uy6w83/P0DPnfNCndaGzWC
nGSACGfmJq/zK4AZwvNY0Y7rvORmbNxry5CnYfMkbT0N66DZuFO18E13XxH84dbUewVicam6Ou3f
bqYZhkHPWC6riNiMocOezTlJMRiISMhFrdbREAvfNiYivJvtA1FuJTXLDOmaoY0zWkerEWpACAim
u3dr5ViUMmVpOU+Td3PI43lQyk9aTJVOE34Px4+28j+O2LuU59NvP/Ogn1ajObMhS7j+cRhVA1EH
Kubu1IDEvqEdxEnq5h9Z40wjG3yRz12xZ9LEnnFzgLp5qpDEE+I37xrgPMeiloSLsdUSfQBhDiYc
Duta8qfm2TkWK20SOxHSH+R84Vg+JWSI7YZ60fWoYz7ADDuYEo//H0AzXa6lSnhD1mqm5b3oY+7i
tfGXOFOImLgblgw2C+oUisU63wQvJJhqGRSQSR4SsXQxKVeYGQKTZad1vB9U6YC3hIOG8cYPfu1u
bB5inQJQlFpGe9+MNqXzF17OS6UFTfWh4ZrzVayuwVW73FZ3t/HwwHsgtkRCg85jUhsP9/vkBH9w
oPaMG4T+cBwIRSnO3v1miUUSNuMO+8lP3EjSJp6XOQzHtUT9iVtH2Vx8YaM5dFELL4nFnAZ1LCFu
OS8jLg5zLiKl0j6MwSuf7AcK9iRzKNGuvJ7eMi46OYvX+b803SEZpr+KeQx4++EKuC3MTeiO/LZD
4kz8DoNA41V8NojPznE/wj0FK5yRV8c54LGz8AVNYwOl96xMxrDRFjRJe3xAaN07cqgVmu76Tlon
37irLb4Ai3RFsbz8383vjb1YzRm24BYBpIo1yjh7d9+2WOoD1OHuHfq9AHSJ54wYmy6VSmdcpsvr
UA6jpH5g0HlPYrxiMHSz9pY7P1a+GaR+jtCmiVJ2JqDF1GKU3k403xqYeQRiUe9YqyEmBnsNszem
hgWEOPyoAwnz1gWICmWpVH3hvaB6qoqIqsoqkBPwOhhRneVR5JXaSdCiIaCEOjJZqp5DdOYevluc
9fd3VPHYQsdnEJ2Zz36IVOp82HA+0N7LT1K09DS8tFPNluUSl9+4JxAJUHvgi1kv35j6Sgxj5UO4
oicpIhWjksaKk04rsL+fH/SZ9taFr21LLpuzfnpQsB6PhQqWVxl1MR2bsYVmb3EJGBRIL6n6nBsj
rrlKZLV2Qf1K6U488jkVWB0eeHW5CnggB/BeK1NNVTvQ6q3cr6l49TN7pJTWcegpAxFaAHJHQ8MO
Y2Ci2Syh4n/ep2oysSgJPmsUZE0otnXcrZ+PI/GhXhpxOPZSiNacndSYo8mB6siq1l/P9sb1mXRU
SGpgTtdZUeToDLdA4K1Kx7eITAZxqSkIXFQdY1OhpjBKW0WPEMOusPhYurhSQ27SVVe0WjK0GlAV
/5ukuYtvasQPIPMiax7wwkRiHQYv8XmnYMhV97PczHdUd+JEPw9UWG/cO0KJD0isGOrn3kn52LCo
DwnaMw0jNyj+x2xquchEJGvSbYBGN3+qDnzVlq3rt1AKZ3fiB4TTxAWKgqB+cksy5O6XU6jAm5sL
Z8V2pReAXdPxNJBN9o4Ougr4VxdzegNoODjYAwOQbzgeuCWcGQfDREy/apNuPW83Ji68xSuWOdU5
NX8cMvOQJihxVRtFrzO8/TMrOmYxuoONjErD9NEjKgD1/LCNi6kiQ6eF53Tvclzot1dVcMf+ytzs
2bV27jIm8huT+z/p9tq8L0gjk+PtBPEuh+yCd8N2TW7bWugzoghax68kY6pb+Dcwjuo7KXNfNYr4
b4Z0Z2R9sAj0mYmatsiTfvfySi85NzCrS/bGMsEcdfhKPXlPPVFic7rIArJsHhpzy6aXFky47pMM
iic25P39ZxLx5SwctA87jI/pjsEgHT1sLIQF/3nhUFeGUKo0arviftSLugMBX6dF9bdtWx4MvDBK
456CtRVwoKX44tcevz8J+ticSJhOd79+5l9nIOw1KLIfWhXbWzx+ngZXqocEJYE2fnk3PFZFuh7U
8vntOs/EfFgW3qXMG8t51sGpELXsEjUqBjEUrnW5hQbybvvCuPOkd0TNkO4qPhwW4BkCTCfR+VpN
rD5pvo6bIrxZAbYa7P0WCfUShcxCJJ1zWP6WC2rsD8rCm5SMOZzvHj5ohtBl10C5c77tQFOfgY/u
DVoo4BOw0xOAnhh0MKcdN71ht235NQwZBrafRRKPllmwzZ5ugC7TldkXAClHyFNDSw9prZgctIhb
RT0kNaKcR4dAvc3nzfe/74hDTZMMKxjrN64fJdY4lgqJwvXbH6hBjrzEi+5PfxJccVLshrmOB4SZ
hc9DZDHBRjLqDMA8ysTqhh2X9ZODfyMtZ4vsvSYx+AlgNU1tNUyBoPcHh7Z62Qkl+aCAX22p+k7X
irmSNKzNq2UsgewyuxhmQ7L4GhH8tqnjI+eWGezm9BCvKg8H07yw1v49fqAh/gjWA3Eq7u8FGR9D
nD80q7TOmA+LjIOXmk2A2442LVLBwmwRaX2gO8O8mMsym5jU6nBxRkMpjDjUeHTzAXMlp5bc3OrY
ZssMY4TF0rOkVyoPbvs+DAsDX3tbAiJTPv3Dot2M3cilNctixY3ChqH++AkTdO0/aYWmjWbrAynb
Is3eSOOnEV3FGGDzM4VGSAqNFGS7mQk0zQranRxApnlfz4pAAdCjnHzvVFKJHNrGAKdhhpXjCCIc
fhaE+EUhbQTXeh8pEW3vdMsmdE46QcOLGQxli5KIUIno8WFXghFXbABx7nAQODsy/miw9j4M1voV
eJrccsE7rTvOTkGODicaI595Cgu5GllKT1d18yCdqs0BlBSs1qtQjqqnwveKjxy3QSbVCd3IOVMh
Ve0ACfSHSPRDO9Ah5nHbGx/xemOIiti7MUI/shLB7472shpqWWH6DKHBcRdxUX0xHKz9jurZjl36
O2iLq03WFjG10auP9ZwA/7I6i4dUo3EabGx84aebzEbB+RnfZmoqM1p2mhiaCUVHJKm7JvRvH6Ig
O/yMW8bl5bd15DP5RJ/X4f0I1pfsVFIguoCOuBPqBbLO6UaYTPj63J6zo+a51wuhYB4J1uYsaKJL
UEHxfwdBlYgNLDraw5bbthMorXeiuvirwRePseS/81eq3AnMgcXsBwg9gYEdOVRrkhDuw7FnYj+j
4YzzjMDcT67+IfcxWlvyltfQ/QUnBU3yL3n0pfoq0bzuSYwnx7ZeVpR2Jgk++mpVg+QpV6ib/ydV
AvAkL1/3LYXoD8JmaNLHHVWZbsEu7aEG4Ys6A8Yg1dSa+olmZBmKYA4Tex6HWDx48OZ+tYJtxmx/
+BmhyDDwmXbWoy09s2sdJYp9gpUtfAev43bqp6/3AkqX3TcZL0T2BuKf038k9CNrd/njvHsyyfnd
1SMuLG/mK43lOR+N0LzyUcrqVcHGDJl789zQjlIiNdzBU0TXYPL9XHvnN/COUsgvR0ETKOZ4K8FN
q8w7AR0YkWoFu5esJKjMIG/bdOeRLVwaUvHs2YFKe5hH+XVNi5IzCzb9WXhkQu8ufLmKTfbKiUN+
qrxAelLNPh4cQDkyIt8a0XgxGYB093PLla2NFoFYs+V/U0QxY9Sexlkp3vPpX53U29UX8W6bHJ3s
9pCRaif0NBouPCIx3SpSQBGeJf8MR5B8pCDxm8x2Q37W7eNYShb75jzJux5LGVLFPw7jxXVrocwp
eI9ifRnOlbCShRxvpJ6EznaTbhpBo2ML5YSjydFVZdOv/xJ2cmbdStGY0YlqS7wmLwnRR2Nmtv7Z
S0CEEY++0tUfWvwkFXZy1R+gSd7FkJ6xJNxqkGDQvdRRMSUwPMxxLF/yt4MI49kmceJd5dvflR/a
2dcjvaHECuPUrxgxPpxDs3CBK7LRCbw1hrRSs5xT5kmlOWyb23sEZicU4qz3iEVa8v3VgK6flBf1
mY7UPTVCtrS5B6wDdyPnELb9KsGvsUBFMHVkYVUFyZ631PJI7LN33NiUkPHuQix+S1w6fsjZoQkc
/KuZz6I/j+S15iX2fKjvF8Y+/RQIgPP5xO8veHzvPDo8OI2nAf+1v53/b8u9P3T4Ft4cndJylxrL
4lkREMH98a6YBr+dx6FB0QGTc2Hox+s7TWaBEVxSt3Ldm3TRexh1oWJ3gIiEbqxuiw1NDwMQhG74
GNZqDW1/gqVPoE/CmiEN75ykPo/O4/SfkoknorDroSR3iGNTDvB6/boWaMCmYJzJlDR+Ba+WrQlO
cmMqMJVVAw8AFyDWQZYi2HSDmkA10Rrn0/0YQWrulfr9fFG7gID1WsvXFs71EKFb3yvn2FS+DAqO
RUWx9bNSBt0RRjLEWj4m2CFlZj+FgNeFmwS+hQfNuRp5XeeTaNwIz0Io21BnAq/y5nnw9Vo8bwa1
nD24p1C5w6IyLvIB2OMggt2pGyGkHDP/DocGgLBQWkoJOesdqeCFg8xVoWMd8DOjbDGIiK7hRbTP
0QUCb9hB3qSF1dQyzR0tLLshU6q4blpYp86yYUEWi/gt5OQS4dWw3ZzazEvK9vOyl6f0HHDvZKuM
fpzwp/q+bvKNNjmr0T9UGZd6ZazoVPh/BDHVGdWF85DT8VWS/VeKRfOF4Caf2BIDLh+9LyX0oULI
j4r1KpK/neVvtME8nlRRCaImu9gZp+chO6XW0EUVGL8pyqBQNa6M/CnTapLhBg4jPoDMyshZBgWq
sHH6hG+0bultbAy17fELYa+ylyko6jIHSirVTeVEpDHW2VZn16uTtZlhwXinwDhFxnEagGObJE1z
5WOqihzUU8ybmpDlQT+08xzsu52azU85BbeZFQTHXqKU/OfPMKBTyopBJd49d562RsW3GKKTndxY
LTEL2WEY5EAj8uYeLeT8rIbaBhGZZDVNdl9HT8qY9RE+5LBxok7BIJusj1vaMbCcSLT11cFqfDtH
n4D4/HBxwa1qB5YtFD9lQfu2Jwnd82JaweJ4Bo2lk8exMhvdV18v529sA/DFoxL3Am2MXeoxW0gj
HAoNFR0nV0dXnqN5t/IgW44Kr+gOiEJK+ZrcCNCZbAQV5YaB/Up01yLd3IUhGZfD1HLJzpWaVU0J
U+DInphcYloPVw2BosZpJfuLMexwqJxGyyjExkRdzXMjaJWcqJ45AN3Nnnu2C3/mH/iUyZzwngq5
u/UzYLa/xFTEAbmBwJDqVdiIQy7JeqguQ9Wz54xQyYS3F3Wl8RD9576EBk6GOEqkWIMzHxT11zIn
uTKZxcb951M9u7Vhn4Z+BAPP0N+tZkHhfLNeCGG+BQ1zFE2ZBC9a2B0S3/x/1oRTqHN9rFUONmB7
4RtMpttKZ4WHdenGiOKvETuheEQfoloHgmSuQiWRltxE6cC9m0sGeKjdzsJfi6AjXw/1Q/KaFe5Q
xFywKi0Z+gSx9ahljxBnXYQWqy6jYzrypIPjTHPhwG/sy1wsEzO+i1iUmw2fVF/X1xW1vbvFEaTh
g1ygNSf6O/xLH9xE4tc1XxFYjl9sG8bnjHB2Csc+Mouo+zPwsFCWs9eqR4KkGD2WgVVmE+km/f8y
3my4nLQ+6cGzti/Yk2ij43LCmRVb1wCXqf78c7JvPMld8I2I3oPIR5ndPy4wEUvlTq4jxbxYnr7F
crVV2K4mfjRD0aybx61G6az+bgfIf+TaR6Ph4pfv/ZnJUalJ76EsqWLXg/TOuuPGV0D1kaCVptN+
qcFNVzR7A/eBc8xZNx2wx2jI+dasD5fkX1lf2G/Z4W95lO1GbfiLyxQOsAX7LQ2rTNn7nOcBxR+v
FvFpgVVfVHz6RX+pRI2WsKibiwCUuPiJ+k4Sd4FqoMQV7Jt7Qr8Rb/jPZH4/luTR/uQtPYyJJpaX
58UZ1zNAjH3HC23nfQzh0D9dglPcQr1QG33O+T1pG/S+zG8tLtSC5h2GuNDUSdkgMnLDqAxIR/RP
I7KbDsaDP0cMry/Jxlko2f07a5v3XXnBp/yl1fz9v1XtooLWkd+P8vqUJdoUQ1A18LGJbl8zBU20
YHDvgRgD6tT+eaKxiUdgHuqSbKF3AgX0fuBjsT6fmcDuAYgzjunUk4NSTEapz+ovlTP8dDxmilNM
vfJfpv0Xadnd2AEuJsbajaPefLEojo5dU/IAisVFN04QJMloJWjW8dKcvohep3p+9GBPqGpVUpys
HJxOh2qJsHbI3Uw2tHbsdii3cWr0P2ZtLumLclJQK1jr973BUO9h/4wijh0ydAQDz6fKf94SHO51
yG/UOtzmpCTVxwfAPSiQS1B0qCeVZJnyzn5rzEy+XUy2bX2rhXRa9g4PGirRheY39yo9237VhRXV
T1PnkoyaW3XiJw/IaKs4kksaU1YfOhRUtN6toA0QnD8rzubGrQxyRK+CTOUlAt0w43JeJgEhPOlP
oVngNVQzlY9XHtcemet53VAe3+9gm6QU/SHAITmhG8ECIPxxrlSO4G3DmpG6+v5TgEib9u2Yc9Br
L4dGqmQ8ZevPD72GzrNivLj5GclMCoiRXlXw7UddWBXusyQxj/Bmqf6WypyF3SQuF3BX2ufkSZiq
6U1HpugIYIXnCu1KzfHlkO4SO5paenJ5uEb8f8l6q3oR/r9P3Z3C6etfPEDQLlE+3dtSjyJXOupL
o6mgYcpTujf0AHf6jCioQq4JGO18M/PHpzoIMAcbozo6sM6Z8K/rDpILHbgX481t0v/SrtHqyJ4n
WJFgLPGTzpDKjVAA4Lf3Sml4jO1myBqAlTx3f80L+Y4lbwqGPeb07UBAxWzstTYCQC5Yin0s7iYJ
bmEzVW5+t5ez+WfyjY6SCoipTdqqRF4jFzYubdTFVn/E5C/c0Ti7dTwNt4Yc9fWlKXFiYULMYPJP
4uW+Hhlpf36TLRiiCV8Ymt5gMByxgtVmsiF4TlFIIa+u+2tX9uymcpf6QKr99oCN9xxnC1uIy4th
i1hm5FBCuvYMQ+J1RjIlV9ETkAhTi+Kh/zLHCaEIy0CGdpJxPO4w01UdMpEu5DSlgLy6wNc7KzJb
YoBCKKUh7CPwAjj4j2El5Xrt9UUmnJbsqEtUX4FJ/TZjULxGy38DWpLG9diNt8viFTaWrK+z1RX8
Obw1pN6AR0OxRq5dJ+1CZ6NTf55hyrD8tC8H514sk+AiR3uPURhUSKN2S72LvaSJ7L+5ijqbi3F2
VZEPuRYnSaQbNxJb7BhLAqTtZojqgwiH3hixq5NYMDctSrJEJffO7b4k6+zW/Lqf9ipPSDFBd/x7
2aq6y+47fzwvqgUTEetB8EYkfs8LpZ9465Rmo37dqlnt6sQsjRBigpDgYYMGjo/iXBkhcCc4ACUg
zmWlINM6Z3HK/wT7JDdzK/AUWX2GiBPft/O7+5R5CgGfzwWYP2sCvD0ZvQ3bn/RcS8eQmq95so8X
Hbojn6nM0Cx1WzFlNwohWMqiAWKQRS+3OTqsbw+ecBMzTFfBFxWXNahU5DXmkitfmlH/x+spJGqZ
QqpUsAmW9pPdMKTCqBdXgUDWN6TEs1U5AwngAnGOmvmNtkM4xmMiXHk2tOhp7eKFeaMeofZbijiA
VLJUJLRDu8tGHb0hkOD4ZookLusLNgKLeyOKtjadGKWdod8cMLXsGw85WWFO+Re3vD2fExSWScmC
TDyR5/GMjl7DCmuIIHwRAiGwutWtzHnevPq5/Gcv3hODi6F71M9Riz72KYsb3jyM9QhBwt8D1PNm
S9NeK3d2NEJVyeT93dJP4WVyitkLwTCWuQlkfAsOIZrZBqxjBhICEawahMpRV/xu9h8AeCKKJ02c
Fmyudk0ZJxJGFZKEYF4giRCBugD6urdbQ+nDfWeIhITHZQYriDCowhsI+obUQaL7Vrq7yIgOcrLg
SO2e/U0pdBX/hbbTniXWsBHPDr1znEIvI2Ijl+nf5BX5FhODmEa4VKv5smduBOP3pqEfHaqB28dY
P9mZADIrDfaIYViPz9S8Fl+yimE/sfDM4fz3nkTwl26unr8f5lK61GY0xesNAeYLLbI32ncrMtq+
w8XJPEGpyeJQXhh7cBHO4dSPLmf9J5kJv+l5xWAhJOri/1R7as4Qog9vb0h6sCDPi8hrHXwxgz5L
Zby6gqCCq6wTkj3FlmVogHchz+kvgb0oenNZr3d2n3g4v86dZwYCw0dOSAhIIoIKBUPls3LDlDX6
x1SeBj/5zUvrBIStlPi6KRv0vz5id98XtAHP6hVgdG1YEZI8zO+wh6OVkfAanwrwVZHUVlZRI7Yy
hgxeWguzq4sTj+4ECBIhoxmh9/+Bw0pCbGGxH4Kzkm4uPvzk2zGzIC/hNDOGmC6LhjQ/NKhz9oD0
oSu6e9dLQE1lHHrK/BSwHPdP+yjL/N4ZdkiqpVJwJmlFhurRMPqjAkUvCLPOFTZwp7CtDUeszb8v
uRMYkMKnjW//MEELFuWH56bD/vYB/W1eiEh3vtx+txsw4tsD09X+QUjfyv2xCsnhiG83eYWvcUMa
RTIMEYzNqvi5HP5chNROFw4odzvfSs/hDlrHoZpDj1AqjWCUQctIRHHMQO/xede3jkgOqVuDnSl+
2fdkqwlwaUVXG8yeskiy7our3ZAk46LIC+SKWDNr0ql/PInpmx641CLZNmFB2J4oiC8UI3PfNE4k
+lEqGos5xSwVrUK8RXpP9zuqxqDONiWrAigkWU6vq5kOjU8/e8Q+MSrpwfNQsN/Q4cp4dT1JohA6
Fr80REbomnbvm6ybfnuFIh10tm1xkDFYZrYjrlMSt5lx7PAe97i92P1FD9m3m4Nph0cgPzf/0YzL
6cmcZvJpaXOw2BpYYTC3CY/iVF+nxW59uFhA5mZF1g/50Z3eSBUw8COZssIA5n0nJNPoRllfDECs
NM9Bf3QwJfLKb8rBr96UIBtMzQmqXaDxMH4skjfOQczMAtOhn7WiDgldiEWYOtEukuoE2xTarO+n
X9hY9PfRht0j+6fvTvUwrxczgBrk/giwyKvIIxiTGEnhfcZwbg34iF57QozytUOdPD0JL+IWr0QH
2s7mmXvx8pmlZCM3x+wttN8JU+uhz94Hp7BKqASo5r/Q0JOhCBc0FS+pE0yWHy5qy6kKSSBor/vu
P0kabr1uYP6igHtUeVwv8VGgj3xNIaSnwv2qGXeKZYgIv9y6eTvaoN2oprzOeILHq5vjeREkTKSy
isLJZnP5dIF+oe+R1oJI74kHJBOwaboSCibuPOHCmSD1Ll/cV+2HQBGRnJCLV3WFp4z+3o3X93q7
1F2q1fOCxFVRO9Ov/7HkDh2NJT3iBz0JOftnqYyKLZbdh0+rbpYB/7fapj9okFMB6mlI5fA9wINt
3xJnw3nmf36+K/UKWsWXVMWR+DrnXdOQNYhm96t5Bxbta9ZONtlgiAPo4aUQbNCXhsXv7Iur1fzZ
TudtA6oSLMx4YnGPuXwzudPeOXhYG3e7O/1rfcTVhU8KUFwsed8UvVhzRzJSX165fyRvKP3/AT2+
4GVL+QgglcN5xfkXOjMnZWy9u3rbBnM7BKYFSnkIsdFIOOs2/pUoV+oq7RIHHJjSjQyuxTf5HMc5
8KKRx2/epTShP9Us3hMd0eCPxfKhrYKBQ9AoC5sZDfL+D0JdPOOHxpzze7ZuCF3TY03vzMrP2UVq
rECSLpE5QbfekKRzl8aYtwdrw7byyDnvxb3/1X1cFyP5QCwRxxr4coQuCZS0fOEoUtfGu2saUgiu
QTHJ8J2cJbPYJD3n+mE3+mkMtworelKE6SjQHND5/+KkAljx4CAQJzmBBmpUXT8t52zxudGVQxuW
NXYepMtYQIzNVNAZgW4VJkDzIi0NVUqgkEli/83VeTn7wmkLtZIczlNPNDxYbLCRNKdE+U/rqUjV
NBDhF/clVLSMKYBWW0boWkG4tWVVyzqIYFLF8+y2qmd0LSU3xEBk6/a42XWc1z39K8EQgCG1Pcpp
xm3HywjoFAMKObiwKr3B7WraqgRb4RmZmACTjzvhDppkYlxBE1hrpkitoFbZZAofDalmB0wFBUem
FLhfMclQSA5sUHOZZr6o58caPIokMiY/9wT3irID5UMr4nVKGJG52zwS8rA1YRN4j5drnHiko3sZ
QRhdyEJ/BxHaFyLiBrcWlV2ChFPSkCNGtDJsc8lsa2SkpDKPNV3jKT32YiLhRFDym4tAxAUwEiwB
m1T4e0x8/M2yJG7rNcK0s6i0RRowlWY3E8Ma+j2YHOb2mzbU2Iu4Oq8AlBm9kJMLadjJQoROx4Ml
jfN++mLcBQ531fLbUx1+LZRTia6Pa8z5yN0zgrI+TR9DrIrDVXD2acjdSnuH0kmYi+iTxASF2Erp
BErIeSOTze8xH8prB7ZTwHqZDfpdxKzDT2iT2Vomhlf9ZAYcy8DHBUp1UbM9okEeo+0uqC1pOpIZ
t5KRxjmyRp5+ANwvRMbQ/67vbLKWhWQq1BS78w6ayfRaGG2NYVKELZYS22GAnxcE1PzgLIPaz1nj
nUWAxD9kLFKQpaVLsqahvOcqH5wKU2Zw5fdNN9SVd6y1ozoC1y90v5loySFNcFyOuRHx4anMLKi2
sadFBiFy5Tg8TtdpKpxWJIXeugxHAm9U5lzjWr3eVrX8AvV159MYGdAWCzIqUTzfxSptFwbXIUZP
264BVIOrzL8ep5VUTYO0htjOmPT147vrPp0jjNI/vG8F2AB/oE7rM3cnS1s8GgoSFoNa7VFjQNXP
TbDMkLfYU+4R/q9GI5kbly4oa0BX2ZKRgIn1MmiAId/xbP7LXQO9YaMlkUhhKBoY9WgmWuuiCdD8
ERKaK6VrlQ9ohUI6uR45rJB5RTcTNF75KZ0vsQ9KDwJ/p2VAFBDX8xyOHTO11khJqBtcolNUooxk
fsfPSjw7Bws55aOM8HwdbpirPpzos2Enk54rsLarmB+iTheaO/UeJ39qKwa98gT5Y4B/ZeKvQKSF
t/yRe1JXiMDkujYMQTwpOSx4mL/ENUniO4IHoOQHaTpd9q3jnOnjD2Qtw1OExmCJLDW+BmwWtHzs
PclCtE3Yu+LwNgRA1cXJUo3LbGY6eJGcJJf5O0emm97EsfO0OMMmIIXO2ohj3C533wShxCP4O1nt
yJ/Y6mv4N2SlBwN0brJmp5efMC5pM4vk3APrs+mA1yOEh42JX0Cj2NDub74b8Sc8DDdxKWh1i44b
4pMiYB1w5YQvKbh8WtpcJxbX6WbLC55XZDxkoAp2igUtMThtxPoxXK3dUFNgyqAnEey7aYT1VMeR
oPAH3cONLrPNW2mkiK/xdtlAgrWe1YeXUwXcaowKSxq2mMZWXz5XI5MOUHEcw2o/sKYWEsciAn/G
q2Q9RmTvfywdCcVBdjRxc77eQ08ki9qVlxTl7JgddMMilv7R0PLB4NE5GgmsfOoCGEM/V6vRgXHF
2nBvd6l0YCl7/9Q4aVyYzurTsQd7ljY/1RW1g70ZSvnbZNzVAu5l5teBEqka46uVEdlsdktTa4t5
SJRG8+mWySRRd2nbvid5omgSdN5udvY2oHRE/s3nQNe/MiGRPuzPXAR9zC/mqyA2MIuvB+f9LV2q
g8D+cdRStvBW80FlGG1iVzhZjSeC+vQ15g2LIqWhwWxXD58dyh++UGnKXXg0tibQ6k1ttqcGuDNY
NOhx1XKUKvr76vmPNAA4l0OuMzHG7hwsEFtYIA/5jYdY8rmkFYQT9pKJopQ5k1PbEi7/9yswp+fY
cY9zO1zjYALUx8dinOiNkl8mVoEbZBCS4UPXCxVW+04lU826wwkha4xL0ZJlqcA64caXHqULznql
q1QjwBEnUPDP3edDLRp7/HGaFUPYPmrBVwtTAdGZ6zlBUMpOGnfdzEPk/ZZZbA/CYofTPqFlacmH
sVJYjgHjcHZTEvJfurxwxEoNhStv7HexDNLabOQqKC+eXdYRU2Om2qaKJoXAwXzUQV03pMGJ+QPg
XkJl76AxkFBZNWL+XuO+wC8bzIinIofYORM+kyQ3/9sVFDzWvXNoX8jI86ya3IE6qzuK/71yKOf/
AREDWWwge7ZnU1z7I8zpZVlj0N3YaYt4PzHarV9KOVQgG2VvfFKWL5G9qokaXsByQKsSWfHIZPc4
1+ufGtBbu98EZI8z7wiR9RiVZ797dFKCM4T8W5h59uURwfcrgCJuOVQzYzqaJUzy+U7heJPORoAY
O225ShHsmbgF5G0CwEp64QYvw9FPvIaCwpbs5u9zkES5Sf4rPKpYxnb2P3zh2ujPnCGo4488oCOU
DVddzZDgWVLCazMrGzGl4ohMh9OP0LYa0dcj+xofxcsSX/y7VWiduvQFfKwGTy6ify6Chk+KFt9N
MJ69SY9O3jNY0pcGTXnxeCHiMztBhpbW65OzFcSiV0S+q5pfMJ1kUM6TWNDeUnIkHrMHWu44IIq+
ghlYa24RTC6sS2vwzhugNcriCA3sq8wWEOLgDDhC5lMKtuAWGc65mAJu/kDiTjhC3NbRv42Exgio
tXeY14Ryh9RX1rFvdJIRlC+6Uzhipq5nhpHN1xdbDz2tKbQE13MvGZT5lt/bGKffPgyWaRQAh6UI
88mbWSiXF5yujQtIuuK2YPiFWR0N/lHll41pdjioBRPnGu1CiJvXYxYEZ4zniAHt64mGENKYpkHx
UgxsKtFjDTgwHTpEyhfFJYrzbwOAMYQiZBs0zUYAcPx6YlDIBPlsvqi6Z/RUKFYpnDeCosbM9z8L
ddSsHgV4LwaGS6aATEtBP7epFtDJ2Vnxun2x1wFLffHC4AB3GBC5ig8C7O5zuUHEKuQZB+E0+MKz
oZdIJl2OADRhcQplvVzWAXyhuuPGvd0HyWb8aT8CsQeJoXY+WFPcENuiSPl6k63Ta12lSpHoYST7
zcvBiaWRv0BajqrQUmhYgVKXjXs7Ibl1W7xcx4qGAXppMJ7Ye9K4kIpq26H9U1aueBGhzQqeGm7d
0gsy1vQ88q6AQVapd7oL5DiFe9+lGBucNOiGvvFLe0DzM1l8BsuxrC0vUUfqlx2gX9jjveqLQ9Wr
BCkCJ+n5tpTjRocOrtOc9uLfoSl2HyRlQh+ZS9pxsCo0f1UEpeLYdN31XSKu24XvKUOkg9Y7eSTG
yOpjNpphEf8xR+RHVU7NRG8JiXOD559R7twu1Di97EcsXedADRGnkw45AMpx0COBBliNhBpzq7fg
kvYYu1tPueSF6ixvaLsXPRqDhoFZSREljuJ+ozqeuSfVktJYeZeB1mup4uTJ8fMUnDGxaG0zhE3X
u0+l/sen+0zt1hKZKdCk8jrZd4678XeD6v30fDQduSx9JgoxJrcmlkTan4MpYIBOVCN1j4n6kc13
NM2TYMq0RTG1X7RKGTiQDZaqdLfr/kgUjqF33jpfVPKzMkumertzyqfzLQrFO5hF3eHCbFT8V+Ic
R6D4s8F8HO+wy31NHtcYhm+2e+LFc6cNUNDfcCJg9wDy2oxvcfxDLXZ7qlcS3r1CeBRQ56xWS1eG
i1u3q2A54ESAJptlAX1XShotGjEngMfK6QQBR6DR/T+KUhbqTag7uB/dTswYHq7NrCw2dlvaiqGb
p+35ih+vhydJllhKWFVwX7Ma407uSdWIDjDp/VnFXLde9Q72RnloQLDdD/NFhDSsw7slx0ZZpuS5
liihnOk4Fr1miOCGjqkLibolp1v0CWAO7fxZ7l6sxbyiaNqC501wWQIJubkkn7DNtNg8VqHoBzqQ
8ZUff569HdLRFr7E18+VCTVILxxLXhK+nzVe0dVr/7dIlhQOQHrGq+N5mm9BbGazJaLoGvL0RVgj
budXx/3e0w7pp4vnPj6D205bJlMMBhee+pu3uvoUlzkCon8BnC3UfcjmfmQEiItTm9Dh9SqDVER5
wK4okQJxzoThR7aSz09HBjiFGN5SQ7KAAuA/1Eq94FQVKquuz6qoXw4XdPhfHhMFJjqNKU9TeQEk
ca69jYgyUXhpPDTLtymBtS6Pk0Zcd6/3driCmraC0Gg8Ntbju2Hl+xzt0QEA0WWg0hbWgyxrcTvd
RbJUR+rFeoI3cuxS3tgM9hYHCQpuFKczAwBB+kgOJ966WupiYGv32xdOQ047HzWvDPp6S9kzY6HO
e8G/PKelnnZAgdSPh8np6e0/NqovHt0T358xXFDXl3HMGv8FazsVtNHDb/Gsga8O9fvUluwaKaiq
HLQ3fP3ee3k7QqkIquxIyGI0dMVinxiAV7uXLx1/x6RKDymHhDx7n+BrDNM8D5vuZ36OMed9zvID
LkG01dige72C3pv9LnUs9oiHLegf9jBHpmDJ1lfqnu+7rZg68XvyNHoiqx0ws94udk8FMyMn+HIl
uwMpInlLWPLSa38duQZDlf7Jwnv7NcJkGz2Oo8QH6zmBABVDcKbiSnVEkmrFtL7367n8cEA4JCAZ
c7Z7608XgMhTAletltUNBYPIWB3c3cVhhGI9+G9kyAXyNSPP8MWOr/p37I1DoB56jEWY2NzogKNz
vrvMv/1taJGsnxT5MA7wxKJCcwnwglhjeqWLmiJ3c4OWVi2HZBvd+UOXgVUSfJUSidLMno2LRPL6
JpmaNkCHpBy4G/qcfs2lre7Mi+ZF+khDvSeVcUDOOvDslVMwREgoLM3qWTQU+XIJe9AaoLLFoyeT
VopS4LDVDgOLTdxrfDPw+F0iF0TH5cu3RXppuAdI3fcZo066YWPbYOq33AEoMBF/k+TbRS8RKu9U
MvjJxd+3j2vI8/eO4g0jgWNqfMQNCquRfv5D2jJWCwjW/gma1yc6HMhofTnu4d64Wv7Z8pOCFrS5
BvWZrRz+Zrwf82tUryTriclbxWr2Qi1G77UZXF0QLFr6dVBB8gXyc6kQaLmDqodNvhc/4op6EaIs
SjZKySIhOQaXqugmElXp6JS4H9c33C3gBgkwRPvzmXJMsuxVGIoemVrT2FWwFVEXNgEudOPVt62Q
SRQok+tAkksyS2obaUAjYs7uiE24BxIPZSaYpV5QbThrMi4D8+V0gJHzUaLQhRvpaO9WfM2slmGm
zF4/Y7d7vwj2Wp9JokxMuSETDIWyeg0WqP3IDkz/4J2TXoWGpWIU9DlcHi0mlPIl3k/CZVuvAn4h
TALjltHBV3kSeAKdkyxtL4B0HIZNZr0R07vrJ03sTgZ+RU+5liodXjo8rnelCk+FKxGeho00eLkT
PruIYw153gY9zkBCG8mqBu7rPuY2g788TaUGoCxhlox7FRFm3z37CKsizsifC3BNsvBDwchZZQX8
6CS7jSRJg3K3gMTF/wj8QAEWbzQ1wepXKfI1q8PwPGsVNXHHbhsf2o/qhjuP65Ca1Zyo5L9QNVd6
a17lxM5soM7IjhOy2bJIEc10JceJ4RTaWAGYQ2gx/+cPdFxc9lmR3ZYX8G+hozIxjVDHW/NKiP76
e3VSuzipavBC1pKkQgXJdOcnI6yT4N9yNDthkncK6tqxmMKyWVN7tVQNAHJjWg9IlfqxRow6kOCL
mhH25syquVJvUG9/pP98B5E5phs5fizDHfGUaggjEr1Ocn4onsqwUVZCoThDYJr/YSb+Evbw0A/1
zV7I1wilBg5Mw/3v706t2x3azZRJAQh+dVhpliFKkVLU2qexRWZ3jjQMCvlmZvOItJP7T+ntAbDc
VxtlliwPuk6lbW0B5JG11jhAft6ScykVKkSvzuoL8wGTPRGBzhFfutueONUYLApzyl0Z2asd/sdf
llNgYKx4o2xkHaHaGDJy6gyO8xdJ46yhV0MWUSEfBvNVbZMFznfWQX/8sNxV+Qaf5iE7w/8/ptSP
XFD2E2VB9Ffr/Gp2yj3LgM/G+vaiQBwfQtaW0ShAtVqHvY/YWOYfLSwG2DcSNmtYo6IrYUfL5PfL
CKiw4u+NQUn95nTnjbFgGrIvSz71K/RcK7/9rcYO8P4EvXPqZgwqOAq/xKXCzAAiSfre/mppHgub
6Oq9phK2EMxYdwtmJZqSxrgisBQlxIZWmw2/0vBTbGJXqlV/KC69ByZgN3H5bTGVILRrAxSR0Hfv
2ZcD81sCc2PDkU/VO85MnMm4Ds+5JT4wJN+NbyDEBaCeSiW43A9wcmevGmabYmzm484l1x3MPwFT
ECihycN7qlSxvk/U6kKe1g1W/FGLE3f9f3zwTjcbW+gDcaVHUuwKS6ZSAqnWSjEMpfR0tNO576bT
RA4hK+lQf3JZXVWePR1FwnwzH1vaz85v+bm7MwawX633NxTPilleElDyuM/s0zWy8wm6DF9wDfE5
b5gQnWKseF9cmagfezIQlh/YoKxgXVH3B4MqTj7wE84SL3UlAtqks67lH7u1nmPgGi2gvNINtViL
BzDz/yoDYb4ERR3HG1P2Azw/IT/0Wdn/WicqKKKqD+93tr7dWZHPL6CsBFLY5GAsW2Jd11sZl0ql
bu7wsUZSwqR/CS4sxQ4imsbZ3MHBfEw22rv4nFL2mg6hIUlT5oCn4lsaPYOTQ5jJp5Sddepirpv+
vkaXKIOgxPuuLHR7Rnj7WR5ftR2lbaXWXTW7LWmuGmwcm5xiocBRAoPJ8uA7CCYT2dZuqYTsQhFU
FxahZb9shNhdI/2nx0s3WyfxyOzsk4KKOSJ8lhpPbwjQivYzLeM/kpXI0BTOAjnE7QxpFteHsfCi
lwjMvNSRAPFBscUTSi4pUYjxS6+/Nt3amqYqzTkYIDZ9lrEKS8IdA/cBkwBlZvPi0CUiuKNhzXBI
AH5g8On+yv1jHp83lYtfLJqi1vaud9jMXzw0RAxFy8CZG6DZXyiVk99wgFg6WCNRDfp9rr1vU4lK
qQONmSvn4e8fjoDNOFOe4MPjGRtlDLcT9MBV6HtUiEwavkbIcZPVm+IAmYzqqA+s1eZpaNKNwmVp
T8etfNZz8XFTnA6BDkGc40evjca501GyjFj/26vx1SCtWtizM3h/AchpcclsP0GckDorgRASVwge
KgPIC/UG9jdNaczcWRVFBIB6PymifaJydnBQ10oPUQ3QqNR3s3R6HDT+85w22gw2XR9gHLCwpVW2
Xc1B0Q6pYJcTpIjvD/OuzDlkVwOEZENldDyxQJTmS67UVHBdrgTNI2I6yIpeZQDtiM3UsbkClq5z
5jNgL7bxA47Puyk8YOMXf+GNg339oqS5Jm5HApvVSoKArzbH/T2TlW+Lo7J3TTn0GpbqfdvhsnO9
7FTRvOTuAhkDRafJhyJsQ7pzcHOytVg+O8NZtRu/OyzoaFSaKjbgO5cIfXWz78TgWGIdZ421mrPQ
HcAFo7evkBF+51tg01NF2+W62S/eHheMoh4seL8dgiJFkYfGOTQdWt8BBwrQ4CtRl0HrxzzuPSWZ
ZGeQxqaYTdqexJpMjVtIwY0EI8fHc94ITfYFRAaCy/kNgH6HA7qcqFKiC7ikOMZtSPwt1mCkFnhq
4K+fs8/B+x4nUEdrchbx08DhwhBMQnIxGT+9ixFydsU/U+FRRQpxxVpi13KtbYW3onwXREKI4ddf
7rJgMA24zkN7bk7zSv/3kg4Y+niXHDs/+eqfYeUsPOJ7GTfdRxBF/I9LB4JJ/R6n74OT8bzUhMDX
deN7r9r3f3mtHI7hke6uOvi/EKJuWpJGfNMXJbcMYArlxn3Gb7Kp84mkp8Mt5jkRdk3HLopPX/vn
ap7fzRjPPj6kRzenGOX8ZqsbYXnvCAOBsSo3su7WSNLN0VF7pdR/eR/2SEi76K49FzS4H2wp/01y
+wi2qje29zJa3sgFQq21KfD62lq6UoPCBnPnZybR/hmKVkZ0BL2KChZNP451HPCUYH5mHsRYy2pO
cNloostItJIQxKDLMxbQHwhcdkDpwoakerJsl2zsJbg4QypQMbLyRVa3vuYKeuU5QX4SCmaM3IVY
GXWMisNtop5LDlGviV7nQ3UKJhGVuveAMn2G5gyMjvOCAMAbVIOviZef1Qs/Iv2SWlUqOz9S+qJV
qTLZXdQ+b8fdsdaDYiseLebcpuy5gm9DeX0lV9HAZTmL0LFujK9F6eCVRC+tAmKK/hjZq6daT7OM
kA5aQ24qeF7v8sJ7k4iTdFTYOgbkH23KWloJy2WBKuo6zdWOURz1VOUbYPcjtZZmqwSuOl5ZndF1
M1cvf3i0MsjQCaDKpq4HedOrU0XtI+3TQ8cHt2Bq74WfhTAhu27YsfiuZEizlqqFcWsVuZFdxsRy
iz6Nuol66PPpFGYf438P0bTV4yQxWUICxSjfy4w5iZYgW2azDItn+ZuhPdNyfH1ObQ3rDZbMHqDf
uI/2NjvROe180dVuD9HqmJbVFNl6afrAi7mkFq0pXoLKh6O+peD+cwSkSYouyZDXoNxXQvLggBRH
siIVmA+owTVC27mK2QtBld58ffxnxPLWvmS3VvrmSI82VHPCuT9/3rSbHZX2VFDjc6r0HUIge8wO
U5pDmM4fVyCI5TPu4lLVkSeQZvQouqELuPs0vpRY15NR5TEBNRATFYgjvhvYgKQy1/kLQuQFvaTF
wULvJgOUhMTRLgYIXVQ/tj88RXOHr94CZ2mlYbYExgpH/Sy+Jz/H49mwLhuSG07aRlHUTPWf6d5O
czO8N30HfbE+dbTY9zEGsr3xo2/cX1el2j3LCvMSQeAMOOrC3zjV0JVgZTVUnoa7zHK+RmIzTQKY
B28ObGI/iKFJJEoBSncc/QMF+5OPDfYBri3V8lfLM/BIPkkd+yB+SfX9cZMVILWEFfi5abHDdqT8
zwLzfQmmGvuneGvhC38p0vokCME3nHktaxoK51JB9AvA8YJBK+K692F1lNUhKcI9fXOc5lqNEPy1
ndYrZ0dm4exAxyFyScJBgilxnGp6pnme/bCr2YCzwZCT4kon8GG6CMHMcGaxVXfkqzLOr+S5kl2X
VtwWeCoun19dFtlXrJJqiwt9QXDqDDE8USaoSuIX4v7RfD3kARzJXUHbmUj0kvt4sKVs2hDpHFkm
VfFgOaDT9/BlD6BFaghDhMM8gj7xq3zl36E5m1CPVpdbkZ3FK1jJE6ftlg/S1YQTrJhPkC9Ai3sT
BbkIfp32urHhDdO7R/PvmvXacjmJzjxVVJH29KpZ2SlmnNxJlZpbyr+NW+7Eb6GePgT57Sgldx4y
Pp7hjtiDFbALUz79SMDcbcVx5kClxB0DZ79ILn2SYICZOucuYbDkuLxq38Q4uHIDCrIYAc7HqZNf
yG4IC5suhdXruVac971hYx34S4Ga+fEz/LRzMRrMJ5So32fb05YZcTo7bZ0/me10VlQn9gXvsc7y
pGGPxNkB+m2BDBQVNWbGVMIlibBMkbB7n1sHfrjss5mg7kkq2LXELiTEF5Ahk3JRSwQvLxEFxRb2
/+irtHxxgl7v46yLdhUUj2exda/COOkrW/NU2/lfdNQRJ9dj7YDyddMoGjWX2P9u+A6v61oLtOc4
EJ6IJGaTnI+OYZt+mM6Ee9VX/RC64pqbJGSrL3cP9cAVg8Q7bXLfU8lcAh+9xoDW5Z3q7VykWsli
MRMz7+h7luerBQybwb9yW4OT7F+rvSXTVm5q5iCNKEfRShY8iSl5XNpjYTI3tJBaJol31dWeWsHP
FakqkmPCy/ed6T0F1AvWltty8lxdiKmscqMV7BOFbteRYu0qRAAZ0rH7QhPjuMJtf3AaxYgE40lj
qNcFkK5sTHKWLEDhXOI6uSMLACGA/YOM8rXwHaRZjOv9cgJ3xr1eCT8cD2LTcw4eH5E7PNhET8qC
4K8+FEteYlO40nBXgc1YLZt6kpnewePn85jp/WTshGhYNw9FQIJTr2J0qEA4mV6IRG2aROM4+slo
6tqVOtJDhm/AIrDqIZsJUyDrYL0MXcoJcqFJgYk45B0AAooOIa6dxqO/6Rir+snGQvkN6WmreWx7
yZnl26CgyucOvVCre9hoBAs7B1PbYw7Un+7mzlhqkMkLY4fMfhPgxZG2/z8EBBFsTfwfZHATr6Q6
roUkJEQUTo2wZUnlOVqED+pK4R+iOf0UBtQMalPhQ0u9lNjz2gk5cq+FuElzSQ6MBLUJd6Mjry3j
Huc3+5XKC1BLLxAd08lcKUMrVwDN8q8SCVlis9iwZD9RRlbl5+BDqYoSkVOSzfWGzoPGNrHHsytA
wCQRRLWoBkeoUma5IZ6nRIx89XtMfZMZc1tCq9/EiKaHRvrZYywgVqXHIuaK1bQDMSNHf9Wpa3Xz
km50CkSvp8DmwpllzMbA11mKYEhPstz0RRF8okhJEo85M96wmEwPjNI02aNqM5Cdy4cUtZXRGrm4
2xrN125D/eYbqaq71C16TkLQ7sdOfDLIu0r8I83Xr0tP8KCvQKechZ5wdrtbbcrbV2iMUbI8mDIE
S16IBs5Cjv+TfrvCGQUTlllAooGM8IEgG9obA7nCCvA8DDCBHEeqwLur2dGX+0YIN955eMLEKTtH
GUlCRp+qiCG8CxRaIv2qXp4Wss6SLV+lgGcURelCpKKYk4BD3ncrPxnrDv8FG4YN5ebtgjzg1dPB
24sV03JYItl+ffaxUVyJv3piC9wqZb+ZezV/7rJKw1N7tM8q/nqZBnTaxgjyvPdTx9Jwwio9RogD
VfYGSDwbZR2wEImpMXDaikL7a62J2M/gFtGdFnEIFf5mW42kf0i4MVGpNwJdo/nQEt2wOpDCK16P
s6jzCHtOUKezzoVd9ajpm/MlnoczQphLEdB5ev488VCSVAgJANXPQvCg5gPp9OCADhWSa++kydL6
ehNAW/7Q/nLn3RqpHwJX3GA8glvxJMWAdFm0ihPJwmM6DVJtOFx8X4DE7kwGBYJ9X82iCqWyAcXb
ytnIiBmlNyDb5xHJhbnK7isgr0W+BjDacwEDTq4pDNax35qmzvTDznTQt2flJ9NuTO0B86n+hBlT
ioiRTX4Hv79ciAOeErZzaiyHMKK9w6dxZIjyV8FXuVtjuvUFhb18pShnxSbwisdDliQOvUexqU+M
JGKuL36O2VJAP7kLDkyCLfnAqXb5pYhmbamatd1vCFVBZIGnA1GXtID4Iorp0jTOw6/1hWOIRMLk
xuAbr6jpyGK+Q6vOP6sOAxg7WVkqcXwVdgELGY2lPgxCq/+t8XNyyolmlLm7WFjzL9ADDv/dfCz1
qQVuEPPFtMQ4bPHRG32BDy8e5xWWgIqcvy/gkwXfTwiIHRfm2IUKrOZBDuVvL/1ysfUM/fRoTxra
jXRfGjNxRBE0G3T7mEX6LZz6X4iWZhtiWYvI7eBkXWzCnONNHasd1R0alry9emboLpnL9mlVCH0r
XXrMFVelWu7cfRZKJR1tNcQN7ionHE5cVCJElpiV8wBnH/497qzFUgOr1AJpIpHh9Ot7c+LEluc+
Fb8fipQ2L4UrKLrqZnysVP7ixsCWE3JLOMIYUOH/BiE2s6YU4pB7z88U7MrSyR4300R6ctVDKSjH
Kzv95Rrb+XRz8rODbqhWM/A/VMpf1pnywAPSSoKsAukLfUBi/GJJhcNOuPW1iivj6V5cRcVQG9Ti
cgHINuRGzWSIup78PdJ1SrfSERbqlGwPblpL23MnbCsn7LGgPGh9mCJM7Tzodzv+9E1oZLM+ETGZ
TzL71JAUeFQ8VD3L2ZGUJXefwcr2Ain2jXuPPB28MDftyrXBRF7Umew3UO+tua48eCYCL9SYvijS
hR3IfvYev/6ff4mqfio8lYmhbHonvzWohAhb5lqLY7+BVV++N6OSFJ/GJtlpDIIwSj9L5IywRNVX
JaRkGHOIr/qJowjnrFONLI0gG72LWXny0VPH/ZWqUqwYMVwbSL44HNK6BzHKY6ewa8KWYDgzegv7
1lhvs75xpif3CBE+K8jUkZdc92FW1eH1ezpiBTHyDafPQJW929XiPdpj/IvpMYfbzmKlfafqE8Wh
1/HLjpTGnE8jYbBisFGyzJ7vHD0MYe6NY9TiZgMzWfMfk+nfZ40LueOfFmn/gokQE5+/jBGnA/0T
y6g98pf/rq6PtkRxuTmGDgAmTZcREa2E0FDU76nhtlRhXKDQxrsZar7Yf/7foQrj6a6Cm8CGInQa
V6nQniMtlhoTr5TYDJO7KyB7dL56Mrt4am1Vc2mqUZAF/v5m3q+uzCBve9Ql9dT3Y7AzPtcE4ECz
5pbqgQGT9kEQ7Cy7NokuSM30PZV8iehjRxIBT76vCVHgYqLjkOtc866IsRPf3inIoNZnYQ1hCs1W
5M8HZrNxVGXqwucQHSJKurhURmRVVxTrRk0JSYVY3arUMgzydSpes6qfbiTYS/lBawiIW4xolz+Q
BmQJTeTAKYF0I6FR+4UyR5Nz5Tg4DXYWNFwrSdl2IaxCi56rZvgLZtJyXZnjoBocBTIO6KtUf2qP
RQmPujXlC7z3M2vd3LPypB9YSV8DilJ0+12vH/y6Tda77Lb9lP2/TDwgxoNqkCG3W7eD+UKtkeBP
xsZEtfUz6K0RfBKXbwDyMrdAndYmJri2kxxqfR1k9oqXr/3KA2AWMP66j6phq+hjrYFAkBrgTzuY
2n/iXfvWTG2kkfKeCERPKBm4tEGRZSLIsGlwuDDxDRF83i63LYVwUpLU1zpMoJL7fgBkHYBdmE+6
TnCtVZoMe6tZSwShHfbbA+jF+qJ+NQApHBeiXzncvodMSZBceLEJ+K4jB1uTaQ2YS7VbMn63wzZy
VwTaj5ucakOOjF3dl2NzfHLdIBzUApzxvX2etfgajxeO8RGcV6J3dU28tnT3NfpF1u++nTUgDm8t
BQ6/pW1NUxhWaC9BGo++8ZBgay7QYzBSG7tYgag4c6PaskCYkQvq0+BG1JjBOqwLwNvlyRKB2chl
yCLLFrkOmbpq0s5+3HOMcIfrBtIRnLnUSl0KYII0DCCGrD4FU2nZnFQkvk8j83ArOI+rcWXNPaCk
oFT/z7ZpKLUJw6ltyfoffW53yF3BtSNnUQamXSc56oBc3FMINBIfsd0cSMNBcGBqTS0vC28G48v2
BLlDvaY9I0MZaQ8CKJv917J3mWr3HsF3/d7Wv/bvnCTLk8e1ZUEscEY+kRKVRAF1RpITI8+7bPiH
9bTYptKeARO0Yq9WbrCQm8jnuiXz9VUf7D4ZHTluKpGOAxFwuJNcPPdjObt5VESM7IbPdRorFXmP
iBGIiAjRKVMihXvhnSgBQMqJek7cuTg5wuJblLt/EbPcnxPz6Pus0uNAjH5xzrYYJSyYYWv8g1jm
kWmFdnPFn+WcXh3r3ael6/9ZYGMEFM0cKd8jOfM3CYUmvjLOOD+e0tK3gvLEkqlM+nAtyaD8DVlw
221ElrfTokBL4Az327loms4qD6yXHKXj1MKDrS1NlkkPX8umZqRNr3qpbudWFw2BFEipfQm4w5Tt
6XMnBxT/1Ei/4XJYy6lxDdkv4o+ehslUN3S1gkzLtBC3GxxLkNpU9rl52d6TWjN8d8WW2mu/7iTJ
v8i9TEk6YH8L2usq+PaYSGCDVd21x/GWhUOCUooy3/z5Pwc7uKp3aQ5XHK9BVzDjbNHf/z8Tk5in
UF+LGS0j/N21pfS+9yrro5CaS8HshWQLyJuvbMyJfZN2pzJLa6gh9+GB0wJR2nfZlFp0TT+ZIUc1
Pf+MCcSqe+nSpNJR8xxZ1q+vhYdFbuyquqig4OqUeA638y+9JEg3R5zlJyDGUYbuGPkJkrjWnbM/
LuzdG4ynV6vLUSxWFCY+8vOljXAW+Fjtiu2+eRD6KmgEonvZ4jXaLlFxrMarC/Q1/wgb69nDdXOS
AuzdMsov3Dz2NeH3e31jXxN1fxRFNx8XqgYer/fTKP0k0uqgSx0c6LDb3GuHTVgjcYxltpINBPzT
Iv9KEEnKA2cYnO/bzzkV7C6JQY4vjyUz+rkEVIAbKs0C4mIIdOoiwzwCxZ18785a0trns7G1JXbD
wC+BBnVR6NUBc8uRSKcpKuwqejGSj5AaYf+eyUEkFIxmGuJ9y+J3j2t7q1XItFN/Hff+5DLy7s1b
42NaV41JtJq/4aoYjyaidel0Vxs1ykTPfmMadtQvyJvJbeLgtrx1TjSzFHR20tvIMYUDqVqWn1uE
u3OY8P4+Xuw8lwsVYeft5y6l1seqAE/gWFIk0kewiwHZpPTe5Ex9zpetj7JciLb2Eel2/Dyb7u2P
1vmiZ9TtOI/j7jPxaE3xDBfziLl6vBD+nkTKG/6EJJZ4KcGHjdNi/TTR6suYYkOFaGLa5nHHjUps
YBUVRX8ULOFltb6pxmLdXVW6iqyDD3zlMvurZ/HPpVcP18jL/Sk8NaplH6dBOD8JppdDwm1Ye7rj
/59274d+78m8YoDb0l8QgxcPv/zK24tLG1cLw1MHirEZtUibDLvrMCeMIU2Ufb/OyfrszkSvmBNN
3dT5gwwrFm1Tv0kS9qme2xDChUHnE72bcKOQCUPTrGqeg/NH1xtza6QYHBqN9QedIFk4lJu1FbY1
qHJvlIGE7UjsiuC8sugMLD18ruKhAM4moI1ph8ZZpkHNTJFiNItS1ya3D8CwlaVDjLoJmXBpcjah
/IvdhV7NIwpk6xNN+AT1f3X/pPUatBL7prff6MhlTlFbIRWz73eII7J3Ou0xgK0WtzH9kyMVIEL1
VVKk0RZHFZ6JdZbjZDErA0puTHNsSNdh8CpBZ66X7rPeex98m9YDll1iM0s+MmajQ0xgxuKXvTyw
qj6+O72NbrtiLrZu0BEdPHRz6SUwycBf3EpFhFT70ad1jbNdx2LT5qAxIunDrKGFVzfmL5Nb5SAV
HoQt9NTjFByepms3/LTTRcpr4W1zkfl32GgOebTkAoANvtokQNoGC0pGl41SNHs1AgLDeZJfte1p
FGzvkbnGHGueD6lSE2hMwJ4VUgTDJXnz4PEjfjzNOWDzIsEq7YSO2e0DytrN2ZdmA5OGGqdKJ8GE
jq5mx3MmIvTlOPKkihuyADZMSl+VLv3K7M2jbOfj8c8+Smfy0laQw0QuNgWC0zu0xdPiSLxoha5s
kUTw9ZRdKENyd9qoNlXGL6eHFFayp1KKo07mWukiGE4JfQq4CQGHvkP02FhRW3jTZidExNUIui4s
o1B2KHhT/pyRPzXvuaYNKcn9A88LN0yuGepxiVLrKeekJExjzlnwDl1jJkXfMN0uLCO5pVtcen0y
2gGLR0BpGuqgRh+orpIZeKHqcBaRLBiMcdSC8aqoyx3RNJ0ssYQBRPGgxRLStIOqyr8OCQxwmay1
Su09XZPwLb8wtr/sLEmyajoro9BgF6LoMyO6OnCtfocq+2fk0+NQ5616aPsNqWSttEpjDrcsTpvW
ATm3bi/8OKr/1S5LcuofYTnKSVlmnAL7njDrFAfFWHJqQ5WjbGHwYkrZogDTPaPYXk23hIXvsq1d
JFWiwKLUgRLmn5nWjRfzi+9zE3RbgAj2JSbuYflZtfY0GB1hwskwgUPeY97foNcTxoR/silUwVjs
KH5eSJnFlrV8flQ0dpGHu2OOla8jDPrKJkkNBBYU5PLSWArKaRanbXw7YA7xHneKDSMD/yMSkeP/
QM8HpyiR1NeKJeC+CfS3expF7BuoeskUglee0RF6ZJGhkNGphZyi+kD7+EmYRtpfKSTdUX8zIG9p
4VPvT/Ehk03jHCrImXZdP9nQEASkdKFfyK+Vk5qpLWZducpcwM1EYCToALrSWwgU1EIXD+TnFu62
jPMJ4UdbZZnmt5BoNTvOFSVB7ZflT2ec5842rtxg4EBkiN38j0tvu7Rd1MXE7w6WPgflr4saOiBy
GigNbe7fCLvyKb7IZLAGyhIVDYuF9NOQ4Y5SctA+U3fjw5rI0aG9u7pGAVAVqDGYxypJJNGuR4Of
+9dwpdJoN5q8EVt74D8b3OFwp1ZhVTA1h1axCclhfmBdmiP6G44YqT8A//eomdUy2hvLK2jAwJ67
Ph5SGi69+Y0wNonzstXiJJG+1mvC9FTuXxoLMfbsju/FYu5vVCGJA2+A9RBnOdhYiFdp4FDz80Gj
K6o1pX1pVaHQV0VBljYH8evT8eFqqop2HOIesY375Typ/0URziY1+kj5URjv9f5i8cYUi+nihGs2
msNk89syyGM9o0dhWpdLTr9bDv3iLQOb7wovnhQ26d99ZpzVLALCpjI0w9DjohhHNvDOlpouapeD
LtvYIGwD0gdJbOptge2mCYltdy4H4o5yzHyseL8/ErWcoXPieTRa/3i7EOkwnPy11pSqQwsxc4Eq
XjBRAj0VHcEGq1uURBWvlby9iua+njUoQNlhpLPfxIVqoFFn3m5LdDB2p+DdBRVKJnPgnKfZhbC+
QXceFHQiybgzMs06rZXCmQ5aZ/7rhFrT14xUU6fI8S+7MfSVRh2nqTQYwbjoBlEysjhonZorjA4O
ExbTomBMtRtErvNCH/CBie7IYxSxBJ2hEZEyhaC+7coJFzfslw2CebdPPPVaRQWR+F4GYzWJTxhs
fudf/tdTiRzY+t8g4/rn0aYWlQni9TSr048dB4hsnWI9/b4CTPEq039Ge/Vc2sGaZH1eD0t4I3Lr
cuhPT26/RQasjuJfJZsAQM98WbcHQkyUJz5AtHoAUEAqHWHJTNFrvzZixENBzTzbOEzTswWmZZH+
G9lM+ibp2AmkyZpd8kaHfQ2iXZbcNk4rrL4AI3d9XFcMWewxoLqDd9recFfzS1xEHpcSv32NqeQB
ijK7SozXSKT+4wXTxqWqhYvRW0AHtB/vEUSrG4Zmz3o89yQ65OEsDrQOJWe5mNwzhjCm45PyRaRr
jUh/Ck+dEk4GWDKCcJAJaqT0APf5V+Pec5+f2U7odk0GF1LmZ6uBJuysaHM6BS8B3/axj8ZvO+7D
+zDzZGCeV9tTjSWtnTk1frV69XEN/KYIyLWS8DA6WZm4UFYk5t3PvD5nflAZarcUDT9SOA5Vpbmf
TzhQmoU8ow818jlBPzObpy99CdGunLf0RyVgASaJXnSHMzNXuc9Hs9Qdm+jKjF2ZBGgr8tO/3X6R
hgbA4NvrZSUunrBv2DD4D+XuVsGZhMTanPt2s6z0ZBMlaLLQHjED9V8fVhWB+bnevJen4EVXHs1o
DfwIQKLURVH+/MMx33zZ0j/Uzu8vi1yEj2P9BsOyH0bPwUxWViJCFBLFWYi+aNVLGFFWKOSfRhL1
s/vixPFZRSKB80RzFqOT3KrwKg8EedHEpxoxThgfLVNwZ6N3Fccz5+kVCevTPHXhw0CDvH3ytJ8k
qa7SYPcyxkk1ZUCQhFRRu0j+eNsKRq9UmQFZajeMvUpKC6bAWLbqYqurvO89dQ4JSIM6+sl+SANX
12gB27ADTz62YqQU57CoeR9etF2d3mYTrAakiZhqfCYz5HqWYYQMoLLjB+P7a/xOP4gceUUmGphk
rc6XtDHXF3lfyOFIxpYvtyFK0nL8oxBg8QHE90+LVNcqSFC8llSPMTtRY0MOPoV/BjGRWLLigIc+
mpocx47uy5OGsOVxpKXKMPpEiBt64KLwPut8AqhQ2pxwkHQ74dsI696Pgj2HwMLOOJbXDRrgXanR
zrqK4FIaSi+VlC+gW3KwxA1Li8q3eA1vuBR3kW30HQ3pMTyaKoAlKtltsR459UYuut/7ri8iqiTJ
L39gmUvTfa+EY2tAk7sn8/4AQpQC7sXcC8IHoCH4y5ovXNkBMfGONRDfxeFVtDCA5AT2vttxGNqp
gMXg6thRrW4vy8aa1Q6Km6VOmQOfEYmZrzYmMKu5Tga0ZcwF0JFi9pjVk0p4mGPCYWJsSPantEpR
myi8D/XvfcqXJGEqkj4426wVaVTLsBiuZ7qjZBst/fPFRmd18JDGJMfhdnbi9c0ztqA8LVgEzdXN
lfka78MVYGDc5suw4bwzv24rucsk3goJ/3Dg8TQepYfDA83VbSu9av8aFfNXfFQgOnyMANDHt0zJ
N56E/bLtEAU0QdkKS2xU3ggp4bG5o1AUM/5CXYckhz8RojpMUXXslSDADkGqrQVKcagODA4Uucq4
pfisClKGLbakPRvra8iEe6uK0Ujm1rU/+wRyV9PBHmdA/3VxYwohVrU1mfKK3El5NdNvJ4d/cT75
dsWJqI6piM4ltLWcmCZcq2urRC1g48wW60O4mNMyX1ZHhplyTKICDe9dH7f6TK3KFLW9apsEYci6
F24L02T8ymeaLqjvNFUYwRN0XnJcH8b95MJkkH80TllihlLZ59kzJoz2Z0WjQ7Tm/KyEJ37jUhVZ
+fJhV5fyMxxK79OJDrjyEsr5kAKhD6pytvRfq5QUvjfybuGEzpNIlexhe7XMFK7mqy15+gYke/Ev
SA1//L1FyJRe5aI1oTQ7f6OQVN0g3JZMy0Q217ArvbcUDuOe32fgDRUm+CBXmsEb1NcDTWfcZ82U
tNk/I/91LjYK8qgEOGUBkCzfFeFZ4W2owY60wBk912TZo3ojJmvA8MPlSBeRTc1bPyWu4tweITOi
f0c22RmfAbYOSpvDcUrwn8kUTFaqURQ+D0kQ+v1rQ6yQNY8Nm385bX4OKze5OpGzlDLKc0OIDLci
2T928L4PadzM/zf8p0L1wjj+xW83yJmGt+sr32WTsV43ov+dgHsO/pRwCOFedfgzBtyjj2N1FADL
TWOfLq2P8Me/h8U+duxxe0kgtJA5cuYli/ibPuwyFVEj0SZD7kFcjeqs0Oz8Z6SIJZ+W1mqK0voO
4aTnOhj53RoLxhxn4jAxEWWWlI9bwNIX/20MjGc9ZuhvsTM6sljSVBZ+BJfxI81ycUlLKuOBx0wy
DvBAbW5uR/CrVDvLAsL5tpfGcfn/wSBHJLzdp2PZum5iiT89glUCIZ6E8Lb5gKb4EgK+/WfoKb9a
ZaGdZapd3cX4xhUzUyiqdxfdYJKfGWtf0C94ZWUoBj9/M/IQQ3zdsFzOF3SoMN4QnbG+LA43bhIG
Gp2BDfH6tDK/Tt8Uun6N8SEqUkFNeIJDfoY/EJIBxVt8irAQ14Pf8lPDj+N3cQZD2c7m7hGScIgT
BK4ZH8zFomg+ZkaWDN3venxkX3YmU3HDrGLNCN1h2m8mdRi5nmL4OetahVkL1PgZnHOBO2vaErIA
hgvsr/fMsXXkfgPNgcMeS2N9teCJnZY2kiTp8MRjQS0dyZe3Me+YUrZA6F5rDOiD9gEVZgZA04e2
eWerAPwZVNpVSO4IDjOlN4kXHwx7X8urjS3y2sAZckmeg12VcQioXIJpmOrgoAzz3zLu/Nt3mqzS
OaA/tNslk6grwEHID7nHj2hL3DvJbNmSEMQJr2CManYxFK2Qd9NwQcwZYuhoO57RbJzUXQHzVLTf
EaRVBlYv9WtE0yrezp8MAej/JUsuJRWYgf4wRzPkNC+c9ININCgB8E8Z0W+/LAzO/ivJ3AbXaBLg
lcy9dE1cD37Fhu3QmJKxlboK9mhY++LVoGcIzGEzIRAUy2Bzyp0RrQFlzr5Bnbjiz22xRJQ3B5+R
SHKVICQPnP6GHYS3yBlXoPHpi5MwUriP2KMF9Pxim/7WaQqSm2VbVpsOFgQ10wSuHvs9KqzmAdEH
eZxH2N+AykuRHqZO+yykkJzs0TMViEYjyePHONfsNv61qMScILKX4k/STbhcZhtOURC/WOuwDLRZ
4lmy7rMVe20JOTPRuUcpWIiggR0Z+i5eGmQVfQmeYgX8YqG4sVaN8Dl8JNKNBhgPv1o5izmCZXYb
y+YhSXz2L1sb4RcYKJ4YiU5+9MPlzkuwN+4uTn39YJKGniN6kTrv4Z0pwdqAfmFgyE5ZmUAHee1B
S/v9ug2O//hLYtJUdvcwKY3eifislivucu4PcZcWXRSrdofw82cZe5wnK8cVJFQx38hy6Zo+rDNN
Fqa3lE1UyGP9ZL+W6KQ8/rlAbNDrxEvOHGV4oB95tLk10Tq25DE2k95cuu910coZUxrDQY2AC5nj
lrslAQOdDqJz5shGTvBBPzvBJRIsNIja/Rcc/pfd6wnqkVEWMCDdSCkiHY/DM4qE4eAn+M5XRNub
zdlUgRTzm5oIPMJwI2QCnwL0tdXp+7NGlLOU1s1ezIAMNFHsXkWFREUZWxIIoT1WqL3OC6cZBPwl
yfodXTQXRI9dKI3I6B0mRrPDfbbEC9bBpf9I0WnmVowbBHv7zdRNZlDo/DFu6BIwQHRqaUFOCnMO
ytMDrZTDa4bdoYIhMm/AEVdpBCS9NfdWMiKSPIdWcVRaANt49dN6lUsQvzhyZSQrJTg8sjXuWrHE
DirVqJWDz47uNO74IbnyEgvshijg5N/vGVBZXbwKbnT+ySwU/fM7mADdItMDKqk//sMIpRH7SkUN
1EjeAwEGUjAFEgr8aXFMSIF0Q8WQKbdDFB3Buo9o4wXlMoCLXoOUQhd7QG2YXWKGV1PgWXCY+UTw
/guenFeoso4ytKJk4WsHb8dUlRcg14488PMRk6Gebqvn8LxJDPDTqSt1nc/Rb0zbo87oSYKLkIHr
SJdrtlUGwvVKKjyyBNjwE5bxtRPVXSXISzjGmp7TURysYHm02u78joSZfeuBH4TFJ4UyibYwOnul
F/qKy8MJkFR2/ixzBvN0qSp815Kd4rPbF8OFqd0HBuuPTvQQqHcAgyYHFmzV+WkQZM3kbvfOGKcL
soXzeVE78eUlvqGRzvuv/jkuGosNY3G9thoiR8UU0YNo9DoRwflxjWZXQQSCB4wHxmJaYa+/RgJR
0yK1b2MO3bku9MnvnKEgFMayArfNsMaU+a/LfVaJZQpDF3hcS/H63Oh5+y+5dr3L0DdsOImOoFYX
RjGciotksRzOTJvQkSga9ZIzsXsPvjJuInwywl3VB91aTOhTZCr8SfoMllGQN5yuoGcpx4S6C3Ty
Av9yfsejuEiYyAHLoG5N77FVLUzEnHVgJMTCKEOvWUesVYyMaIkilop+w2RuyknQaRsSa3gE1SjY
Zjb80SFuOd8zUBEh5h7188LcPW62nbDmJdRUJMCWIu9aJMPPw8FTYD5IjuCjoh7nkrrhSYaI6eI+
hnCNOWRQqn17v/WSOkPhgT6PIOxzujIMaVPvffpkwLzsa+jmnFF/2I5MwL1R+aZzSzvz8CBxhuCk
F8USWM56b/VnZ5GlCzKhUJv9pT8BAvG3E5qZq9Fx06rNUAsKK9/KGM3V4E/+gmURwDZR4ajWLH2C
NZ0oaZaMMNwuUGmtNll+sEjNTGfFaijOWVJDmty8UUcTs4EC/E2MVOWghoew3NSQncTih0eOHQrQ
PBBbdRLyhDEoNTX7QF/pjqRB0LEARmUpa3179Miu4osYfEvbioG/tmHAma4J/gwDeG306CT1ILyr
enhWsO9b5FhMu3fYSGz/hvQEDmJB9cdodcNT6lxukWdl5LgVBXcZZKpB+DnEXC3PA68dSeA6Iqx6
jb4vvz2uRhwQGeSlnWOaJtlwaQFbxS1qb52agvlnn2wMc/+f1XLvTyFduphNMNxSS8NRRhHotdPy
QhGdE455Hma4eUCwO7IE5axWZeks65t08mrHSTUx0Vmb3tPCbXZ2zRtUuUztfpdATeMSnAgfwY/A
Whfch33C78Nl7yfFggrmJAA6vPVQvhwf3B2vdrRw0/yQxctFVrLPtySk/+SPgPRv4f2qSF5UpZ6B
fcFiDq1FwWtswkKU7n33Ar92eDJvS+nIWt7KzEx44qw7G1o0q7sx6dhZedQfUZskVNKFylMXn59V
ZZv23eG3hNkxo2xLyJPwqPYNvqhbWY3MPRECRov35fNnPWrkPdMuR3DHENz2DP2KhFCWCk7S2zOi
wyDCA+ExaXEYw29nfNDn7KXfYPV1hiGDdejYf69Hm9/1okUwa3pIWKfovayiwNAEFC6MSl6xITUx
llpRtEz69UBqlzgDpmVKh4AbCPDUul9k8Y4BYeJEo+fwRx9ARmAqeRWnSMe2UvjK8SJUIlFPJMCX
2XTNyRnrGTOtqd7a1wocDHIGg/1s6jJoK3h6e82sB/Ol4nhNE30v0yuptYkE/NvGRyrQVXNq6I10
wjxIghvoyeBXBBgY5TkRVXL3fFwOBwyaxSIVJwMXrHwZsxNAc5d8nXUkxUpyoMCZODEn8SXSGP01
7YhTowlaCd04S+6d4ErXSo+f9jqhU0sG3SnWXbjULWTVIsUd5pmS9DY22INuRWHnzpNL6vlh6VNa
HN1Pi3+4LC5iELbJgaOhhrzPK+EXpMnqVPdmh+01US06iyohuRYy4r907qtZ8h4UFfqLP2QIuwXr
MRtbw2ZTByFA/fJyYUYPYvmScEpFTxyaPMnTRfCOtHMq+u8/w87HO1x6SMgkDGuSOOJ/yCBGPjVf
w1z5szfCHrCPyRCKq3yah08/5dOWj0iaskDxuvu2Agzljld+HvrijSg13JLUcwx7uEvjdktwcHCy
Sj/wNaRH4vUbkbrdHMoPEFvFMAc8KDy/ObnF5rkauzYSOgE0+rWgBqDmUcqVOVptSjh+sfgfbjiQ
qm9EqfuyfxYA+FXzmu/6wf/Pmdex0ud2Q6nHntB1hTJwwvv4AqxCI5/WZf8WKOjs8JWPZ0UqNZnk
E39HOlcUtVQ41InFjVpDSwH9UhxcGeafWxKM+kM9cURbwG70921WydFdM1w2eJhJgXRs/NMMxyGP
Sq9jdArMB+F8iiKjmhXjtEU06Ir6ZEUxxc8mMmMdmAq+b3fqkO3BJmiklSFe4gMj2AO4RV5B8EYn
LbMN3syNndvpbfcWRSf9pw/xrtN1woboWLkQ1Biwnaz1AsI2RmZKL30/cQO+5RRHziMZhtnn1x53
H/TmLBVZmENSkCY6a5t+ywX6HkOoZgecefpoLrFuN61sSdfwOEu+onvWGC9udaV3br0K5eOrVPE9
+E7yo2nDx1RctFHR+bDrbrS22wsBG7DlUepCugKaCM5Pze8q5zxXINyH449T7dEEsvfjE9jdAg0m
+zvhiVe1V1jbP+CzWv7Gtki9UgsthJyNbjpeN4BHIkIltKeSzPpFBUq2sDVY0i8STk2UPUZWX7wk
OEliNiUGt/K4f1jkt+6DP/+L18GXt8yEH5DS1M0xs8rc01xQAU+SGZ8/dySvR/FhqaMfbKrSV4xB
OJ7uBqghQEu1hQ70/Drx4jQBS5qQGsoYw77c42WvZVCNRrwwuhqYO/ehI68Y/QPeM9XjVP4fZum0
J+OhAJyv6+tvaIbb97OKepAaA2QjGkxTLfUDZqJ3I/XoK8spLdBqlVJDtoRTtvxy7UduuXw7/Hub
hEfD6709vZVoNJb06MWUH98fabNTY7GHh03/dphmALLYsLNDhISwUxp6SWL4fcqr7B541qcU3tj4
X3qgmseI+wuL52FUE4QSr8N3y77/9Bmg+fv+EB87fQpEimVvMM543bfoTdHidbxGnNWq5Ldfvrgl
+7Y54a4O961qqlmmH738wusW5R8ifB/E7oO/3DC1GRahNadgz9TKs5EQ+cqTtrK5IF2NutJy+sU5
S/LymzVN4m4dB8YrR1etnsMPMFvg4nXpvuJCvuiDn6MKmFwSFkWaWgefCfGBkyz/CLW0rcVoM9KY
qHK1f7x0tf4Q0gm158Zkgi4HijIRaHTAnl2EoQG0NiUY/j4UO5sWjF/4VSFhQlxA/ASYDmr+TwSy
SMpvBTF/Fka+UAvj6IleRiH7I7Wf5s5a2u70sfwtVyfrLtBgmC641JpaPgbKHUnT42zUWq3+3z0D
CdSvDbV6Vhgbkxu3su6AELnP7Q4cFjFkH1rbjJ7GAfVto+omjPmfnGIxB+dHPCiwz3AdLplP8Gzv
XZJBbj9cjJlCORQGrVLoeZXc1Wwz1CwNLi41kEZPbbxj062BTH89sY/qpYM2EhPnidflqgThDN8j
HTTUr3bYBQME/2M176A3Y3+QaCBth8nx0Etu2DHD3DjbEbCrhMkKFL1w0FQ3t0iB09MZkfyFZPRf
uPSy5AxEdJSoGKjPlO2qVcCU+xEUNe5YVv85JSPcRj1Qj7Gt0IHfCV14nXXBj4N8Soo5HQ/j4ZdU
OqKjHfuPFX7yFN3/jBjg89DIYUCAKGviou/C0r1zNPTxN+UownpsJw430NRBl0V3knn9gqQjFikS
55QMRzhRUkzlDjKPwcAk+gFYmhUxp80Orycjc+5pFAvQhquGGyFds86oxgp9tmX+t0NwUPp9w/f9
71sKee6d/ET9GhC/9+zvQnnCAZzJ50e9vXHWDuMxr2Gnw3p/2TG8dzKK4RS/JnZWLwocq3MsaOXZ
zYWrDO2tUIIFRdHNlD37wLTdXYvEo1s/Zdt5oT9iKqpukWDbQdYLapE5RsAuIs2AvEXIxAYjOM1O
7e2DnVd80XWrzuJBI2U2lfrQqHYzfqpmuz6wQ/BVka93/hznU+rteey0+rVyCVkE1NTPwJuc1LFD
4UEbJtLN4BICYbQJzwj1HZq3ll7haBnm+aFNigUNJKJpMZUcQNuEwFz/ekTnkVmGki8xHGh6esgl
fI/s1wgyqh9r/4nHGtlN367FN8980vKlZv2GmI6ArZAN5t5L9fmCAOPEtK7NLG0JmxFy7E9gaaEe
0dhbr/+pl61IDfQikp80tt3quut/ukP8tG4UTadp3FvPXpHMrFMzGt/Fk4/zyuBflqTH19495eRn
wNxgw8R4DKnzFI3x25+/dh7m2YQEwXFKh+8bZrGiu2yeX+VE2dwwD6FRdesQdmLlcMQndobFsQJC
AGRJQmX9awIKKqK6kB95dVeIysUNgyoYLRPn1kTMqSt199/ntEDLHwZYWXEvJLDI72aMhU33JFyZ
ByPQWNSb03CtdfKwy9iTptEktJYnrooqHS8XhxtNXHkFFogxhw0EL2y57PI8eZQ/6j9UMWNAm6Ye
IiI/wVjWCbC6rr62/b3yPH+Oc3xlJZBEfoAIQCBkNzoHlpSdEXLvgsPy/MAG8yUQcsdFKMYxFxDn
+DfElxFuqIIQfDTvd0XZiqV9dVgjiNsrY0DsI9TulaAZa72ual4CqT5g6Ul/Vzwl5RnrAgL+UzK6
O+JJoD4ZM9cHKUB3tKbLwf7diFNytOUdwBnoxKKsDEkMUKHXVmzwI/17+K77rYG3N1OPW9tJBc0Y
h+1Jyq9BloEDLLOinVRmHZItxWFs+Q/J7/XCK1PiPxEry8UvYhhT+sv6xK6oFtSzp50EchKY6iAt
jvyjGjJ4oXz4BGPWDXgzQ4WlzurvNyPdvTWy4ED1U41je6TguEFMcGsyozhuTYwqGI8xIQRtzjSR
LZDn8HzfrZ9GJERDCPTnqTDqvqEE6RejfDi5FezQXtH6GjCktQDz6azE6YPxkh5XWXVOywLdSLA8
Bhgq6n9mYCOqHIwtO8r7nZwiuvWTg4zXXNuISs2KilLEnGIYgviPnx+yMp7XuleCh3Fc/4YoRVeX
uwul+rlq8ZtgLpWtROWMERvr+SIhWhlH26TRAl9j5u3byxPYiZWsB7LR5HNPbKj6pH/B8ItdboBp
ZLcgXfaERVBM/H2SxjCA7pdxlJW922T3bEw6K/hBPJCTHOAJtPl3Ge9lKAUURmI6QfZWUoCcHNuh
FEXfV5SDuJcSrEf/5yFOZ1X5RpEspQ7X40H8nx1kBdiOBRmY5QtS6QvXk4GtKoPECshMYnhK8YTe
v5yyCEzX5jCy9kBTfgoCYCLrmsPi7+E6Jgo3iRG55W0kDsmpto1+RG4C468o4oLzWnPPrVrm8phL
kd4nWIt3kFOmfmgNq7ff6VonHOo63MrvtECNVNFe32HnhK+cO2siwwt/+84a69F8lBfv2+kanGAZ
UqMsshxASa7mpN/9oZrVpy/CRJzygzHSbUwcpKhuuj37zWAFxyF90713E3ArlA9TjgPtG5dqtk8T
I9wTgIzOsu9xXxFiAHGAx3bJkQgRIpb/QJZlzdsb1LElOCsp2lJZB759lSQkYOJzO8IMEQHFtKcs
eUbzmbJWVnrwg2dBklyWW2nRfM1v+mv5gAlMbWopaKaB8SJ+sFGxdjpDW5gSToNubGsRKGwess7v
e2ulTE4NWnQmGO7+6rnoQCmSZtQ1QnKeZVJPy7oJH5a+268E+d+eZYXi8rdcsqbobAq3QxSMQQ7I
Fp0qsaS9JlPw+rN147X+jEaqnLJrg5I7p++9Fv/jokcmiKcMcVnN5Fx0nxy82Ukkpt/tUY7RiXBr
rDGRCU4qR2cHFQrFwt3jNgyC5k8llKQQN2fAwtMvsVcL0D8rQXkFyJMySWi04JEhyBkwDxHNjhpn
hFEQDkkOl2xM+ZNURkGeYKMGfAKJ1xEtt4H9UxgiCojjndanPHz9ZqcO6jpp/DgrZGqoRrvdtNc/
EvT6/fB/xQW5ihYbYSvZIUGrTNeCvdX4z6wjJ+YNpWFlO8kBd7e4rNRNywWKQUlNfUZUQwoTmLxd
BOce0WuR2p0VVDuammjNrCmyxn94LlYnR9YYgaTeYu1xxtQiqnbUu2R125oLoWEq/dNUMgpHnihQ
Cth4teo1MDOJ8Ac78FK/VYlnviEXKdvOw3yQuIMvON0snoz0iXdhNc4ThXKubPzGSpJq2LU0i/Lh
lq9eg9c4BdNAu+P16Lg1oH4F6ZJ4iXFrc8hEeDWiMtn7gfFKlRMm1Xkn14QEYe/v2Su76APGalxA
Xo+zsVYUtB9gRhL3ozY/bnw5ShMfEyQv+uvcqpbBwdMB0yhbALvlpox1bvgJ9zj8NGYz1N5u+40D
TY1NX6D1bYjxz+DGcWIxwcWFs6CWr7ZE2OIh2dHGPTB+ko9geVx2dwHV/XVuahxeURZzAjq6IpYe
OvgMcK60orlnjMSKTfjIskbNTf7nUTnBpdFr2V3bXcIIZj6wU+F7sXkpBM0boGsb9FVRumc31oc1
ODgKr78xa039WRyTCz6IYoSIskozrdIzT4kQO1IsE4IcgKgk34MfCHhyVVxRY1h6I5vIiO/veB2s
8A7xEqlOww9xum/8nUefBXDbfJdmqt+Rhv2KCxyFGBlG5sDIhpjUIVrnsGC9hIiMYWMpSsihxgxY
MQXkWr7ajzgXunA2JFgSdyrCS6TZkUsY8lAmFI5koDdsSpN5QIWueRsZVdsl21QF8DluLdT0s8Yn
2Eon+nla/g27+S0OAAYf1TrF+glpGQXvlUxq7v/EjJABxJ4MtjcD8uNYdA+2d34RlTqMUiazXvk+
I1gyI2Dha9ZS1CLGC56+NFDHERqWH1AdmJSvHFHitAUZDRGVjb8H9ZEmI3E2sxQdty14oFhfswez
2ze62BZIeEJE3VXhzAiQ9FMrVmvrIBZOWYBGD3UHqawsLSxW8Y/kYuNZM8KVCx2tP9Qz9jwtT0iJ
OM1jeK6Gx/BfrGzlgphrgkQh4vFimdPQW91f/eo6eywKfPnf4nV6bPMEIY1WBynhy3b51roaGCkL
2acRrU0ujli08soa8z/+ToYzgsBGZLGL4viKlfHp5duUgp+S/i6zC2C+iLEL6iUjCyerdHuFdpU5
M4DBSlG+MZgk/pp8j2BHc36jP1SSm8sZTKx6WW8KEyJGtdDGJ231UWx2ZrovB71goA4A1iztqoRh
F8fWD7n2Jh1aHjQyIwqw59LWf/fiLzQbh1J3fUm0BmN4WJFHxP+VXBBjZ0Idqyx++dvs8Sk5B0wu
hm79ipCUYt215YhceSMgYKw2WMXU0r6n6k5VWTtTXddzQlCddkdWAZZE4nfrMVKZ41GWRJKepNTL
uO568g7c7VoYe5FXZAOwvKD1qZtmY/geXWVlF1p7Ehm5tjbuLLPEfVjHTlKhZ1SVXZrxQvinEgSX
ySxooUym+oCVYvejG6XfbkvBsQjLpZGK9TdYaBXbDLlFtn5Z7g3RPJ/pVL3TItQaLw/TUjVrsQEk
MNEQI51ufJAcWxSTwFNH8/4KUQUJWad95sz45MTt0QVx12MMJsXzzylHV9JrzIn4RzQ22EcFvDWf
sPOYK4hJrFYsm61A6FtQR/4mKqO0rmeciuFKad7MiEYrDPHQUnUWhm4IfMF+Cd4OqPaIQ1PQlNL0
m34ZinZ73VANo7/oJ1EfBO8gz6fXwVoGxOdhGPqC0LjWAkl0LMfZueKa9xCByo7kn1Ye6qT99h+9
D17uSo4sb7ABPOolKFEVsFTlNIzz3B8/UxQDaJ+Fx24qtJt3mtqsvLmKg+GzuYSErORCPb+ICHq/
OcVhlMugDYetWGb/uILR9j2dFQ3XFPfzlssvxXoHxuzbSF1tFMeja7Zmq3y8b4q7McMBM+EoOy1P
6jPTLO5VJXrqtiQZn1J1C/lyicWLGHDr5IyEBfq2IYT/+UkeHLZyE6svTe/pOgUoRXEBewP8Qpsm
mdx9fBrmYaE7pFJ0MpMcgiy66ZY0qJVBOPQXUkgRGl88qUEiWugWwitP1cjqaHhCVtZ4b3E4ZWOc
uHaYeP9cThOfFt8ZC6+Aveo8lZ6/x+4Lsw4n0AN76Tpxev3fE/Tlh4KeS+Ga0T12197VXYVnvevN
xujmYLp49ScT8ZFzpEcXSrIUaz7+p+TlHrbr4pkseyWXNt9gefilWuvtaJNSkzKkgczrENDsP0b9
qquws3ApJLhDhWs61+/csqloGBMjUhu3DsTnTigCL+x9udV8tgUSYyeb7uozaiU9GhaQvpbUbnPe
CaTZ+k91D4cKJt0L3BQWtsBvLwrKb1QhpdnGSLWre0kq4uco+9Xx7xfRln/9vmQcv56I9TW/xJLC
Zmqx/ZtUrLRdcw2bERPSNlCcifgnGFg2g5D1FMZn9mB/0MZppn8/EJknirwLvAaAC1pt8l3fRREy
8Lo6BLq/kHH4OKaozxmHgEIO3fp2jy9N8EaIiqEdSpcONN7FGvbz6atxRSEZOccf2NYNGEFuiTtQ
gFArK7OwmmfDmUfqbIHFJE1AuWSUNRKkxif21YMkyVUCnRa2l0l5bBoYh0Xu8wGmjJNOIawR61kc
vxJRe669/++TDxgj6HrRXAjL1wgmWZwSaJDzJMxxO3h9mQGnCvclrH/stdJHAWOIp6fMIcgUThMU
ouM6Sr8w6IYWH/e8MVBsU6RkKCMRfz6HZzlAbbvnb4uw5llcjFIph2V8wjo5mwe7vLSH4amjvkVB
7r+q6YwZKLDN6fhuDH1qPenhrXG6GXTwn/kxcz3lAWFjfFs0WFFkMGK0YCmy4JYaqpNIqSRZ/ktK
7m8TccxcDuUVSIwpUR0/x77IOb63Gx+BUVafzRyaaXrDfrzNtecqT85wGotkdKLhtQqgSd7KgV8p
07pTIBGY4yaQK5Sg/YWv25cBhSZLBpsrZtXarlveaK1Mujw4SQ2L+0wa8qFhLgbfFyx5cPJY1wtX
c3Sj5c4t1+vUaKdK3wIfq6S5g5uT+L+w4X1U2wWJN6MmqldR4Xu9hc+mTUGZspqoa1MVK/+oWbCk
oUPcnomPf5KCUeAW2yP4FDh5QHB1Dt5DoiNSVZTPE2K+okTwEdxQ4eSvnNSYPRvvkelcoSmVukD5
bBwxLdGKE6JhzHmKiHP6PJEUYpMSNI3Wou878MYNcAF9w8C4K5zst2/sl0WvueJV8Yuqke325mJy
GKj1YoBL3Wyf4zvCZIxBpxMG2Eq+C8h007t5QCNnOd592azp+0p04Rcw5iV28Fak+K7KyrxuajGs
3564y8j5Kfo8iJq0yIikyLUQVosNh9u+18qE68mRf/g9D3bq4WQYt/uoRiGcNri9luPaZP7sAB0x
SC6hY/DF/fDhfiSUXSy9NPcYeUL3OQh09pQfSLG6wNOwthL/Z4KRao/LF1QdFeCotCx9hSw0HPpM
d7VHAGWr1HaiwAfNA5dPSToLQfHG5/kEKr5+2Lm4R7XB3PmKW1xZBqB8JKdusimofXQ1XrTeIx4d
3LeLoBocd/b+nvDepCbDI4twvsSQcySpGDgQZ5/UraPQr5Be1vpD+rHRs6P17lNT9Tm9Os4zZVdN
PKdiT0FVTpq5CTjHmRkF3PdOPR4P7De+TnQa4BnrqK37JiX26vr5WyPnP/pVFANQe5AKwWPV3tdb
5nqMqo5Ziw4EXQmrhmsPXZvsy4Rw9ZKmYhQC++baXSi8UjkYOt6SmMGH+SEnbvdYwHOw0skNj2Pl
Z+eebZ2fYdxYRcz7p5IygfO/Girz4tcU859lp31XqWwrSFY5gL/fBSc1qRfqsFfwwObqZXxJZ0Ae
WyNlqCH2y8QFiRLDs3oLxc6fOKC4hx+dXr5Eu0iAZ56VCH4rebty0Qh9YOaoabJc55HxJ4DhYYKN
iuO3+4pbG4JhLRkxQmM/5bfi2q6mYkYlOhJT4cLqQELjPrq+3DTyA6rMpQE5NCORqwfuVEhut7mH
fObWYjUeq8Y05eEThENh19ActcPlmy/aLeM6DJOeWmK9WKbAKZ1l1o+P6Xb45N0LFlaW1e/DCAMx
cuSHWkum4cuVzdvqe4QXbiZLS+Ro0Tt36qPxd/00TAP63Ok30W7y279PGqJzTbPCgc21bncdA7sg
si25RIzfAJP3bcQFq0LF2bTKSkkGfRMM2OffhbrIupQe9x+hfBPMofjUsxz+dJ8MfXpIGkFSDFGs
VUiT7xFIK2r5EIEVd8ysce10rOU2dx05vSBqKzdt+nMwPAVWPA0NiwwKP46UZnBAcgw8x6sAi73j
3xoKiFsPU9nbpdqFS7y10Fn3H1VsG2wALm1JMZsSNnm0Scyc6hfCljuecnEseY4poinNbbfR7xSo
nh6SLTa9of0fW3tdbCUvwuitWM0/fIIhY97x7c2E/9HrK2K/u9em3bf63jgVFNDOCuBtDfVeEgv9
2p9/LvJfGtzQ3cQBqKjPWVmXljyI9nB+uIkqS+XClvq71h6j49XA2Qld/XrTZZJjsr1AQq3Fy+9q
mDQqq5+Sc6I2wukbyymg2TsDXLb7H0bHOxRIotqsp2qxH5mkppPbLZvlE+cAF4QFuLYGmI1RDdAq
f0L+5KyCINoywpze9jV8XVuFKx9ZTdDeM5xYNu0PoiAicQOJYx1QKwSRXR3hWsMCFNs7q6TcE60M
EHZOFKVyUMwz85+pRn/k9q98Gdns4Y2nbPDjK932BUQHck4LJIvzYyg6rmzpNQheDidYUcDQzIkO
NnpNGT9/HRFde1BE3NBlGF57gUnjn9en/4UcjRMAjUMYRmxQUATqX/3DhOowk5ggV3ismPNMzHEN
WNs9/nqOKzh9icLMlf7Q2OsEI+VxASsQy0G1fPzpgWTETrhBB6F//VX5Yi+pj2TlKw4+P2qRSdSp
Eo0ifRDzSVpXta+MRDuZgtvspu9MwRtVI9bOMt8gUCaTXuETnVxIL01zXw0Is6h6iKYYIajYIrmT
4z+/Etr/JkXYnH+JfUfjUl/8RcMXimrNGCCkm2b6gCfaMK6Fo9KP3o87JGerZ3x86EUM066kLGZs
8bwFt+ZGtrDf251T6Qxme20aBZD54ja0YaZ0MHD9KF3gpbfn5KAeGoke4NqeeRPvQyEitl0IX724
B/Jr4wKBFQEDWaEgawkgzosQDqLZ6mD96kQrTTD+ORhqOND+d+FfkUCd7EYGm1ZFzdsDTaQYGdsM
RLPaOs4IH0Kb4XKuYSHlMxUMPtM07vEQ1tNyf3zSZpwLh535UnxznIplXmumoAQQwTgi+WNiTgHy
6z2gA0h12i3Ab6e09rn8KJt/EcvQhNgUILl943FM/97706Fx+28j2PjwX+kvrGP8w3GNussZhzpV
5Zelro6Oy3xgHD4U2GEKJIaqMG2c6HdOtjIoS16u68GBDGB3I/5opz5+/AM+4FP44Au67s7MXtMe
cyb4rLqT2qlWSmpfRAJr/mc2pq18VyTuGBFpQQ0OACo4sA+cJMj5QJBZlWyPLOEpoQoYje9kH1ny
CMcq7X0lXzF1e9Ll/9ya5ght26lLFAtYLNatZIF0qREgqctai/GdXZ2gNg7Z6EmcFZP2MKWZcVLe
9Z9xwnwv+lnZTm1R0QD7BeU0SPsoCv+9+kDuNzf7e9D6vEZHR9arDw7nWf1V/IW0aPwCObs79oKy
evGNIcWEACHUTEra+poAMg79j/6TYmM0bd8n6k5qQgkAi9o77YH1e0yX4uwMDVfBFb+bZl3r/p2i
nWT+oO/Va1i1fC5C5JMGG8flVTxn/lQREF13l/43vBvmnJTjRjmPZ3+ZWRMFZpeyOzrzH9VfN3t/
gEmz0WiKiuvoMG+0fTn7vaI3CKbdYFX1SSQqWH1UnBiAJc3Wrzpqucgjp19tv6zF0Y1FxtphPTkv
qxNWSxSG9XQUaKbxlyMto6pwE+XHtRyZTcR+zPisX+Lto/I2mcZzP2PzqLkJ+qe2M7bHECFgAVIM
aRvz7cwMJM9qpODXkjARFSaXIBfQwutqLxS3c8ijG93qPF2vQlTlZaUpDwJbsR1hwpHz8AIA2rMI
h9z85qXMZwE8cyyrHN4OytA3Zh7tiXIIL49Alsrv5ZY2/TcRfOwh7PczWeXzanSmKKgd/H6RUgel
PqzXIw+3wGY59/VvgAKOte5oKPWKMZurjhP7lnLqTwCNmS5CC64awSOxXgQ3YsgdWTECBcp02TWa
cdXDTh7mbaj9WmGQS47s2xiCCxVKie3uR4lJL1aCqHJMgNV7H6MvJ/672Df2AoXtSQYH5UVbV5wz
oGAPVuumP0Julv2teM0HcEx6Zbgk6guAwBd0jQPLnlLjl08i1EPH6f+j4fE6ZgzJtPRgN13ao3Sd
kMShF/WQ051qrUBTnsjcGev/0YcpDI/+9S8aoKQ5AHdgPvwGvsVNKlimJNrne0PkBIvbjqe4DPDV
EsOODYuKgemeZalC91iUT8fusLH5XPRwcgagNPky+2mpbx4SlWes8rqsHgXwhG5xnKZtX3VMtx0e
DDaEmvS8GjH0ezRBn11Lo9dRvkfDWD8z3fakE5XZuSfxFdML2KN2UJKivG/8WD6IsdfLlqPVHjP9
MkxXNjUKdKSgTUmjIvuKgcnW6hgPYcEVxG2iQoKStb9HjrOnocHW13eaGR0hUJTo8ZKwaUY5Fxbf
nlfGyj3nqHcWYE2UF14pFldPRUqpF2quJ5Lo1aq/e0KHu7K9kBIPjE5/KYHgRlBbrMXJc9JsOKHo
pKDs023jsW/IUYE5L/Bgu7EA4uERz60mhsuGgajpMYHqIiS89WEJwXF8Zgeiaj+zlmrI1xmZxahH
8urvQNkPfUE0Cdt+k51J7E8wUBoEUrKvRksVCXeD2kwSCMjzkBPWuTSSe5UQCRhAbfklMkygwVe3
8I57WipiWDPLEfs33mM+z0aUd+oz1FV3Wmx6eOsacU1LTAafTEIqIyxJn72wPsFWbNlGrutjryor
qPDe9/kyJ2lVzsG+9Dy1A5F68HlcDgx0/BI8ienXkp2r51vEZNRTyKMzdMucd3vlJYhQzGXDWYgQ
1ZhSZiNpI2f/w1mhVQAWqNDnV886WicWJAEqLSxoTXK5FYnFJsW9Ha9Z3D4BPhGfROWhzhHebPAn
RG30WH+54XUmr4H5gMwTv1jUox0MvJ+KSGrQZP+oJ30agqZ3vq3mO/WI9oh5xbzFSVKyppf2mpAD
MsIAdCBOVt5n5x24XacWToZpct6AtEnMms+Vtgu55TNW00NdbQbTLpznDlqQS1hansV/0lMvuZaf
XpihZwXkPL5DAtI8n6NW2ZPLzLWKwKGoMXa3dHJiPgX13f/gv9Cs/nMEfED6oF87jmXoAvzYBcfo
H2qAExDd5KcKcdkEAvMqnR2YmZWzvLc0EjplA4fNAF+eyCtdBoS3U+BLlYkTlq69EfL4Z56UHuV5
9gNM7yqCii3JlIJMwdWhFjTcc3sw+tnjyX2JDNlUpTPAtCSpXhLIFaGiKs9QODa9KVoyCKBvwHhR
MrJQFxqIGJdYnYc/XK6HnER5o2GACzzUSiEn0QZkjzUA5BHU7YjOG30KHWDfLxogMxeF5ltW0JH2
fJZhlU7HlaH9ILivJbxavVAD5vautPN2p1mnEj89DaxQorTggTkM4Q1vWyGkDsrQWpbxOUB3k9mp
pj3UKcK1EVwT8GwNz+zlq4FzdzYkLYp7NEUPlGVAud0qw0OQdZJJ1amZzKGYTJTBxynsyLowLdvo
12v2UyXyUDTelKf6HoAv1YkiDAgO2OO1yrTEZZaEk6v6+tIgfo9Rvwwhnx7hNta8sMwhstPyt6dp
iAcA/EVhhp4hOIBFdwCqp67dKsPBt4hf01hL/JJ3QizNKZU1BhPCy34xdhhAMkU2F+Fx1Jg8IchY
S4+MpGWiZKP1CdO6kQ0g+9FQxkPtN1cA5X9TQLsolE1tL+SvGx0iDpbA16AetRryuzE6OrYFNTIu
3n3CA2iRr52fQSYPTUZ6zPKQu2yppYm1U1yMkHeD1KjH04r0olpUsRPsjiAi8+tjHQ73pASClxCe
rQKUdxDA8agEExnxfaJmvEqpY+FWD73SrvrrCM5K1qm3VAvFUPO51O1nFYOo2RrCltus+LEj+B0i
QtfQV9nAJg6G2/QYgtpavwK7fvB3UT+/PS3oBjw9YjY6SUR6JxNqtCbY7k0nF/5SRqGU9T82HoaG
5ZnJrT/VK/E2uWFO3Px1S9ytF3rbVfTLA6rI7tP+UfzDzUbQeWILbj0IAUKhIm5Kb4whElSa48zt
305YxJMuc0DR7AW4ADZaLcscEjMtxpQm+qTjjO6uwRkuSaVFXQB+YvSZYBuiZQ8SrWdjdlPSSlm3
Ac2VlvhTbQ8VuD9P+PF8ro1M+iWZtfohr9ZLjL+OFK3u+HIfruMzXpahuOX4eNOMbZ8ZNixBqQ2Q
5amEegZCo1nv/PdWS7jxuO0FZrKd+X4FV1xGQN1fbPYN68qPX7IAW82eaTCEBE0kM8rY44XMviDj
bKP67h7pFSZ2BarVEgdvL4mtb/WE7ZAvkUKLxTt0UPn9lqmZnZ8y15QRfKyaeAAw8CswrY2sFoSt
J/ViyzrkOLkpWngyhjLBHcCKMYAkGp3ln6jlGvjvj/uvJIOjCBD5kiMklQCdGQAENp/4DAE/FrCC
02NLGAr8Vinam7hO6N17WqUARDW46EdyUamfquL2JwxZMsvmdf2IvnPu9m4vbwE3QKCR3iiy8waC
4PFpSrjEVqPyFjeS9LI9/XQYh9pSCzQTVqDn0PbhDNtDkmt6cvsmyVw6w5WdRDsU1ts8z3NYwTjP
kVQOj9usIpGxo3oOUQbmD5pSII0oMe+hjKmWZYI7pVk2YFlG5J5+hjrYU40FDbEZ/tOs9woVE9qp
AwrwzSPkJk0G4CdT5R7+5qwPnnUkYDW38x8OsBd2Pjwe6XnJyFioZiBAET8noi7bNanxU2T4ZMVU
WugrsISQiQI23fHAyhNfvRA4izoOTFpPbwcsWVwZjew88WjhXJa7Bohrok5whmZc44I6zsDTL13O
vUfpRsnzvrhkpMwQX2Qonxk3roHI7isxSYDq6T93GHRtjpsWj3sz8FLNbLJ6RKQWRII+Pu0PpyNr
y4IK1bEymqiq2rl0V4kxU3DO++rkZPxb0RpIOfC4tQiQCl459RB/xazYVOewbLPmoJyRIJQ8oG0O
9ZHQNfHOfBvlGkQTmSpDuY50261bA4IhgychZpdM8I9z7D1Y1AMPnM1PnJo0f7xWYClpzEeXlCfV
2VhY60BstDSG1Gra6jxT+dAlcD1wKCVVl102HOJJILj+7B9lt3LF5/lwPH2dBPKQ0WD4ZxUq4617
Z30yij8iosD0ArB4AOSwEsSR9NJTRDBGCfZHQIz950heo0qjg41TDy+kyBetJXI3kWNbhKsKpN4E
r8HKa7gQGfmYYUGlzpbaaCMEgfZajt6BbYFBOFG34KVYn2/ce+vJVin1gingroy2rGHr0ZWqpohc
so0I17nyyXJo60Y59k5fr5XFI4iH3GjbsdqFqIX7yi+HN+uAB3YpeE3BkEOoBaP8QcTzUKpoJc1Y
/zbqgW2gGcYSR6D9PBcK8IANDmJdFXudh3Fk4yknKQYpKCBF/yZkzh5BEjpropTPnzU7ZQaOKaTk
LxdA/TkZcorPWRhEm4cHf128cxY0KdYHJinDc+0Odwa43TE+y77Bz+4MCk3aBhmTkDP145pkIg/9
VK+RDGLyx5BsMxNhi+9OsAWpOHw1wNXSwdTaJFH/QVPcVOIMrjcrtEmk28xp9arkuxsP/clocKqt
n1mCDjShdMspowxQxlnyRPLTmOca7KgH6ptA1aHssdZMdWz5QR25Y9LMEI6LNiooT8xjvRAX/oP5
xLsxO/v+tkW6aD3aH36Z0IQBakwc50/401IU/TQHhbGltJZ4t5uOLK2b/QgQPH1TkdTUoJ2LQHAu
5qwpktKS0CC6WZgVMc5iktY+PRW0fCrJ6k2dTvEApzahu+dYKctQdwh+g3fQiBr2YwZj1xuM5Ygf
pB0C6BzzCyCbnJfbVD7+VBQHN2Bq/bVnczCak5XwmZut3djtfMbSlZoZzr1MDiDyUn9NoS7RT2r/
ymFdeZ04BMOLZnqQjgGZ8cBWENCCWvmgzcpjaYV26fnLPha/x7rHCK1z8f9b897Fhmjkea/yeior
VANpmpj568mrpoYGZlQef3t/1KZ6JO7kHSgYjRl1l8/CoNjMNg80FV6Ze3P2qfseHjUbKV9jWFlV
DJx3U6exqbjWob+Nn6Ty+YW0lVU9tXayiN0l5JLnIUb6wOZw3AdkGLHLUGQquu6QDQOwfIz5Uj5q
YmFbR4B6ahojzNgpCkvP+7ZKD6YAK2aF4qTcGOZz8VQWLUkkWVN1m/ElCG/48KBstX8hTodoMRcN
O0C882g267daqT1ITga3xsS7A296fe1Fd8oVlp6DhcvVITrFXebSkG6twriNoR09+mfpWnAI4CDA
IyOqoLBrwXiu/wNJ4gA+f/KRWk//uyxhosMCopKGSgupkIgD0WDfs4LaWfqCX/+41R0zhu4jEJPg
34BGnSbUr65uaHVP2UQTa/bWijiIW06fH0S3rR+mdC/IUmZjfKLomOvGxsT4eF1O22KcXAhwCirH
GHHy4cK8CsG91MIQOT3u/gr014ZA/XCYi+Xl7z9ixXPQkCdkVBBCppI1VQ0bOw2Cz2fSGIzicXqH
pSqOEyg718ZTGBq3gi7miiJAazQwrOllsUemoNjvU81sj9lDAjWU9mgEym/Ciy1cJ6SPPg1a1pPn
RblFKRTiAWFLhz6bGgJBWnsXGsqtCr9NE+9A6+fyVZzXHEa9puATlZbwPZAiHgXKfmPtbd/fPTJz
9m6DGQ3CtL3AmQRRho6wH2I52hl85CUWE1wniGrWP3KVEi66sATTzrQT54Kp3U73yAirEDcMMdub
q5AbWoTNda1JiXgwnEm5+BX6YBs/lWrSRnJSbefyFXyjjOx0OMmto0tD7Z+Y8c80z4lpwxph9jcb
B+E7NF4H2tEIJdJHtf99ATfshVWPf3MxjtwG7WiXsPVRRXlV+2R0/naIv2rRaUVt+cwmpvPyneB1
h+gk+vs69ZO/yu+e+ziB2ZyM7PS66qYFwaVwNfCdt8yY69pABZ5ZlNgkgDO7Xc2sazEn6KnB95Sr
h04i/+68rs5faF5hmk6wYotPYgxiIa9beR/9SIFk9LJO5UOwfhbCM7ZzqA73NZbpmPL0QaiJ7wHz
Iy72Np65fxrXOZWsS2azZPfLfQ9NmMgZh/4ED4ZGFpVpOjhEW5sJtx2Pq+zJtDv5M+P4nH7KAndZ
dMwM97iiS9xikOzblQXK+HEloXTm8pTae7mELqGtX600nA4l6xs958UJBYPZck5X7cyn68iOOJzY
K/4WH4VXbPxKG79OsFjE3oX6P5RndT4JqNmsoTW69AU3VBWL+y4Hm8beM7h1kCe5FBU1T5tHhFT1
z2UcYN0jy8aOmBwZUotUlvEe3czmm9PJQIQHSQmuFhWJFuhUtmQOarBpjThV8bNABBofc9a+6/zp
tXc95x5w3KAs6L3IgOBM3DxKR9xJA0mYNzGUP/8hQl1LhZRBDKFgjNyRiq84SvDd28cNHoh1SbXX
oxk9Zp2nxhUUxaQey+J+Vvum/tcjIdxl/4AYDWL4u0myInfPK8v9kM1+HPSqiSZjmTFz8DgOIOtl
Xwz6y9NB29QTZPsvYlmbZr90ZGjA6XgH8NPeVWsWnsys+wZn2AsnBMQvFFziQYwpcF9k1iZvQDrA
mwQCtuGEuqsPf2gRQs78rrdk5d1oq5sCzpYHoiJtIN+qtvgSpNnLHwnXwqYar02wY1F/5cPzz4UO
x03715XOqaAffH+3Bw6mk2gnGLQQpfSrNGbf31f6973Cr2JrUvpWdm95Oot8/2n9alQ52xgAcWNF
pW4PqbJ35Nk6N0X1KxFR6XyNdo/2wiHBPHW4mHudBAzh2i331/hs5ZIt0gpRugDi5K38S0MjSsJ9
Ik1NBsP2d4AJY8Nf2Z5C0rUSJ8LKjDsW9BOPGyJn79FPzNoJGtvymeyuiorg7Rw92yVf/atNfiNS
hrbKN+b+38Fa0vSyRSsbI7qeJaz9n81BKJmoX3fSL1oPcMSR5r7MSxARPDBoYhVbyk1Hpq2wW/3Q
0KJaM9U1qVJN9MUscJS/e6lXIbflNvZ0ucxQLdNZ+OrsFP4vf41NWGzeYYqFjZuVpKwFrorqEi5p
ui6drlsz7DcEhBuyIP/UeDIXA+jLvOMBJ0mggv4v0uXl6gQocEYSkB+Oq4shDjrdFK66vWDaO9bR
HIk8a/nz/Euv5c5gXJmlmGOWCa5N2a3w8BKLTzb/P/RASna94D4Uv79jkrJ8FKDAygV+K3xqPf9C
sDHxr6/n5jB8qCbTRi55IhfThn6SYm+Jc8Gyj/iYKJgFqFEw3lJN8nvOBC1u/yMvCn6Z5nXPJsNY
fhXXxt5OyFe7WuD4Uarhql2gV/gJPN3eVxUG5CbU36skRK7ORj0DbMlRQYjaOx1yBU4/x3hT7mEO
TCajJ8j1yoeE4z08/sSY0mE6w7GcDo0RT/o+KNvN4lktOcreY1JJr7AW/aBm6iwONReVPLqsA45D
zO9rSO0l6qQIo88oCPx3iKuEo9AiwNn6tOSEmX04nin+xpfIavjGxZ+H7vJqAYUlS7IYEqa7+7BF
K+3f0tS9G7bg/YIzXzmlYT12dQivv9dYUyufBEnYBYujdHy5fQM8hesPz7mqsO8wyQhjZoFhfODH
Sevu+JG7fOHeb/t4d3pP3lRMtzdWl7vUYhhIUFYZ/V/qhFNss6iM+R1pd9TQDOMrggQa1cz6bIL0
Vo6hBO/S/EWKSVVWxJOrcZKkDb8OqF++4oY/j9cU5BS11cUXqDcj0k24pvD5zKEg0myigOvhO+sm
h8KIHcym5Jnoo+nA65HJAPpEu41lJqR2DNpGdz38EyrrcPAl0z6hRBL5kI379Uq3mf1JXWT3u3pS
h8r2ZjvidHOesxCy7XCY43ZIAyi1QKzhMwMHGQ5C0ZS825eIP/CuL8jOTScI72pnRQo9NOh6iAde
j1Q6GTG614AzFNyU0Zl72QbeYFbTPK6P4PKUQ9e1b5/2TfCIaczC9p/9g8fKxv9LGFT1LD9i7yeb
Z2xWRCYTNocUZFAwx6XXvc4ts6dRrbjAhH5lICHvpoczZoLsHBBub8mYrlMDOIdQoUVj9+FXNCvY
GHTTMqg5gIBwM2sAvCxBYjTFzwJoxhv+lz8tGwYzaNT0xNkvXO/3ocFQAn7ULXIufu+93epg5VjA
Byhbek8BjCJMiGSNV1K02w1NDeS+b+QSo+axgSCCghsApDG48+4h2tnlgE+CJWiB5jTSyTdT249H
rMZJ6pOuIFyLO+X6ZrDXvYyCQSskVJjgan8z8BORvn/pjMO0bFF5ojwFVZg372vS8/xzLmbfOG/m
UGQxJuPUZ6wIyJmnzTbgEDbx6TeUj3aQCRDS/DDvaRhy1CMaQrlvOvPc3FqJ/T8POOFjyehmm9sL
xjyZ7BdCuyZsP2Dn7PUiHoYFHtU9RI90uc9TPohOpzb8cm2BZV1iqFOBNarX3qsLfY8f7TQ5Mamc
4r4CRAGMgcMPkULjRvHtRlKsdWFvt6Pe40IE4Y0hOKP13sKxh9UMcXfivP+AIgJzaQdJIsajP3Oa
THop0CoQPxdmdeOZAKNKRdmlktNbXY2cuesZRegxFfuv+pUqBChF2eeZPMkmi25SrCnx8izElLl1
SVU8E+Ah4em5is875fhE6XkK55rUf2cP1gUvHb1aeh6+B9zIPRVwvPB6edNKsWDg6BzpGMVvtQ5l
BLXXqZ6k6d3Npa80GvcyIFMLd4+XNVPfcD4Ap3J9rd7F8HhN4ADJ7iHpjfCXCfo7oDbWQUNi8Bl/
WgZ5GrNdeGVdaDXDX6hCQcotoh2tjxlfYmVD6e0K1HdqgRL83+GTupi3MGrRGbKieEYBrIR+iijT
pNHgWirkfY2MFwxtnAt321VkZ3LzzPxALj13fsOV/CguSNp9ER/Mgvr6Senn8/6KNYegMFAQecZO
ixJMeRXN73itudRf0IEX9SZj6tm7VnMFfMeBNp8V19S/It3O/GpGzu9qSPKFsbhyr8vIp3ZtOc6G
pjIFOMkAzgl59pXFJgXsv/63XPhlveQEhm7pBRbuB9L9FedywPFrIpgJRA5FfbkhE4AdyCUHbzDX
c58eWI8n94fKP3v3aFDGzxJc0vQpQ1WMd07Xmj/IPfomKBKGLxx68pE268z5WjBL6FJSLO+Y1gD3
x85JiaXVipReF8z8B5ETS0p8OXwatFEdaBiFyivHd28NfU9x/+0K1nUe9pI45d458P2RVb3u/NjT
GBhiEFqUCeWsNtCjgVg72K9pziqHggHaUo0IJnDWuA6DMYm/2u9HDn0WVPdrsk4LDrCN72kgUlv/
XcFPHH2tD1Rzc7LuIX8ebqryPQYjWbBZ05hT9JRKHGtmgiqEvG9EO7SK47+H3YtnkjuPDdDPSGDv
VAY7Spv/YRH1EYXhhn4Qhrw2mYnKuNmTSlI62RC7xaoktcjzUHV+/fdAj8nU2I4e3iNgVbUo8Kwb
WmGA2ks6/8fWM3G65velWcy7SCmBrqWUJy+iGQ38pW7KTBmbAShIgZEfPuM1wDOsfABSF5ncb2uv
XC7ZX4BtohDnCSlLVDZ68e0frC1azN1YfDHS4iMdrnsxypejJBvnpnmklEpozgqqekCnZtNmllkp
UsXSfk+cvKwekXlRFVc6hO5k9m8a7LXoocTrpwzUx2Al7bBr+sOeQullHmcC1/2nMDXVta3jnY98
pGrJKH3jUdYI6h3GYQSL89kRdVWlPVa6uqy9IEC+M4v5/yyReKIFGTTZfph9TjFtmnx3Q/XxmhhM
qhpfSYVFpKRKDhYU9UrZKsVnPrXh7HaD/RvA0Hp1T2seYGQFkparlNUfLKuun1VHwNIvlVOh7wZP
34XQFSVN1zpewDCXb/Zj/RgQc2SlbmfWNer6Ktlz1V9OZv6OBR2Cf1mSAQghkyc6nP6x07lwSAgO
mKJJgi5VVukQOjn+VYgqDihOFK0b8tLJDDNb+RRppwIblVH141F8D4Ak4z8mjP25RSlvbI6r3vwX
Hy+Iu7+W1tLIKukMt5hl9FaIjLlyuLLvDg+7oyv8wLF/USXcnYI//ElIAwArCED8um7qIJDCLQnb
2lhxaeSMZ7IGIScjsWm/NX5QW7I+NkVYKI/4CMWfbEitef1F5sMUazFWRY3c2ZBLrf6nLQObVM+p
hSZBnZELh1ALpr+rC4T7jUXQmppYxhUkVn4IU3iIMcoQhSQTkPALKSGyWcbzfq2otp2EJDBd89zI
E/UqSY1YV/BZeUQKm/XhwGxANhDz5h0N9ysmnXDe8znvpR6DMac3pIQHzzb+9Q4Aw99nI9w3t7lb
CIqZwJnI/5QIbBFtXJUjUqWWclgyAF2h5rAMV2QNrwUVrMQGoLZDGAnIAdiYeJC8xJ6oDu80xBHL
4+C+Vv42lutZxWjgzhM+NVTkCXUI7OWnjUS4T1WN/GPTm+uM2ws72qj8aP8YeHuwMLCajzDsLSv6
VDyNWGOBNaSb10OIyM3bcaVi5bkzHrzjIn+YI+poLS7GtgF7z0qOxMFhIg4bsxOdPLKN3nMIg2oS
GNYsmNkH/I/GOflLe6aKTWYAFwA3Yi+1eHVr3R4NardUsGCpXFm2ZkaZlpGLvQyhbY0HchkvhhG8
OvIq9bY1nGpIQdBMgH+kRzmkP8Wlkp2VJCVZNi5VV74Qmv4WITzvy+F54evq6+RDer3zSD8SViRX
L6gMToCYgM25EUcgx51PaUT5+9L7/7QCWEG2E5kmYwv44BHYDQQiFOQP888WYgFaBe80m7Dm+5GE
tv6SAr2vIc92+tMEj2rVI0rLHwZe4sx3ex1JOzgk2WMKwIKEXmMvfKaSepDyac2nbPbK+cBVVpu5
F/6riZay/X6NGv1at3RRsMNXAcrrf+QTzVbCOqSyCWhlPflfQDlez5ZV7ZIZ9Z/eznB93F3am32f
NG04Wb6oLrluCCONJo4Vv83sDmXp73FwO4CNQwhY0fNlzGplBxDQjCsWAPl1oiIsfQRgreVZt+vO
6PbxEhNFXJEdDREtYtZer5ne7ZjkFAwzr/FFTxwYo6aKTLFfa8dxwvaHxXYIc6h7s9EWTR0q2S68
c/rcqqtKSz72E8pf5HNYtQdgH3ciGytypBKkXIt26XVujGqUWuaRgsaq7ZzNS4ez4zqI1c5yQEC/
uy4qjXF6R0LiFKiy3bEx3kx//qwiWk8Jr4Ntn6AsA8KCjv2Uyvy4s6FYkaeg7t9QTk7fVQPcsK0K
RV/hei8l79HJ3J2rHKs6k/ztXeqbyVWK7gjfF1q4ZCH2rjEBvubJZjkvdwhwUvxv2LbPMUtl60Q1
fPEJ2W5gTcUFT1J/pw4QdqRDZUZrPmr+i0iffaVNtA3Eks35OsB22sSj7xvCLHpaPm/s3qQclpW9
Ze1MET9Unai9JP0M6WU5K4cauOevuKgh992nOuZ4VC3+kGQ5upFZjaRXhQgLnS0GzBWYmnAxQlxj
lNYxAConZWoFLsXoP7yryipwLjDNpd7m+ZFcISewKijqCdJwCHODNy1B72Z8d96TC8NhnJUZB0lk
PD7czGHIIMW3mIQ6RNwkYq7oaSCcN6Rw0GI8JD+QzCyrK9NUcBcd7vcz0MEno6UlrQKnHou/06B0
Q8cmot5bvQiJNuyuQk2U5AtgkPjzvW+bDgViWoMJJzB4BPzgmMuDXbLk5vam+htehel037Bb4YrA
ekN7F3j6fPnxfJ/X3HsFszrjBC1BGg0e2ixrrGGJ3MKqzNT4vPP5Qm6jfHR5u9t29tFLdXkA1JXR
7aPdnED/f//Epx3HOVvO19FYrizJrdQgtaCDLfLIiEZgwgBi+ZY7lKeKVXrnzKM7fmbQ0y/Yvl2l
psKPVGNh6zZ4zz8tcFQofIz9dCR4UHbBHWPdNieClypClZDtXi5QP8FYWVdYzgmfmmnJpRe/UrUv
3k+a6sp4wqmZIEaRLEjl6EGhtgwJtbOoaSZYKyWy7wdA967rrIaJj/F4yvMXQS2HP29nL/naU7US
aGHxKthKqqEzc5qHZWgm/5ZLQQCpBJuki6+kGTFt+11tyqBv9qyRbROeBbl1r0EPFCDUowKwUpLr
NCStSAsdd3BQ9P4fceuQBuA+x6wDO+ElGAOs2Cm/ZyPgSuKazTXeYIDrm8JzXhToNEEWlWCBQw+G
70SkAe8SUJ2n4cwoLq6WPxdFj1B9piqpqiyMoqVUrVM8/tTsTkMIk4kPz2V0FwAAiM0dVMyIxulI
iFLYzb7VcnG/yjmhfTRigPeqpW7w6O5aGdaqSo/SGR9bn+gBphHt3XlkgsHSTvFGbepnOhryBd9b
W+1Qwv1wG5wk09NA+6ySz1xobWyoFNuIEk2mulJFj5DiDQmakVjob4+33yQWMH/jQUzHsQCEgvfU
V9vOtZxgrHzBzCwjs1ajSZb3Iw3DZ/nc1kUHpn1LRr8L8N7cHK6y24/vYN0Xqd/jHfb9vB4YRGnx
xRyr+euKwzUqyV5vlLISaQW4D2aDW/pDdQ4jgEaH4lWcewvs+81XVeVZGvJbr9LTqw1XT/UMMMWM
3n8rLiZI5XrUQztyET2906ZY8/jXmg/sYviW6G+D1ALXnxDB4F9y81eA5nTLOXxBFbscoKUXA9dE
xN6bwW1S1CFiDt4alLjeEwdfpwwzdj6wvhnLuP8wjpP4pIOhRCLfSXN0VH8l41z/ngSLTGm8/VLF
/yInjhIhHkY/d+h4kaYgMaQ4b0qiZdZ6TF7vqqlOCijADXimG5G1BQFCZhyjBCj//LQTMPt7uZGC
98pIOnUqViJY334ofyy5d2xi2rpW6lgrOlPqWkO0yTTYagbV9Ums3lv/A1qJrz1i4zGdGtBgD9H+
gc9CsjFc0/DdiOndwSyDgtvFxbG9CtILw4ofcSv6Usc4sVNyTsHr4QmIHUWa5T9BonfwXlvG2Lxo
NRNmOMWwe3TOINV79wQF+3Zn2mLN67SYpLcgIZwqfLovaPMCHS72HayDPsTnAR1JJIBF+uESbpAB
sVPi5HrvvGQzrwhKgrD4k+9e6IgazYh7n4EAo0EkdfX/x/3LX/tvZGxNbrw4ccP4LUR+mxY1vAHd
ZZ+jk3Mm4MwSa9hZUrlEqG4EI61d+M6ms3uSKp9BnnWKmKjEUGnF1G/nZFN+6vqLMNibhhoSWdrp
0nbySUzgnJ0KYOeVpCAF0r55pFuaI4mt05gbzm3IafmpGWUEBLxarxhi62fv6uOMe3LwhicgUSlp
34x74IPnIW7H3KuEwLNMSBdzdiFfnS6G82jmHMQYy5oZBlql9Ra46NWI1D29FHSdc2VgWEEkfLhg
0iUKTh8fHb0Q50gionamllgBFmesEViCIDIIj7s3tO5h2ElT/B5W86JlrNE7KxJbymDO/sr3NG6H
n14EjxtkP3A1pTQmJk6Fev3nw2Hh3rw/EbVMO20RTUAa5pQjdc7Dbh1EI70j8fkQj3oBcxIat5id
81Rx++E2x3/G/dsEuGfoNMHhPhN0GhtlkoGasqOmOI4N+ajykg9Z8pEqY9TcSDHnizbDPfqGnIZy
GMzY0dScEeykEgQRuXIWc2GjKGdhEbgN+yXJF9AE1SpjaZCt7QgV9ZSB8zZrD9cIgs98LaG4R9vh
m6mqjjsCEf/+ww+bc6Hkut9/o9Qeu+2zEUsFpAvY28+CYo8rgJUTEmjYzJOrbQkn1uIH56OmyVaI
OT4AqvjbyFzDbN1nvtXlSWJh13U0paGego+hWOwu+1lyzxHR2p20pIMiRS3LoP0E91fHu5Shkfsy
lfslCW+qBo8l59TZAGYAT2yEA2XOyvtGbIT5anwb6P4tivOdf6wuMHYQOX7gCQwq7SD6QDvKxTbk
osS+p9cTXq/shCeNKvFmvY0KrWPGekV35u9yk3y/ndoFnHVDhGbtijeMHRxEnfArclehedJaLLVk
nA/2G8FaQC77gjv6mc+/sVtlP2/O4X2zbDdYAnoDfkTp1TwQxwDyzkb0V3+FiSVYrK/LftuiguqO
kExnUxdjUhdO0Vl2S7T8dvgJqwj3FLwvhWL+7nI7DB7jG7sd8VOQlC6yvkNM5o/XQB2kjMw+FQ2T
hjcc0SmfC9jzrrjjd0xQggxwCKBlvr0l5Ur12H34keUOekly4ZJFCwEDbtftxra4uddJ4PM0Q5V0
jGHqejAKRSM1gMW8wnu4JKVSK4+/TnItabD3gMsycv7AkizVmcTkcNYHMInyPO4Q2gZmKR1r9OFy
onLyVPl/LAGeMgp5KoEMEFGCcxSUgBsdFYz6TDTIZTK2mRS6+3LdWgdtCNoeDdhAuOHzQndFPKEz
6qbMS/3KPJrz3QsWlPXK88uUe5YjPfwq1dT+TfDKzAPSGd3NFnJ+6Dt3yaLeBQ4M73jVU4Ujke2e
Cld6bgnvNLP2TmSYPGO9DCukeGBLUNtdPurbb7CGmecfLP1fZYd8+fMCO1m97UIBCwVvgksVO5Yl
GPZfVmFbJuK93hsJJ7OPYio+A6DNXeyES8UwjiUpZKcPFGNx7fTvW0ipy7G72a3K+OM71nzYn4Py
UIIvAvVTsjNIoxo2I224uL1SNXjtZnDBCguO/riGaT5+6+nXR3WvGJOu/wJReJmXbrUbABnshTyD
g4BYTIhdTjI8r84X5spt7gsYuT4633TEykILECnJYyQovL6lH8IWr6tlwSbdAlzNFe+PieWc3f+H
V/Ssjxb6atdQJqciFnY1UAZXZG9pLPioL8hNhncCjUDQfmxHEM4ywiPV19+6slYywFsdAZ1ENW4V
MtNtF93W1APN4wt6ic2ZVvKYKxqft5eMkQIy9BU98NOxqDLaU+yYE2SRYTrqioaQKGO99pvnyyWP
OmYL0RAMuB61XZ346obUkl7NHEhqjL0ISKx5Y+nnaJhCfED+DD9G6Gd4p5opo7uDMQNuRlMCk4nu
6EseJw9LLTyuMArTV2/4ZZRDJHojd4YKG9JRMojdbaoT/aoKhSCxKzh5yMSFkPIP42+q+ZGPGeuE
kECFedyVk8k6XJdt0jojeCvQ/GOJmH+LRjp3BvuvhnFvAFo6pP7BFHAK4qIpd/3HrMUAx50lGgSF
mFqUJK2FbNhYjmK6nZNGlFK1D4yVGdNbkVXdQgrKj6R7THlWPI8HuVC2lki929m6Rtuj4M32Tmam
TbK6vYvQpPfss4Ke9/XmPDbH2C/0tS8M7UmGYQwghrfz3N5uB2qxH1UgjROA+E5f0MHb8CwiJRG4
WB7xZPkUz5lB3c9hVfrSbPSWNr/w7vEJ3GF6q+w4ECLje7BO+DFPM7cdN0mQcsn9cf2tNrEru9ld
N+eWuAro42iEgGjjJTxfJGOPjUf7cTugCbPHS72p5a1F9Q6A0saynrnZ0ZcK0bRucGAyhq8CMXAq
8i7kMk9C0IaSKrjgsxDG3XdFq091/tRzHB64cbxOAoGulO+oPxudbYqdm/4pqsT4zgUyYTC92cFT
LzLtoEVH8fuiS0/PqtF3n+0EUDht2lWXtiUzC3posOghfRVmPGgcYyJ8yTzlGmvlhcLFaFt1c4ms
45WlI4eV0mgWbgZVXKsmtw/2Q7McNGMVsrdbIlb0q4LhnjO2tAkR+sYDdI+mUl8xE80AcoB1XDtL
oWE0z6j2sev6LrWhPmjx3z3X2YdzCcqpA5Qly4qRURb48/vwPaI3IEA90u616ve7wVOxsAFilYSN
9GzGrixuBnmpqjkBpT/K1OAAyHDZb4Ctvgk8U6C/ONeR3YdwDEl2xsxY3/zPuTIsS6F0Oa5j4Pm5
67zlp15jgBfs+WUhu9ud0B7KqRC6bZul4mHcK7YHaE6a03a6vQoFfxJa2lJADBWvOKzPEsyiEKOj
gzfpjWafu1Ahbyt8dc13wWw+a/HHexxs8qB89pRckaoorsBIZeXhDNtAmclE/kpJtpZHaAtPsKmM
12Lk5M9Pyi7PeC8/MH9Tux0PtRL6LYM+KoGXvkTNTyWtgzdI/1FwuMaXl4pIBfZOw1YD87YWshw4
WpcK2q5AIXwZp6AYQCKB5xE9lM5H8SMvoswWcIv8ctyFc/hcxnqtY+LLTXCInA5AAcDrDSSQ6J6L
cSZj5TTePkNG0swqCWjie7kzGpxltqahx3S2UmKxvL6Uh87ClQzRpxOXr5KSXv5Oo1BNAd1+qAEU
+ZlgpFGkgqoJ8GqH1T28/YPmjqmtgkqECEuAmWAIVf21dGU8FRkXWzcoQhVKjV9oK3RrxGf2SooH
hFOKionREZauPBb0fLlktPkw6zx8pkrLAZ3L0RrMEYheyYQaC8rirIad8F04aygZoQTYKknjqKRt
fO+XorPnbbe+RxJ/LE40HXfj6Z+b55CRPs6CUUe8oGswNSmhYCqty0DRZJwovj1DzYNmvwLDurw1
MXXPQVwfyf8GxB4GkPLXV6YSUDAcaYmZHOG0sEeJGVXDw/BMxzw6dwADaVWANb7cjnPFUui1aGkf
WIim9S6yMczQyE6s6GCSY2sELO8ywcndFPHbKDwUmII69/SZABmLynWk9qfY7TjMa3ZSdf0eZbSh
ADD9Lkhk6T8EUBNeHJiVvl6Enbo23FmqF7LGFgvXkki5+qBZ92up+fV+SG/gWv6qlQbq4k/6yQh6
sDM5OkKzr1e2KUDzOPvdb/ZXiNeblIPPzYchDvYOXi8UbjH+Lr/zDH+NCskHF2Iwkm0rem/bqCVf
2fak96ke2q7pVSLMGu8+tBpGk3J5bp2ROCswRMXpsEQDwvmdeQ6Q65mXPOp80atdEEymIMaoig5c
NRpDu1see2PpBQtvIkzWcSL6HDaU4CEnFiiAjT7oV14tZFhTZVvz3y0fW1TPhuyuVswsipz4gtlQ
Cv9MgTut689IndqUVIptHDvLwYRZ3LyYtQS3AoWVwzFHfeRU1ZtvB+E+1zpdh99OODvn5I5XcK1z
+DMycvnaEgT4cjmRCFu4edOAHWO9vD8Qmedye1AO7V53RqKFGuHzL5H9rEhtm7qdLBiC3nuS9uBI
wbhNZD/zCrXwjjgt98QSNpzEo97lCqTZN/DyRhXY2NIVjGUb4AFb8k4QcdilWy7zE6bDtCxQ3TVy
jI7PZgCuksd8MCQBwWrIsXXP2B5aTKuAj7yd6zTDWfKn7Lh3yt1ATDrl6PTDtD8jzqbqGSS9fZBq
3LB9wU5XgZlNHGGu7OeYb4HF3Y3asPHsgKylvO/LfOc1Q0szSqhhNvemNQYE72vnZeSf3uw3R/wv
gf+rzOcmsl6/TVldmjxziPLYPAbhPJ+pdiDqGG24r/8KaSn0THT2PcFPGpPQqoGRPKCYFat0Q0Rv
/MnUQpeQuAzBHfrqWVbAtytnK/w7dDiWZyAMMJ1xrDGKgJtekp5nwT6nBHpmntLsUgFy9rQjzO9o
7irl97qziHczqc3XjG1BA43DIttRW272wuNziRAv0tdYyY3zlucKeQJ31kkwvNhPJl0zVffC1CrA
d7zPWXKiJfMyEjmOXb5nGceF0S+DL2hHf4J1UwtImTKg/rxU9ipUqf+47MkU1eH3yI01JPkabrn9
Tyo71+bIAOFtaYXkIotlQ77zfO4lhFR3d1/5/o/zerYd6LrUOLbjX70JC1AodWYYWeyeY479DVYU
HnR/7xQF4uupJuOYvCy5RYlnnNTy8ti6lkn64Vg8ATcJOe8j4O8/TVVF0yAGA14RenBr1+jCstu0
7zLJTPlSix9uXBJJycTu1Cm2TBbKwi6iXSCTJz5PhjaJH43WYE0aKw/7OXeiw+yV07YS7zjLJcbT
nA/2D1RrBmXQT6Nc6J1cji1uCgYuF7Zf+Gnj4DelZ6MSwMHRptJO8KtGayYaUs9w95WjVjeU6Xg0
CMjhYwhlx3WZalLkww8T2b/XBtXkJ8CG0E0j1bRSKmWoEOZXs6cq9PZiOBw+ylj1oUz5HP8N9aVz
0fEIxPYEfbXy/9AzJZT9pYbPNhFWEINNgcD4JoXfV+azP+IPUiNTqqx7hbSV448dl+lyix+eeSe+
pxrsH87lgjT2uZkzu0+eZQ+pmV3qAI6Ye8eNww26wHucfCQSHGjELBl4ZARSSOROzhk+AZwVsL7Z
yIBqqKnpkaYslKx1zqZ4v8AYNu8II5sE4OX0xj0rJ5i19GZuz0fmPERlkAeSJ+qBo//nSFWL93Ia
oqsoL1HBACT/6o4vXU8dG6bE8gBSsq09rzjYHuZpJqNCYyrl+bIMVsvA/d1SODaVHr8maFKOODyT
XKdCw4oGVspkegG7pBkqyP72VxLL3FpHt55XJ8dLT+XBh+JmtsFxbfdJGTdvtDBhuepciFk5zWDM
iqEtho6HCDIl7knyMfZQ7QdvCAtfwaN5lE3YA7to0oDY3z1yTTJTpjNLXZMd4wUgPmP98ZFLzBOk
pRE7Oz91M+WLidDh1Vk3hkHYqYVkN32W5rYMUXpnOSPD/OnX+FBX8GfM+kvBSINHkot1cKqTYyLv
L7wJpQDKZfezFNk8gyQejlM9wURuBizOr8yTHmzsKgkS7iF6qjMjtqqEOOjQbrCHnWjJrSRspNyi
ZwiS4pzumvtQGd/gCvg08nx9OF4AB9FDqF4XyFr9m92+/U7ovq6Rv6+kF75XnEyaPkG2gz0bEw5Z
jeNh4+UTKLUd0dp+6gloeOYGBusD/i1RnzvBUJJXeKThdfuGoZhZHHaqHDNuuU/H/KNHRLdvLY/I
yyABIFuUcpUsBnqWAVqRThANaIxo4gXNE8bx6LZLZBOCxzYAH+g7pItfTOQUuT3DMX6x6Zdhuviu
Dtjeh6mdUZTD284rtR6CXfsM1r3RljmDRHpc4zubwG5BSOBEWgpk1hzjfZlMt09DUJ2VKkF5BQ05
p3s6mHYNMBJTT8FU847gr6hO4vSftpkI8elZuB/XTlWaR4EOoDfQWW7vCMiR8z+aLRGgvX3bHf0q
pUty9vSOAf7AKeBSY463V6M8kz9MGTrLknP8eZsJRsaGEY58HeOLppfImxUpVJMRS7iIXevKwZuC
IJgE80V5v3hmi2pdNQYRi/Ei2zrWI7WJAgTiIvHTikBaoQ89Occ6K5M1T/4OsBEZK4xzghi/A/TM
CuROApL6bj386Xcw9o1rjaxvQlURq/HD/jMZJDM2d91M7hjijWbO6DZjQfwqz/PKljSfcS2/SuaE
Ob5s4ACoBaMErIKBQhyhmw72Mo1ampmdV2TKLcwnqBVD/TV4IVx+amsmyRgncZ5uXdvT2y99c6dI
adBYsxXn/q7nGl5LHVmKGlCPQvFZ+QceLqCp2bCGei/s68CI7fSzh/WF8HUw5F9oy8KOY6pEC85A
wcxZ6e6LMJykzZJh9FuZXW74HZBn2FCaOiDvVfgJKNiXC9tgM97cu/ZcMiFQV+uVYqN0ZE7jy8ha
M47pZiNMdtTlq7pf1rTpj7nFhrFzgaf8HYEQMkL+CtuMbhDzqa20LIVo84/QzajrH1jFPNJGYKp0
olLHHNJnNIzG6Mu0KHEUL4Y+Ahpeibx2PU/QTdCt0uPEEJcUgjjyWmGkxLPTopGBKLOZMNMVyKEM
jvPgxGRyF70eGlxZkPyQUKN2hiaOFFi3WehWaPBaxL7oTqtcLeIbpSjo1OAFlPs5sOmzeT5wovqf
JGZTBT5TzHqOtOV0jS6+LPKlBIMg3hR6pL/RAcmwCh1931+F18wJgZlAkLPnGARqSjaM2A6xcX4C
SJYdT2ZL6ctAuSk6dnHs70QZxqaflRqlspY219Fs9jwHsXSUxf9GATjG4gYkz8nBKWyUPrg1KWpH
klv+sB8KrOty8dVz4eQS28sguFiBGrV8WgYw5VWkAlGjo50uvge6lsWmEVlg0+EvIZ/iwK2oyH+L
1LxFP4O96AJCB8w1dUNrjwrClsN7G+ZEcngctzkDuzZLEEjqUt0CECO1AlIV7XueNY9yO1w25/am
FI7SzDEMpdEoZkWDaRWRv4CYQo/6Az+Jj6V8w79wt4PrJO/irXyWSEuGRMgCTgM3lHf9/LeRnY1k
1lbUP+3en+u0yuP83nZwoZWOmsF0M4pXeIAZnwLxRpg2TXiNW4uKiEwc0YxznVkJwrB6bbgQR6oY
OD/Y+gC2ppYRsA4gqI+gKL/C/bvU9AHcKonWq9iNeezwr2ekdVievHSmC9LJgkGVvsFh5zZIajS9
ahCRhw6lnohfTjsxl3z56eNkDEpRiG9xhwoSJtGVU0iymQxOjber5flPhtWctaivSKCjTQQDfFjI
7KZlAZALZ1/1Pj1ciy08/Q9Ivn9cx7Sdjm37z2uJoH7CgFsuJ3AvxaYfcxDf4jQG6xgS2yZATSmh
Nqc6KBjWyijmecfzVpzSoHtTzboAzEiRA63pK5qpKGHi/8qAncQnFsThtreOPS8mmMzPlu1S7iTe
xczCnFyJrcnZRwAtOntbAjGozuyosUL3mmbF4hYUOhIxYlHGEY1YvFUTG/tWrxGVJzDcJH4RbFjx
GNCa07nBifcv8ChmsiUqMwezkm1DE7eWphdPLzkqVPX3k83YpjwLNP9iFhhMjRDeDXqrsnSCSauU
sAhBERHU259mxRoZ/E19vpP/ITThn9tuLGz82Tw7l07XIyiFpUd3zSGgs/7tJqtBnSR9lCVqrz8P
T9zcRDq8KVVt0PPKN/3/eSeWnIboGzpheWVJg99mPhL4jbqFmzF4SQTd1DU14bP3tTwwdDdzfMBT
6263bPDgK9tloelbcoc1BTvzhNiyftYAmgOnY56DShJcQngwJzuYKXnweJIBQDOYpS+w6F+4Hfgo
WbHlDohzK0YsTqcPpdqbHPgForCFCnpJBo8Aej0hPkfOIKCAVO4beHmZYkpIsWJZMsYYIPjrEOpL
SSlMa1PEht2ZO39TawOnjPQSUZnEyuYYs6tgriptoTBzb8Ov7rj9/iVSbOnPzMX5cnNYmALPkd89
kPjPMMXkXNQw1e7czoO2KUkAOyAQeNXIK0/0bgSu8WDeCYNnuEBL0OIo5vWBJiVppHcO4dPEW450
YWusP88ZVkYbsH1uqmxEL7fr46wlBAvQCy0gevWaJAP/qSEjoMSISx339+IbriadFDUWNbPA614Q
XieaVngpj++K/C/0Ztj3cwG2C8ndhQb1jEyFa5J/MMmdbmCnq8fE7zgcsujET1BF6aW5q4jYi676
I5xjvk9Qt9H/THRtJ28sBIpqbBXP+7vIIgHbs5s75UbplFOSXtj+GaNMW+/j8GC+CHQDDB6bMwww
4Ni0n0LioARK+FGypaDUGhK/NyCeiJFVK9HDT7MSSM97z6r5JSXe13Ps2i2hxk3zSQeU2HXayg9B
km27WGwPT7eqoGCWhZODBh1RWkRDv3sLMP/6aIY+q7wgL9qJgH6FZMBnb1BfbndJ3idmcRFU92k3
TKwsCWV+6klJOZZ+z/gJjcJOSnFGEGHxd84YFXjJRi19FLc/oPgsCl+AbZ+eyGyHXCDqjKQc7z0x
0hZ7JueDXq/DZJQJcBOotvjFZo3C7wOI7mv6vppB4EnpQFy67a7w9ufYOseFKklNoPIk1LDp727G
FLrd/zUskZom0neLs38hKiABfSKpXqAAFjeDfgyrEeqZ+cudG8nuNBPw+0FzrQhyqqrx/JRqywCZ
YcU1dkkN6qMeSj3VSXWkY3XBXrF9/meiI5O9e3A/FwdmTz/Sw4T7yklA8VulYspIvXPwpPCJcRO3
Gj6+fw+f51Lm+bxsYfzOyhYB4JMPhbRSKKphjzgLbZB1cHWhsUZ3MKgXWKtKc9thxpdxI+/cUJFn
kMGKoznbrsm5jywj714PvruMG9EXS5MYCR7DcbLegH3Hu9kEIIIkal66SvxCIYTVKMkRyl1ss2UV
n9O/4fraZWXe1c3OEW9GGPCDyBDH8/tfToYF+waaoYrp9XlyUmgl9+IjRs6xXZO+hTkjPsRwvOAJ
IxwQ/HRM7CvNMxb+1q2wJ17xKCQ0mAh4PYdVRbf7flNeh14YHIBn8f6SzQ9gxg/8pcBGJld8Jy2u
g8STr/1aQMEucvp3TUbxhCZhQkksyzST+Yf+cp+3hLV3+dY2wO2caeYWYMRB0dXYlkSYqGB4Ju5m
JwECVI+eT+eynC7q33vYiEYziC48rw7gDeDtmYR/b9wcTj/UOqe6F2gUh7Gy4MH4UCgln/1OvAXs
1nzqSXcOG5FJPq4I/rWO2GImYAzxPfzQ37DAa0EU+WBNuE4eGJlMCCsLB6qRqXmr4k4xxRjgTNlS
y8dirL15CyS4DbKqAQFyO5Dqp7fX7JZLydKbJ9IyamD88umQOpCp8ghYcZvLF0qD9aFQMVjLXFOB
QhDON78tH0g3atTnedk/fBqO+xIyyC0SuQrUVGRsqkimkity1QU2aPRXCPTkvP9qHWQxOy/mj3hM
kaPu/mskzw+8PZGcmvLnNJsBo+F+EJB+YBO2EZSEa5wLO5MUST5yotHOM7YHE7HI2pJXSPOfZL/R
awFXOVRp0RhjBJGWiqXg0L08T0NE4ctXkepnjzulUC3u4rTVzOhhTSzBBFZijA6+ftF+XmrZY3Aa
ZeP/RC0vIH0hpqJpNt87v4l06jtG7lv/s6CxRrvgkzFr7cXScdA8A55kEbAamDlyjqZPZ7Hxbk4P
G5A2o6foXDOrUR7x3fyuO7LL19754QHOrHmzOvBfzK1Gk+OzzbFIp9X3ZkuhN6hLp8uu5kjYxkJz
1/8Y5nMksIi1NozR8wwWK9BEaeJA4XupVkz86LQ8kq5TAmCYeMHo5w7exEV80XG/Zub+i4tl6Dam
gSNfnNMB6L+ko0fxko5r4/oqaeDzR2FgkZedG3Bh+9Kwfu0NM+nUT0YIlFDJnexcjDz9TvqHua8d
hZoHfrGv676fV5PEIf0qZFFCAJGZnQOGTY8IUipIHFvn/RH77ju6q+Gf/gC/QN1+Q3EXa7n2HLuo
v8qDFQ+qyuxwv/6GZxajDikhhwcQNkeOuSEvjLAUjv7D5ggcIcg9yJHfq+e1DurSCZAr1X71eg7F
riSLKN+924ns214JDbR5VZwYQNiDMbDW/C+HY6sW9BwxuA6A8Xp6MOLjthjB8JYJRKwZmUU0PlJy
10pjfTOSJa/JYXLPcsFl1hxLqndk09NFyG+nb6fOpo3PQIaH+ReKBnSJFaVQjAg3W/Wgqg2Gxar1
OhQxfXwGG/tdLQZ2lm/nF4E3rHUqg8L4Je1NeIo9pF91r4qBDy/03KNgcIFvIZQ4sLaRnjt4J9q1
vKD6Yc+m1rLrT2k6sZjEaaWh6mdwZ8fgJ4ephPr8IAH0+LSnQ7goZQFmD99RedneeaaJld/HeUbl
NHHsIVzHqJGfrcydSlyQeLX0wiGi1ACeASA2thF2obW+vvPDovMlZn0pP13Xzo4XZ/mzUa1eC4mc
d3e302pQtjwjezEtJuq4D+BjFNgEYZnd3Jf5+R3FoZezLHMkQ3LgtsdHls1s4XXWbm36fpr38EE4
7H1Fru2UI0In58Vh3Y15jaMcZVMm2ybvyfAOoMdILYLyYg3kYFAxogHN+t5bdIAu5pYjak1Xjw+f
r9qGJtsfI/LGYtNSx5zu9MkFfjxxIWcd0TB0ZNlNQ+vlmlXA1iZ62+u5JjWXQ9FZODFV6sFJ7Hc/
F7YduxIi5wOVYwFRwN3NIr614ngn9JP5grNmljJcv5cTz09JOOduSJiHn8ktkhYfoxfCEUXztss3
iRoNyT8w9JIYjZbj9pm5G88S8xr3g5k9RK2UdbetHnYEK/OeaJ/5UKzOQa9bZEx4JecFHSK+EbfR
cm1Y263aLapkh110bGLZRI9JtvgPzpZq9fHTIQlC0S+OqZF30t5PKKI08BU1XQHL6NeG1AYaFUZy
M5qZJMZmUhRsDI38wDaKWG+yCeyiWA7/SWT8f913STOd+b4ememCXSQUZX6tTg6roYtKZAxoCp61
/HBUIljuD9+bBBhlue1AbBS8DoCMOSBn7W5/GdxmIuu8lHdSJtje8KG6PT6mpS7uQJxdHnA0yid5
Vqx3OKMrUdliiAA5vFt4zml6E6aLAaqObyX4gvYhRzQSdnwc3rWb7Mspm5PM1cARQjOaLj6RsOYs
8CmniohMlqZDGXLJXdhYoWNEmNN40NiT99hDtjiIOFEKvu0dAQh2zUGyLKGUlIV8wTlu9OefSR4W
riXsbgM2nixeelNStCcblXEkd5yTL/sP3ZtkkvuFLIkxXRBp31xMiWC6FBt685Qm3z6hqOl5tE0q
R2JbNqWch6TtUBcVsvxjC/ox4HtqUxtmajWj/QY3KKdwUVtO6x2Bsy0wKvE2/YDZ+++iVyJ/183u
1wSjj8zMIppMtI49hwThoLI8AF+bCLaKQ5dzY7yeMp75VC6RZ2f5vl35lRuI9A609Ed52GBjzLoB
OYaQDwcBItoOAL0EFJfUODyoGnlaHpGUgbRx6nRs4pRm69u2Oryl+bUFaq37+IK/UYlBG5Jka+cY
D61xtaPs8RvnGzy9TvelanxVUML4VjTXEp0dBriimpwBrrnXtIPXDcwq6o+Hd8kMl5L/iMeoAap9
gP3ucedKIdiAwdY/JnSGX5FOg5NLrpJlpv67c/2oybKBZwFumsp2rJv4XOlFq2RlBhhqE5rhOYey
KxlOuRcbMaLit5u1tIZsKnJXGS+oCTLRbbWYVjJWDf+EkDSZQwSBO5lCaBs9FvcONPpjFtAj29mi
MhQr2C/RDBbkpFfm3DlVYxzTkcIhh8Gf08gM0zX0gF5BiDxI2dTX7IjrJiHJdvySH2T2uKTraWtE
Xuhm5YIkERVLzJCQeY60hPo+7zxTJmVfAwYi1cYuszhKYVoXPCvu7Om2rqc4nKNeEfEv75Hy3Gz1
jhenvTaBV8HEMhYnev6BVaTaPcbV8qVZxdtq1DVsOqU43G255G0lWexqgW+cZcYpMR+UCupamaZG
PbJhSTVuXU+NggxYkNXA+VstoKixjOsK+hTe+erxE+c1acjzqkKuAaJPCYkrphOarTfbxztNBeWJ
a7LYRm5P2UyVedJgWJNv8vpD8U02/9xeYov9jpEF3gfnlFrZUCAdShG8ApAatPnWydtj38Ao7PtF
XM3kECJXsJHV4d8pMrzBbNu7EJARZjUSSpDeCSR1SVrkEUAfNxhLywTlZkWvVt0+xTNAvdFIWOaz
3KCCJ/aKTw2lLzaNZ6bBWrHZEKlH/g25TB9mJ4NsBug0F6DWeK2ynj4rEGhC7k+m6FZFxqo37xDP
y+MmvtsqSc0rdmJxGSvXoUE7a814erjpK/ogjvODoqDfUSUQ4DeH/pz0DhD8jg/hnmwqqQ8ie1eE
6kl/jb5jPamsrLSyvWAYp++jom6nezrI/lbvXztG2gOJWFIwb9lSn/+7DJYGZ/uKpo0LH9CZpvMv
yUdhT9uIfNh6EoR90YVy+OQ4zr2XpoRUGJDENOCTM+Z3l0vvlU9ae3rlh7VESjXdn3wglrNNNSN2
akjwMwmcssvqHqyOA8oYwPOkiYmMv6hchh7qDLfE3+jYQnXTly9toCvtl5CizjbiGFF5uMSr3bXB
k/dpjBRUJ3hnECPA3nHxHH2JmjXsllzJvXojJ9mopvJXIUKbuL0BNGoxYRSDuZ6wBM4VtvAOVKDG
pyjbu+fDBbKeO0FO1WOYSBZbm8iDJ36VaAXNiOIwBFAl25MaK3TFIrt3nzQswfMDskyxl0i2Gl2X
URRQ7Y6vTxer7Xc2iOtFD50Bzt0AxxJVNJP1BX+2D0/Xmv7JBJVOQjAuKPCtyjgGfg/fuQoKqZER
3ZaiSYxpUo1npKL6X7bFKIMs9N7VzsJ2JIs25HMm0SR2mwPadx0velWPNOLA/jhDjrO+TvzIHpUo
8ULBfqH2hQYfBsER8DHQoHS0RVUQfje5iHeDL9eHO/xFHgmAttvFkOoagNnP9R6R+InoYQ/Nm1jM
fOL17UWD2buPn06yIuXzLbhv4ds7VJ6TJ9yyTQT+gUtL1nH74zULw+U/24SWappoC//Jacq8ilbl
OU6oHCXIz3jrjYMmYoiJFT01lkZN57BjptEjhlVzWE/UzwZ1BgvkrV1r/rZQiUQuVrgTPpiehjrD
P9TFrIUoazz6HQMQKAVIm1cvm3RtMtrSB1SvfqsBgsBLwoqHhTfWx+01j+C4rVpffwCKXffShuzC
FwIgyCwbd5sEoupGKAfpt7fTJh1pzKhjC0bg5BUirL8qVcmKc/EKpOGMwEZKx4Lygg6tLpzsEt2y
HpgMvXBLyChG708SKjEb7cPc+gcXs/Z3GYz4y+C1cHED0BdVVyxWnDWB2XcgDUv1+fVKDiQpbK7o
/gE4XdVzrJ8m8v4VNQKu3bd/Opisrk7HqHzLt7wg8Z61X2lPMPVq4AnicK/7rmWnbwiKtq55xoEW
ZY3pxewAvvs0jRcZEPzoYG5z75T2PxFpZIGgJMEw4eD+dWnQ63zUs1QGVcRiFNm25LiFzaulitk0
hVgaUmJzSBkMt7Sf3oC3dS9zEb58lO5rKuwF3dOL8aaRRtF2eb3frBCaJu8iQZIiexpAoznWpAjk
f9aFq6W22GZm1YcKMB4QTg+9nx/iUKo8aZPmkqZMfdSmbw5lY8I0WeCrFEBi4wTfFNTm9WZhV/7+
Qf/qPKYKEZtr/5wxAj+c2/G2jWVPWarCUcjDjFLWjeTd69dOONAM9D7Zdab5dRnHM+9cSZAcWh/Z
5c/lKnOcxs/y835AFCxbZukH8ahcDLwttg/IroaQz6DKDdRtqctX+uwOjlG2pEIT192BRJ3y1DKt
Vc87DZWiKqmYr9rmDhzPUNgJpY/YoYsSGc6hDu+yo6Ibd/KZMuyEPK5ZLis3Ht4dbXgp2KxDtqSU
jREqh7jCxgZbd/uKOvmzQzm6gDhGMDEJ0o+cA9kXINmijTeR1QyzOej6Ty0Q1EU8ehKhsQQpC8TM
KPYLPs2SVM2boV+PWimEzjSOVK2aFj1mW94FeKKeHQ/k5Vnh9WfrhA4C1h2zxqMTpmhfftic7Tan
JKyX/qf09ISJ+3vITDbqT0C+KlaJ3hh819dXe21H0PRMgk/alexUHy7fqG44gbKrVNViPdvY6xK3
nY+0zOk+V1lctynmplixpwR13OsCaZrBhlnrQnJ1emyES9+8+IWThb4L9O1z74sQqxguYZY3OgJ6
WZJ5dozvJiBlZ5PKqGxLXf0UyPP97k1rruXu2P0hCl3WaQO6s3jv4ZDCigFAGX5YTxSBFFcXr9wK
cP+zw/3OzHVs2miLm/oOY+J0pM86sOJNa57xNytavi/gGPjzCd736I4zIYdLH1HlYDy3+FSn8tdk
KDPgIw5DNAbWrhTy6Umr27TBqStJcMz/9hhixioSeQbXLIFrAhyaVGGL4sA5jGmA4rWkNk64tyZa
kVteI3G5ju+afN+DAapfmcs4MIOjKteH3PYvakpIG96xpHJopleqoxlxml65dcoTnwkumZVZjJBF
HJpno/eX04gduaAzsbubPC3PN0XSde/RuMBZlh72YWYjWbrt561dlScN/lQg/mz5VJrVM5EHXB0a
7xTnn+MSInyiCXQzOqYm5v7hxlQRglrFKXEmrJTGAvHBMZLvRmlqgiDRiy45j1GN8k2miSZWoqPh
6FonnT/bDO8Nf1URh90nubkn7ZAhA883vteCnlMB/MGpXDhtMrtV6CmH1G7b4f2e427qRy14ylL9
8VtPgAet9HzMVnzqV9VG5LkeXZLS2tBMlCM/CHy8NYnXziKl7hzqDKfrnUWypbU7murl5pdQF3cL
HT+Y9tXL9V9H60JKYbA9091VQFRE8L0cP9kzesdAaeuZ1xJcuoizPcbf7MJVMkts93EP10YobG+T
WYeJnwGXKqI5ssT7vDzx8qpGpO1KLuXxuuQHJfBDo8SQ1SqMCMJGyT2+SULllLXPvx2BWDHp1Iip
VnLB+US5mj3PIAZe+g34hzNHgiJ1Ukc33E2BMjej4jPaEpqelyMvYdEtt4pRn+PX8kanWxeiYZBg
0BvnB/UO5/8B5NTnIpNFlAEGorN0DsycHKAol3A6oYUOvnsWgNCtk7rkpGxhK4X2aibs+avwONOg
06thGtVuPkiDuwiPEJsmJe2oNMfXzr5JLOpjS2lAmt24mvMW6GC3djMqZx3XjGToDO9FyNLJKUI3
XJdmJNirSswd/qLgFWS0a/G05Lmo6DJsRsD5xGH9pZw96Q+5Zm49zlVeKg/DiJQf21DvILF49HKT
EPlWK/44ahP8aL8pSzby0kKVXfIG0Dwla8tlOatkzdPq8XcxyE8jjClqRz0n6rv1ldLI2wLG3Brh
WyWfweIPTCmHbWPKshDMi/UeHtbE9QX0nPwr0mwFk8qMWHze2GcxA7dyvJ+Z+3y1XX/3Ld+0kVVC
ZXu08s7eWx0k/BLlAepU1nsvj9BC8T/PtBVAl41h8ZKFLLjOsFGXU3vd4i6vC1csqkqahQm9xBmo
usOrK6PjC8yM5Iuiv9t8BeWbeok4nMzurb4/BlekZK6Gf9WMMjSybrrJl5UFsYajdVjm0RCA8FQV
+h9WLMrS/5TIZPxwcqorTf/JGmQpMO09RNpCcig22BA2MSbl/qxIRAps8dTOvMNsZBrpTClvSVo6
TteCLoFJaTBDXgijB3oGNPpNLMPrEcYwZzRIryj9CJTYDhlqY1UcLxHn+iHGNoOt+N6rQnn6sos8
2UfGE6LDpbn+708QFaPfL9vBIf++/OPxpg4Qbrzcjnw/uRH/GuF3lVde64aQ1IQHOx3gQY0OVUI4
1qjWcAIC2Ju4lxfAA8y0OPsZJBnBtleWw4rYazoyMc/i5nrh1pCsYvodRPfyFn7rJcxJ6arpVyOi
DsHMDbI3egUpgjYUuz1Tx69mjjxfO3EGEPDICxZOq/ujWrA3fyCKPqB4V0meegWKVvq+RAGuAkNk
481dNJvWAixFnW2J35upgf+VmCjyypHSAFgoju/8SGOVngM3rezMD7uUhwyy2dh0cOulitK397J3
LnMHpEs2BvBOm9U/m4WeIexZebCD3AofUBykCnNldk8wncJLXTbYB/gNduyA1eN4scZ1Owv3HsSZ
k95CiXofEWBazRjAmrHuWPRMdOg2/HxtHf8HF8CNxyE5p130rN4FGSEKNCIbo+oiS/SDCdhhOEwz
NAdEbKf7mO7wm4iZa3a1o40UL2AlZkTf8lsqqRsktpgXCnMQvTVEfPYiukOl3yBLo4JMmg/46vpU
dEfV93lj4qYOvYYWLgze5h3SI8Q5yXtQcBLFS1/OoARPM8c9PIRUZQ196Lakos7ni/wNtGFsQg4n
tib6bWOAFCPimwYIGKQBW4in/0nhx/3vt8hRuWkhrOQ6B9RltfhX0KVh5y+no/jXNj3mr4TElhK8
TApfFGt8mVIIuWqT0O/2vAOmRHwZx14FNgqiq7dyeKljWeDqecgP9ug18kJOJO9LFomGQt10vtJW
Ts2VCggjIe+LrVesUhZa/sVZ73s7ErsJ/r2gC1WmFbFoKM+F0fUwNmAyEqr+HhINNJNPQhk+/FyX
a/GLUoIVt08MApFprSPSZ20lATVJxxGqTtAsC56vrKA2HoK+fur967jQSQlQ5oaKifyGslO8669J
36NfMyJ5OqcqrUb8ovgMj11QbTpR0zkMdLwMsVIe0YnYJzIL354CyoV6ipbJJSyXCT6V9DcI5C1q
MWII5S0z5BJT7VZ2SHXlTpFgBxSW3tdw1pzvaJJvWSqGG6i8F2NPAhaHrmPCYbB10V2/n54o+yIm
EWWMoK6c3gYtM1Gwavnz+QwIgLQuJE0IUXiiKDEoXDGFflfKyIy9ALhhGfQez4Y2HbGE0CsaCx+x
gpalKwGJ+tT9BI5b8cdDXaeP0H8/58awk7Vx+xv8Aq4wKRl8PM9Tr4xfwz4kosEif2BhCb5dv3/W
IXI9cvyxkm+2bdBC9V1OtcPFTHd/wTyX1bZFFhDbsbiL/Nt/5wcpQLtjk+NbxWBBdSF59sCgyfoz
sTEGqZVwZYG0ojB/KzUffyVAqxgSOokXYrEW4atBNLQBxzLXr5qhj/nexUWxjho/NRaTq/ohZOOJ
ItI7Byh63qTGy3E6iY1EM0geCkb9DHa/AVsZFH68pPsFB8Oieu3O1YUuWi1gzfiGEw7Ta3dbD/rO
ls6Y6V7LPA5Ny5Iclew1fCf9/zZnENK5WoA4DGGRmfHi5VL3IF6sSEK+vWRnRBERecYQXAi+q60w
da2diBFEnjhzu6iQ2kky+WNepZUbIuN0aA8HB/5A3o33pmhjX6JKsWjfKFgV9jFwPG/XwjvWOV7r
WPYBf3sW2E4G3FOWEUcyJWqrpUD0eOh4+hPGCDnXa8BvSjvSVh7yk4/RhfVlWkPbjlFn77s+TQO3
VifYMfsCcRAuQja9aKCXihy9XM+rvvq709zLGv1fY+OLKxyiXkByeOSjwiUXgQq4BUs57c5A8/F7
xDx9rRbu+PkNN83BKnTj9XIfgLrZl9qSpPrvVeQskybHZvsVoUzetpQ7Zzt3CIGVMnkj3BS+pioA
btGaf4ozO2o8fsHIbCgSUz9TAsuYdwm4mRkqHNQ3OSiucOxMUtafFJ9tAqvGPyIuWaYVkSwiVVhO
d0pSOSe6Il/BCBNE/EwgyraGadueEsPoyHTJfnwa9E++25toCXeipJrx2HADnQjDHlLp/xEhVemx
exSfDg5qRO/jfhQksNDf67z2ddGMYH0L83np/RFCGKj2abmVoAvP+m3u5yHKFYc/VK48xFf5TfJf
7zZpr6sV9xMKAAk1YnOa90GDU8cWCVBRle94bX8Au3+ROXh1no0zApjkbhabQNRlyF205ypn+HgV
6gVy+5OV+vqi7GFVA99Snjyws5W5ukQMI97SgncucnfhDyGbbCD/58Keh+hSbGcd9GCziv6qUhUr
43oKp+uePUqln1wjzSfo221MV1zJhY97reUyWpXBhxsQ4J6EBcyAetqwxyE7POKJbH2xacBZlJsM
vMvX3IFhib5Tlluibzq98c5Ks5D5Zatqjd3KqJuS4uRUDOiZWePpWHh4/+droLveeGzkJrFv77Sl
J58G4PQkJ5DJ/chtVIv+Y8MlFJJUmoxkulgiQHZ+JraMGE7tDdeiZt57d5Ywr809x4IJ39BDYNoI
9dTzXh1LanEl9bwPapszHB5zoqiczdx4rDuwfLC2xQeBxrp/U7UwUh5VHJOJl2jyQduAw8vJeeOv
0ik1U87gOo5yiKAjTHNc96qvOboDoVs1nzun0mfnaxQathn6DCWct0uBlH3ZTQFG6RfHWGnINnl3
ebXaA8XjQqE8skJS/oBr5KeysjZkivW+t/HKCupQ+h9FNOaAHjYky8RdtFRCukbZdBbO+hHyMZJf
kEl4lAbQDm8jmXzTrmEYuoEOd3PKXsm/fWaRXoVFuFkxTqQhrzZM7GO0OkQaNe5x2NLQHWeoy1lQ
et1vECxcT0rkmmFh1YcO369BzvCF3fjLMYCjwrRVRMan0K6B6mDskYeKf3Di8IVFKI4DsUyXfXTx
WGuEpI6bSvIAqnf8VH/DVgdsynurav49KzoGw/y4bWHWIW+2vKzUhfh+syvb69yyB2Oh0sS9gbeY
0X0zCwIjxI3Q+qWQAh2j75ZfUnpv/0xEdUvp4tHBqh/V8DMxzIQ+f/eoYKX8hdgtThwz+wL33gIJ
+9ueu28BiZlVzZl4Kc+KgEDub67dR1gq1dreOutXy8idMViPqC3uvM1Z4PrQNjl/53gxmYp+uoEF
9c4+/x61UVFpmCg/2PAYcmrlaFvd4rTEYn8Da+HdGL8Ma5FhWUhlqlCsteGvRj8LOdBwxm6RzWK4
BuB67EKMoyjnwSsxtLQO3ILgiqakAAndFlrVxqYJwt1Xt0PA4JTNORI84zCNC9KhUbDc1/4gA9oF
YVLU97hrCJpTJ0azK01Dzi/vMwi98PQzWlugqYDw71WGcznOQTwt/W2lXI5QIxdA4LSU/xmuS8Xu
FmYPk9zHXQUzv3nYFpfR77tTG7dof93MfxZh1gW7rB4I6NCHLcKDnjsit98zcz5NpzoOpZVTEIyN
dBu2FFbyqADJ/N1qCi4JRKokiDTMHdIhbFtR4cz3KEDKUBmyqxQ0tMZZceGW7q3bFKzm/z+XFoje
4V8SazJ7Rv+EK/phNbxTe8U4rSywqmrjTeRiCEiKJ5HZyuKitJ1P0ttS+fNnD6JLZd/8XgsKob7k
uv939ejfPiAwl0xoG6DFqF/578NDuASaxMNr8SDKcQMENxvoXZzIZFxGYmjlY3HeUvrPYmx+jWWu
aoAy+b75jLSZf1SIa8mhrS3l7C+jApLEU7YV4cS8BrRIjvvooaOy034mNTd20ms00JJmk4lUJZpk
2OQnsOIOzmgoA6Ei9gpmpZcA5UqdU8E+a/wdEzYOuuHfakoOZ4zc7z5Rbs1u2Qd0jFzT2CnTHjIY
jGgPssJccH77qRcHqOzpZcrXsKBDO40sVvX4yF1xh36PEj4wJMHpWlL/7n6QsKq+BJIRhJOzdM7i
zfZr//ACcHA3yZsQE0w83DLFcIvBE5CHjmlp4JdLjEChZitpqhkNXrCjj2GYilSI//HADUVZ+uhw
T6IfKVlsiKJsXFBeUo80DkuTL2towVZpTq+15t+LihOamh2S8+B7UM9nv5RToFCcBWo2BI5yKoaq
RGfFWHDXBrqQ5gs1ME5w+XTTegchTfBJR7mV1B2VUySfGAwuzsuhJqtcXIwNpJd0v4XyV+d1iS25
MO45/YbX1cdgHRrLcFifNaiBHY2CVl9oZ08M0vbyWioiJMZKUnt02vpyJYKeS7mNGDRTzsr4Qgib
iYetDR0wZ9bCQgf0v4J6OYYMyuD+6dlqpMxqVDkzCz1oku06M/eG1r6IVJCL1vnTHwjKkJFdvnqC
4knOPstIpdG9MNUIBOZlFwpz/Mqj/rTdMT1QwqLRAvW4tE9lXIn4NH6WxiM9shqEKN+zlWYHfz6V
Gx9moGtAmzzMbNTA3edkKaVpCaZhnfb/ny+epgl6EOkZN64nlJ5THgI3HehoWKFWWNc1Y4GCMjKW
9EnHki8mVBbQ/2ci3Y0W7zZ7b4b0m7QILz44bDMidD/jsfEL1cQxjoSp4Tg9Gd2UWRLKD7Ijc7RO
i9MLXpOdzFRfrIMdbbVkss9iNTdPpPywYIgmLBBuWglQjNjxvbmR26jCzecVYoZMLo4IIb/RdtiL
52AcbwYuf4ZNGfFO5yRfAf2FzIyDQsOE8BBDNLMWEL3v9ossu4KeSSDXcWTKKmWcEO3fbzJ4Yia6
8Ohl9jxavPxMydmLz6dwGQvV5QCDGlbL/Rl4xPfjkQbToJ/OhgHzPgDVyGEai2zJB+DeWd8QjvLd
HuRWDiEvpUbF/Q4yyyc3WKRsN2JL6JgV6O+TNIZjZ7ku/M0ZJLwrTfVFlXVUOYTXda2WXJQUbprw
VfMSwFUpwZnTy4vKrkTgOPGQx0eqWPDj4Mo92fXujed4pdlIhwgUKmtdHbFyDr9Ht7U6GS49ityW
0FAmKfeBIVZrhROeyUxpT1AVRzqRg1ZafRLNi3JBbwuemAY7H4lFig3IGq6cbbTGMGXAVU2GS308
g385Me+eNoSVdUXYExTVA7Sgq8YRI9dLrA9SUbKj/FmGQQXDlrW8HXUvqMDO6VUcSlRcIeDQbOPP
oez9q9KhZWA3MYgDwUh+9dZUVf+aiBZ2L7+zsWVK3w1z7iU6hzCCD2Scbb6RtXwQyLawl2Z0rTNy
AfkkLwi9O9qAPCb3/Wrfgwf1vu1+LdbkjytXAmeI0ABw8Za3F/ZFa3/b7HlK/aUbdYi1+7qr+H8T
iKu6MzpaFBNbfZBQhbMAXXaiaT7441Z06irL4hD1oD8fso7rShwYhb4DWGvJ8A/w0bxZSSwTCpye
K0gOpzb2kG6HaFa+k36TAesDN7ZR87L3BDhT7cTtXSRW+udLBMdi8oSwdSidKteX5VB7hRJ+R1LI
GeDPU/POgNNTvejxqc7giB3McTGvOq8uyVRN7P5fHSmPV1V0ge1XSxxwY+FRyZzDxPCcVue1m+rc
v6ugT5Pb/kBuv7ZlpBU86vmKKTiR+0QfMSIFn53ZTnqDTlk7RPKrx7cA4Vz0o/MJmFHzYm8Wd0D3
BKNnN5UrjZMeBFXOfSy3y7XsFMBZvIouvX3RFpw1cucHV0h4G4uPDbZO5mXiLnOsk6Nlg60Ci6fJ
4g9ZOBPS30G0UJxAwdtfRJrH4+iXAqq4t4HOXodQdc65TWIK+esHiWRkoePgxychccDiR+ZavEyl
Fvk9ugHHq+qHvEOmdXQXHch50nkY97HOV6Cuqpoy+npeQBCnPVIBsV0jpGFcVvt2wkMB9ckKPPVG
h+UaHVlXJ7RwlmG2oyIES/FFwec1AKuIZcsoxetESBCEMovrDD0V1P6nzOR6dVC/hTs470soQHc9
qlIZl3vqjc5Jwv4vUz/VYQToi6+wxcohGCRlMvmsQvoiI9dvb2S55Xu0t1840HpNaxT/RCyLfYcF
f2Jr2ecpZMwcv+HUa87r3dD8Kp/I1lpKOEOfomSW0kX8l2NVxhrhMWn7vyXSc1ewU12htUFbc11E
QkgiOSwXGAS9ohO3xc0xsfuPERhW/52u7yMMyIX63EEysfsuPt1d7Nh0q+DbmvEnS80FwNtQqDNi
j7fxLtDXGYCtn+W6of53CjIJYJ/MleF5AIDUxAR8bHFU2MHO15hcriCnY+FEunw82OOTYNq6qhhy
letWYdagu1uZ1fOSooVEjth+JgDFWALvfhH3TVSPW7ehihe6R8SXFKTY7bd1sddauFV157PUt3Xh
ANUkDAdsCHmtvgB5A5d+xXVIwLwQGVV0mKVb2CwE1DJ83ub0AdKElstk512wKGdJucyLANmJ+Eb3
CRIYA21ZSsh02q0GMPB55SSm0UhJrEqcpA4u1marCBKSvk6W9QDYeVGxuznFU4DulEOEi4+Oo+38
iqZZ4MzjsgM8PnroMBQqJs5PFU5VHeHfB+sxm4ReymbXanjVgm0+8oacljm4ImX7Wj3sbaBIYFg3
ap/6BGpte+yZl8XLP4kQdLIl3czy322+VsXwq4AxluXexYsDPkY9EwurS62ONxdG1qNRGPqIvZiv
UJrfptblQhi/7nIe6cI6xQdxSgRkm8H8mW09WnzXI2w3djB4eu4PxPMg1kEeAMp96ukpIuwGkyNo
ooouxlEKnZ3KLQ+e8N47LQCcGo2hYG6LpRKJwpzyvYwCqiQ0ksj5iYujHPPq9y+ahVTZ+Ak3pjS2
1ZpG7K3dyw0MRrX+Q4ZRcufVJ1P2zJuObetmzLK9PKLwyfpotMFNW+nbWey69tJyKQD4A0suAAxy
VJlkCQHg87YtGuUCjwQNWSo+P0QHX7qN1Zkr/j6T7V6xLBU/aGvfTenj0/61BoJHUu6Y3Y+//Nyg
C84Wc4W+vCtPFTzujJhpJ0F49HQeuSRmed+0DxHVOnfVwy89a5xSGCcu1vzpTWIaYXayHUVa4lP6
M04RtvLE524vJhZ3MGJzsO94LdexA2sbkIrfBJu0gJIKHl64QacTbc87hoXWn2X9X0xRAGEKuJfS
yhY5o6nI7BqsHumffGcE9pZi6HTgT/5iNKzXPDJdIAH4k5lVbGEdhJRa7SopyqM1b8lcMMHAr8vG
vc8fOAs3/2FM/ZudFxaYBezwGjFZVVos2Hd+4i9pxfpyrFhED3uK5EF+7Dh5gaelWCDgI49gmoTh
Fk0vQ3z54yX5zcerSVk1pVzhGpPsgt+FPmwXgGrJDzO747i6iSpa4a8FpFzy6VVzR/mhLRbikuh4
urQdYGIzckaWdZe5KXRq+03J+z5gVTrN/feQSh1s1cGBMlYAiaLDpiCna8YWb/4IDnsPGD62304w
PQ6d7+7mzCfW3Nr92VeehYENKI39KoTxoePqK7PHxOuXpcnCyBAuB/3XPDRtg1kdVDf8gfdvgWIi
wm2Z2DNNpzebBDd+tFTn8w0SLs6giq2/c2hzO+n7qV/IA2dDbCPgcuHCQ7MwPsuGaFBc5aRCZ9al
9QkEed3xZbUZUpiA4OzpSi6TLob4gmd3cOgZneKQr6T6+IXZz2sv0xXyqgwq5ofEh3L71a/NehWS
yZRsfFsHEEypXX0yl5VpQd3QyUFHtMspGK4ETE6OreW06EfBco5XPQqjTNz+8dBjz0yoMJSMwHKp
lbAULVjQClFM8wI6NCmIpJLN3BFxJnU6680H8o/tTAGVu+OjV0MVTkAfuFZknJRVx2Im60m6ulea
hep2RBlgZ5KbpScdFBQLN8IbIr9dc5J+H+TE5fjhLWvDzXf85Rz8MxofLV+vBd2ig0j+Ct9kK63/
Mj+8BUhrp/a2NUnDHuO5YtNjTUcD4XMiP7RhgfscxZEYeP2fv6DsH8fXrJ4T8ZAn/tDh20TELIQq
WUKIpnA3eDVICsa9TFz89Jpth58jIJe2GGHXWaKnVJOQRqTb6lSu77li0Hp6lXF99tVU0e9tZJgl
L25XZdlBj835mLZ29hNGElZVJ8S+oYb++KcDRlY9mW4amms+ApmUnggdylyqZvAc7s2SfMwHLmR1
RWlxt7C62e5z7xx7l3rTT3gCb9wix58/kK8eyGM09NGYltXHCW7oBP/2MIjdt5ui9SKBHkHNlDB4
zSsSoqQ25pJeMjU/EzsceX5RQ85o/h/5W3Sdw1UX1Zrty015MZySB+DpP1e9kByhF5QUoIpjvAN9
3FSlfTpb+GEOxP5IdWAZQKc4CBnhKrr0kzW/+KTlo3J3q6GHr2yY0eQ4wY7FngGKkJDImAOWJahD
qPeMqKkvf3BieSjdWTjRnQervqlQpsbC+LRujxrPlV6mMqTi+fdJDdQRHEXDWNjgDnyQ971N/VOv
ZUog92ksB4UqsO/oGGKPWSay+JCmldjIBA/NsAZb4vWQ4rHMi5vmuwN4CZOth6MCGtj47vNniGle
Iz8tdRiWhM5rCzjnvpiV+HnfO6HlBPAAow7V00f7rbHecirbEHM06XFwlGkjdvPcE6RP09wkMhLu
ZvMJb7C/y95WMKnZ/wV1oOap56iCghC7XJTisRp9kcWDXj0ARFpwIJmB+ON7b75rHXTBTGIb0OJF
JOAAFQXyVHh3D+lxZiwf6Ms6U4iF93yiQqNJt4Qxy2g3BlksvlvFScKoA6z4bEigbU3peiTB/wWE
OJkuPTUCtPv6bc7MNcMDxctaxHJUEI+JopD+tuivuKnlBn2NlfFZmCWJ5IqNRUqaDjIWVM0hmeap
QeRDtDKluQAIe/SB4904e21LHEKpVHNtLiCKsMTLy7P1jacAryxoxl0sAAavfNHFzbIC2Q+e3OZL
27DYikqVkoFy632GMqkTvtIi6fkrakumH3ZMA3ADG75gu6yzUNuuVFeR4FKTpCxdCYf/wxwXTSL4
OPmegH1zeqqRoBOeWqW3uGXUtUo8OU1nENUyHyvro29pP1Q2zrYlD+T8genEGR0Iv7KbnUua6mdS
MCS8IdYBNMnNOZfJjqNuRPCcYukhIwSJ255T5mfKgr3WO6mQ59ot5Gthq6+KBxeLD+uat5PrUx+G
QV9L8Dx0KtaS8GP3Pzgm+E5e3LWMVrnz+wgiBBhk4PGZFuQAYWL+MjPb6Jyq8/XSplcaB3W4aHF3
DWJPu+8C0ZIjqoTwYTD41OMq5FLbc8Uw3+2/9CiZPy/3EHgC6u/Xh7o2mbdXA3w9hZiKLl4Xpy7z
iSssiAWv1OLXwR3Mno5dNH7Y1EdEICMit48XVa50TEStpi+/PMFK2PQfMrFttllS5Zho+ImkVOPE
eG3gZ7IiZZlbnwasl9sW0Rxqu2WYMJZLaRe+2Sc2c5fGOhfV858vkqPSgK9qN7+d0RDXQtETdPhs
21Aogz4dCpxFIbdCgmaPLRsbHkrQWNJUpf0/zptHLlkURRognsKjj1GJwDMfVfWBe4TAyEUvnUG/
W2BuTKCYrgUFicF0VwGFeifaRDPpIn164GFjoXRiF+taUnScDJYPNox0EW/PLvYLp7SWVAoVPO0j
NsDgf6i4F1SPkDoNcz0GAT+48jUEAMN5yDETLlQcwQuC11a5ttAbbEFCddlAkw3BRzdXO6yjYDQS
9+jjEklgCOshqZO9HTmBuZ3H6MoK4lzjEnXXTStbPIRPJ+QOKOVZ12YSPHUTZEAGdGUDYPn0khki
aTNWIOOM8QCgYOhxgv5cIKyHEiPWsEbF5L+yBj8FlMc7n1ee+DpFjUJ+z5pPuKngAYPGnLcqkStv
O6ZiNkx2ydxnZulRwGyQ4PKgyOnNzPCGrwqoTYkM3AI++ENQwoEqqDPJOWWPsxBMxholZ6m04pfC
+3PSDPQtXguGjpsDuQwjD/kVlcm/aKJlnko10TaFCSpUxQXmpPIAKg6fwkdpqzbYB8tqNz9KHG0B
ts47r+j/LCSWQq4xua97s2wXP88YY7mKNFZ8Zkh2953+ou/IyuI/BfPR+K2zOyA0J8lanypLqdDl
46jmRczD3hos8BDRT4G1cCA0KYLIzYXNv5g7pcM2EYsW3d9/qyfL78OlSdSt75VFtFVpBNtj90t4
UQEhNjerwg13x13vUAYzy7V0sgQ0ixLpISS/JD/eAhaGNEYNbOIVemywRGXzDnpW/pyx2uNyDLG4
3LwYVeVj2LPgFfua30BQ+vtATu9kGY/of9dVjM4rotUbiq832bt3KNsvbfeSQ4dMqAokxKQoBuR7
mdT8f+UQcfPYE+WJ00a24RBXxM3RIPs/GGZXQ/NNDntREqCA+iAoHPTH0GgnGplpM5h/RuK0FY5h
wBTURCDHm2Rahd8ryGG6UBkp3+HF7h+nxKkKWMjH9li5YEUTajYSCxASXR3oCjHcTVO1raJaGPED
rN4ofp+Zn/KwEVdwoAePdqBgR6J5Us/ehW4GvgE5/8cDvYB+G+9hBxS73heV9bulpPRPuM56WUZV
7fOfrv1I0Z972Rz2FMELRXtrkMr7YWZSjkJNkIfJuf/Bj4sZDKzshxMCEUB2gGqS3HPNJRvl4tCq
UDrZxy8wNCn+/4Jx3JW+q8NZrESLnqQirSnvcqEtGFAVfk4QjN+vhiu5hZbPUaox6kSXVO9bsmyI
uk5hMMqqFYrXPJdrqYk92DsPEsHC2GVdAVuqeC8w8hF4DAx+cBdf8xVdA3M1c6DWUTxEyS3+59c+
Udq3h+KBX2MsJbC9T3eYo98eVU+XM1oyYZ1gb8hHBms8vNyRGfnfvD00UsrlYzcG2sX6zyinIZe6
SMJJmcKph0JPlqgsJwkXRKsETDCEZEY5QxIUzLRsaB/k852SPJt1WqgIkvIB43MawKfWXbGLrFzg
LgE0vZjAGRy1qasxFI8dbrs5/osMwrGpLfPM70TnnjoLdHX4y6+rD2Nv4Ydlbje7Z10ogc9PXoLf
DXDAQkoSwJJ+IhafGIDS0nHyubFW0FNeDoWrmUQ0f8weD7MHkbZtlcQv6zwD5Mu3xe2RVMkeLfe0
KmUtAyu0SoHzwxdlQTAHEhpnTHS+gYspycgAcESwtBpPQIJHnrb5Ga4XrOzSsQGBv3iQtP4Kb2az
6WEYANnZEaKUPXA7x1p0ynugfJAHBPXcCamxgdOOR4Uy8HIleirNU5AocSCzwJ9L2cgisScwgNF+
3pEx/5tqEOuFH0wkwf6M+s5A5+mQvfDdBr9oRQqGMq8XbnyOPUtl0vFmox03TE3SE40EyOXupJOH
42AGpwOkWlCaeGWBktYdViPX6UpZlnmHIf819fbFU3uWWKVT0fK4aGMI4AoMEMBCGT8kdJ1XX2Il
hOU6+yJUml3vNH6RQKDMd/Y0TGIUiknNXFasTfGDGFgrXE1yU6+yswOh55O9u1xEO+N2Vjs0qf0E
tsc3146RJf0yGQnqjl6aVm1QGFJp/ZogvKXzQkfFeLGnBlZorfwambU2/cVmMpv5cDSaYYQnL9WN
Yc1AO6orLcJSMNLFbkWBy3ExpxlGC54t5Fg60Ppd1FMiC1johTMZdqVSevCZBGhdog6mj/HYCypW
UxmQX7Nywsu9Eu9zQaN7kYenh7kqUlU+CL5hOwoJE4jY7GcDtxfx4Eb1+HVrT/LxR23LHMDnjoMI
HktGpHfz6iA7ciPIEFtdqQB9bOhGb9detn/tNUkdCu82/3tFf8Kjpla5K2AEyAhYB5NcA2UrXaOV
9UMBplcdcavxggJ9AaYW7TMQNOCby/dLLXCxjufhbe/mo21XidiIQY+iKjMW/XW8RYYSUMvN2UrM
599Zrxar4+m52+I451LWkvO8zXxC+gdMSHiSJAxuKjI+fS3951YJISnFtEsw4Qaf91K8LTMaXZIj
k/oyZXMnFi+1YlE/OToSC2YuLljZBquCC1PRfFLE1a5TS1/7zXKI/sjgsVgGCILzxVlRGeJN8N1B
sMJyzYCgFVU/RZUd2X8a3q6+Ws28xsijwxHwtcNKL0LdaSovh4WOFORDCxKuQiakZB47+orKXx4Z
fBtjU0lliReLWJSbxy96qw1wMvKPs5aIqpC+eEWEGxmvuvWpaCQnoQL1JuoZoLhNH2VrL2IP3eWS
Qai54cKucA5eMt0FPdS2G5IErLMWT7o0PkAgjq/6rzf+6/PbH69xiEZPWTxU/I+M+AHaN4TsJ3vX
dlOuoJb+0t7q9Y8f1s/QmzC82VFxVftpp1uzviBKPkuWYphqs36P0Nsz7WYsMyxKeOh8701hmWtY
8GtsKWNpEdNWxZMCwtSqy+JS/ZaLYrcElpvsjVdPyGmow6iu60Nc3FFBIHkJrJVEYygEQyHiiNnx
c17SAVaNpudOH/Y5WrB3RFTtmR5UqMm5oZyAYR0LOf9qbdtV9jsGWTdSRFI7NGAKq7Eu5J9ATiCA
Ej9umwO+p4Hg1YNfOGg/Q6endNsJA6m/p7e8D9n38tNjFMWTm8y5HSbu7B0Zs0cluvrsp6jzUPwZ
s6LjCkrvVKEeT4teEHczVngY3ukBvSr7zh+z4DJ7QOgkdDUYUmSotOe5bY8CHhgRUlYPr/v0dFwI
y5amuEimbX384cM0DDEVaEz0PvSuFwA2DSsJIRxmCgKCqLyw5sE8+LCjq9FEwkaL9eA4SYl16RwK
SrhWy4h2W/GUh6In9WWdWigA/Ocz5aqUrc1ooVqdIyWSMkcyDcp/QPhZ2nRADW1h7UrRNfyECHWV
wKVQvDi1qRaQqLXzvkpkGLcg+o0RhvsHYIKLNzKmnthCSVB9vCG/gbppqL0eRpNJskRGUjLKnzo2
LR5xp99L8n6ZS+p+7MUGlqmHtiylBJQCeEfk7wQCGcoZXxxzSYGAiG7mimAY9WDMhPH12i2ilntn
sQdmWwBpYdF4EBSeegK+2wiq1StSIkmJLnjN342J41FV1zF5biSk5d+9S6qIQ6pZHulwT29mHBEG
xyujQDlxlZmw9u3QNNP88loAo8xLXyAsynGKUagzDfoln8KDN81aGBsJMl3o5jga8slis0QnMOvW
YvJz0B3iYNGyfF/l3Zm67VNB3Lz2Xif7kKoaCd6pEC+pP2ZvqtLvbAvepfxQ9nHYpaen/jRr4LPm
MWz8cGkUxtZkKt9Ka9xca6I9hQPpPvbVOGn2lkhsose++q6iUPM3lqbx6xN2PGU4i8HcWm3ysLP0
2JemrDbQqqn9pniwvDQyVJd3qCfS1ywe9FIL7Iml2hW/ppGS21HXadtZCUudB8YtmFx/G1lArl4O
MxIHp8LyNKNrvsr5cgPV56DvZaagmRMvzz9ufKZwTDz/LFP2fIp2jIJkR20+iv2/PIeYH2YMVX/X
rex8wQQuAAZtXmBf/jJbCS/C05nxDJsNsk9wTmWdp8YrLtv5fRaAdI8kPpiQdhLR+/JXqv0q6JEC
2lk7AEhENghMKS7CG1SZnHKLdOS+EAPobKmWLVpZ72VIZckVrgRHxJbCSP/m10sSf796vQ1iiKrK
txXs45lNbvputznyOsThCwhp0h4MEuBv65k6R7mNU9DZuFJq8Yv1L25HkYv/ZGiLOGJyydpSUFrm
Fj9c0EYxgyQ81ct2rTIs8YRhULm0It3k/9jqH3gh/nMTphkeLPaBnGJs9Snn92ONTWD23dVlJ988
/lJzgsrudvnRNabZnRG5h3qQ7n+nAnh6qmvVrUTcCkmTazogC0QVuJpYn0TEUXdlbCP+lb4Cry6A
CuiWEQkZnFIlEox071K7Nt6fRsLB9I/BsaXVTK5uKAGdK9hXhgqkEPlRO01z6btMtbLVk17Y3H51
mNuQExRfk0ZZzpjBh7jybmkeshpwOL+2q8XdHPvx/NNqSh0QqM5WO32JpQ5G2+RaN+kOpbNoaCtg
Kj809RtjGhWNPIYH7FfG0Lg/2d5QkG9b+EkVAF2UFqSKELlYEXxe9rU6XJplzV8JBaQAnRr0pK2J
9QWbv0nPQPp8NGHyMX6SCxfB5nOy+fDLusiDHB3D1FEbItrC9KvHRfJBgWPOqdk3+r8eSAOdHQgu
1gAmr92VuNHSxwoG8Lw/tQ4WPCTJ2/gJI6Cgw6+TSNK9gvmfSng67tVR5uPoOSj7Gl1qjSUM8BBb
uvQw7XOgHM8jHmcjSn8pye7JEufq24AlK9xAT4OelfXVZIqaFFgH2/nMsb6sesgL9mhWVUHcAinL
4LDd5T4lk0BCtIVkUcdkJu3hqj9O/K+kF7yRZPV6q/jUiMQT4A5HAOVsODIqqUVc5FwYlMvq+6Pc
fhpMUN93Qh5vRDPeRgE2Uhd61dkhROj0lFcJ77QiqqHlwiVOWHAGIXB54jdyyFKW6OPLQg35PQiL
sAdMvKiOAjLnTyTVZZ4yiPqlF05cAvxH+50bX97vuidJX0NUrWgy1YAq+WCMQd1KcWm50V1gHGRF
8FCUppC/oko+fKBZb/RvwxZ4rtymQD5CuHJEnA9yvssC2VRtBIIUxnn/ozg0hgyhc66/2q0PvMvU
kiYVimtjIQjNjsNGbvUqToTE6YCWbPDPVHhiG0tNCGSFP149gBrzBcSv91o13tC5hYxjQa1z25be
+vpIe04E7W7YZanC9YWJdnX+xleTV2wJJ/oAURRu+JoDEMgCmKF1wF8RB5jmSDpKMpjrQL25lNFq
YSWwmPT6z/X95tY1qt+Hd8a7sNdxftnEIpwrXU1Y7Jfz2jC8QMA+Cg83iJ43wIbPyTUTrwsg9r4/
PvAAX2Qg5z7UPJg9HZ3tQPXX1/qTp1ykA90ir0yXzaXFuVN+fGtnX04MLtkOC/gv9zX/xsTm/A1y
Axygnx+mayQLmTe69QceeFNe1cRVQZh9Uzw0jeZ4sgef2GdTLm+ITvikPv5a+K443ikWt55HM+M7
+gN7cQOcmugVXkWFRbHJcLgNhy+x6vP8VMv2yge2o4Dgn8f6fWngz/IKqGiCpF5ltD/EzMiV8YGi
BAw6tAMm74T6EBOd3VKFUA8qkAqhdxFHXQ3r0KSCfG5yyzNZA1ZC+8qbDfHgUrt/NcySekbSofMO
R6A5ERurtrYElzRrccHzuzWTuK745bPpIXE3ZmNB53RCSzvQwT8zub7C4iIH/oWlj9wDQ/+HPXjl
zIRNdpUB5Hmk3I5H4hbqFOjtbgZT+sIXzS13P15fTSF5FbIrMUVd/2IxEQYpViokgGo7OcsKQX9y
Zq3e/8xSFL+zGUqJZshX3ySunYY1q7GGkhTNQsi0zxUsce6j9eNAGu5yVW7e83f1xE2gDGfGOQqp
RlJyXS8u0wahRqzS0NoZhGXbxg9qx5d36UzGuIARFYSn/N0+in0CLx54BN2i7+TUbW7EjMT77YmM
5VB1YGu9nre99R3TvlpFH094UCF5JyrCoA1UNrRdBrbs65TeNML2C1bqJXYzKDaLo8vo2MfExW6e
0QrAcIc+0V1WIsfPqjQslWHw7vxXIL/y4hiLmBCi9It+7JrPxD12NdnMokyfH7NWKnxKirwBTcSy
C66qJIhs6J0CeT3chdK3GGEzbAb9I/tUr8cC2K0ghKt6L9Hzmpi9RtS9QBohr7G4dX1XB41JoDFd
EpEqqhVBJH5esXy6O9UySZM8jrXWHS9sWzmtWd6WOcV6cmSrOlReB/HTpMtcKCYgIKLmvzd40x7d
u+7v7KXZ3n9ptxKdWRbgkZrDqzrZU2SoB8/YVFPMIrgEc9OF6s4eK7mPHMLu9M6K/SGzOHXSWz+b
YAi9UeEW90sEfsqRAAEncPAt+G2cmajt9s0CJfcZnI1hex0l2y6h0qBmpY065gst//QeG4DWId/A
hFoMXbDDtBcS1FJI/BCo7iDN2lq2fmcgI00ZPWV1zzgk6jlFmw3CjqhKSg0Ry5RNZcoY24/X38fi
vLLgBOjMYW1Yx/loBNvuZ/VGzCntiY/evkP2FA2faMFRLtC64jExkjFtw0TK+Za9LWvpktqG1h7h
kpOP1rrCsB/JZKy6Klncaia3+Dm1bv5A3XJYtohWcOKJRQFjvWJUNJ071N4HjcwG6o17Le76cpl8
aNBmkTQOpKNOcj7q3upsWIoOyrsRZ91KBYsQ0oW9uzAupMYI5TIj0GPkPtzCTQ60iw6oWtaUL5b2
GppUvZIqTxeZJpG853WmIRZvBtIkqV88dH6w/Vua3e0S95TL+ZUGwYpbh2V0MV0SSeYV8a5OHAu3
jKnQl8uWnjfVNkcz7ip9ohwhis606PtGGxZinCCT+v9fftGylemZ/Reh7qlNu5svdBJzGdeyLG01
6ZuoQ5Y9OV3M/V9VcELq+wwrRcJiuWT2xB30SLIKSQ1niqKXOeVeu9bK3tC97R3wvt0dhUbnuYKU
wBXmpH102vp6dSJYyzJqMEPEtiptxjGc/4qFTubJnVCOLZmmAMQmdJ7pdnCgs2JqMBq+y3S6s2Vl
Db1rP+xv1K1pSWZ4qDhURWp6KdQWLlPTC7k/4gJ4IdKjHcwUemDBlBT8Y5KRSrhPoo+B5RUbFp5u
+Pf+tspf5gmKJe1HDNZD6fIPpLvQcz+5OIh3PXPD/sLWFaiv7LkrO556e7uCVzRy1SINNnAWsb4M
JfVDPp+lPxRCV48eyV3I0qJwlcQ2VilRHTPjRu9dYCjdQhMKrgfwbr4Sh/8RpffuPxUZm+veLrxH
TKr4sBxeFFlMlCbAphiJaCHi5ANFMsRSuRLMLRSl8Meq9OCztdeowwS3czfDC5Uk5Cx5zraWgEgR
2UussiWnxOtiBdV04+5gMWX/I2HQDZI+hX77q1frski/4LFnrmM3KPqXp0BZShJ4+TarLjsg6UR8
bRa3PnVRv+ImXwCG7V9VwkwZ6GF0qwemFAW8vv6cYVzjYjIatf3EhobSkjdIrSVf813UaWDNUBZ6
wuJXqhw7W98m+1KYBk+s8BLeNJu33NqMMTY7GaMl/pFN9HN+BOkSBAQBAVlWzGQ2WJS9JOvDHkIq
/yFqweo3AbUIG81igB5bsfxq+Uv1CImCw08LEWATt9SF1q0rs9ULb+Y/UrzhPdlgHtpwDRGUEep/
hqf+ivSP363TYIF0J6/fg0mlMdOa/R6a2hHY/t1l/vWzQm1pzpUthU7coo5xMin/s1RukMEANVqV
0Ft04kOhPeJm7UFX5ZIa+xXKkAKGqrqPPCT5LHKhSuXL2/sCuHlojtwJBSdT2BCRu2h5ER/OMicz
hhGjXmAptrjrzAxZtByNF7uO50ahkkFOlOUZAbZC7ZVjsnS7v0mCWwFGjt5J6CjLLAohGFfgELPj
XKFkFfqG9ORsj6QTHLDMElhVsUO26cjCyid+QJacFjTrr/VdA3IwpJMkuPoHcXvfx9UXVMr8/fex
B5iAEFgcAZkYb72RqbzUceZcFFYgD0mLUgRsPFo1Mkw2sMQrbp34cDwRttqRPYbhcxEztl1wvbCK
xv5PMPaZGE/kW9raY17/jPQ1Hwy+wsEk4wK+fFGbuyZmtf/W8MtEeHS6dvdSAFvpSOI9kkoV4EOa
He28aS8g6rSZ6bb6jzXoyukWbN+m/CC+Ge6837EGbQuhvaFUo0bBfozMR4g77/Tgs0d3j7pt9rkS
KjT2Bo9Xe6QAPeNtykOZ37vbs2X4HPwjzL+pJk+Uy3vK3uDBiCN6+00nTSV5ff1K/hH883TQLtdB
yjQFzwG9aYaPcXD7xkQ5erTzW3IGUhrYD1TuGd4m8WYGoYs00Nmb28SLJkLQUP7RXs/LCrCLfhAn
cOYcZU5QqkAQRQVc9ltacgdbCUrm2vY8RaLIn4wlDHeN9A2iefmvBRSC3vCJ/Y6jvLuxp+FdLP/h
XCR+cbjXhuFWJlH08QdJpVZnmlA3KSIWGaS7zFpiHsJ2ZA4Dhor5D3xGFzuDhHxzs3gDJwfoqSV4
v23MaDlqayASP9qwEFonA/BngFBAfzpZqC5ltZQ6iWZ42iXJlOpWjSJTwhID3mB+rDvvdGpHH8Lj
90M+cPJT5QZ/+PgiVYzCk0MO2luU8Rhgql4/zGGph1d2/cnKA57JZ0FV1wbSmDJyIvpLKWeN3gcx
QlgDe+7EguPNNRghsOefWcCUTa3fKs1vuRtiBIdzLkp7qGCaejUjhK5rk6z6q80wYOsoL0a6V1+v
iPD9OKx4weLI4pF8STXLlajuRuYm/gaSH4AQdOGHJToj2IOcxcN4wYSzq27Mjl+uldqe8ZkXYWko
B8aso/OZMScLLJZRv6tC3U12kCZRsqBpqBuQWgbqVum5wcgCFOqfRiy8yQC7mK4Q9IfyGeHG3g13
EL8AYwpG1wJtEiooS1ab5mgb6DKFnCvyHiOt23fuJRT1T6SYfw+NZYJ++45jE2Sr3ulhYvu0YAkv
cTryAFk0JxDlhQvwQNfRiDv7+59co3G1NWd6J+aLytjR3I23GfY8wCGPflxbDHRqroWHSJEV6mh3
iqTbjMNXJ2BeAL+MCSQnMcNVSYLPuGgovrAuV1mPePfCYb/LALwzLHmLKkFb/DDT8C3h+nsXgljq
RJf4zuQHJUS0C8y2xsWQn2IYs2mFOBS0eYs3CA/QgOkUMxkUHtrbME7uPwtgmeYE93z2OnrKWqbl
cXkqHjfCTfeLR9mbnmtECpYPMNtfSLaNA7JpOoPgzzmcfEC50s25nbqhwMXLpskXPbxe43uYisds
jf60Brde+y9eV6RA3SUKTg5OSic9wCzZ4mgKAATQjZqoPhHHHIsP7rKMxUB14AaZnBgezLsbp+TS
D1BrXsMUdz4aeW4Qx07OaKvg8jCZ3W09pWcHVJNj+kyb5QCjVy6b03Tk13rR5Io5zJa7/iRan2Ya
qcdfvToMAOliAtm9XODJY23MF6/to4u7UB0l9kL9O8vuMlUA8t+gOMkuPjZ+5gd6AkL3SDkxr10l
GTUEuyB5V0Tz8vsonVeXL9O+sN7zclQHIrWR1zpLYmXOmoG8OkWcQxxDxRyQd/wmZoz6/GQDRHE/
5sspFSFmCJDn9/ip4BKVPVCXHklco3oW00sVtLPZHd/0KmBxY6MjyU1B9v1OKUHZMIooumX0C9BE
HaGP+vj2B28fmUII/r0REPK0MyhUlzRpx6ITdayv0+gymTxa1ihsGycVP7+3g5z2ZWr6DfgCZQ3E
7l0iy4le/QdIQr4//PMJPPW8IPNwpwjxroMpDlSVw4pFuEuKgVSwztGtGuVfB1IsRnMgQI3fUspF
jSSxzMuMVYOcIc+63up+3u9WB6se6GW3nSmUlSXEIZxy93jIBTZ6xStZiK/t7i1Tnkcg6B3YHY3s
s85h1hDOa3y4fu/kddSiTxCfJYHO8tNwyutFpzIi6uZ36+T1i8Ivtrz2DiMq4D2YlPO9RstHpZw5
2xGcn/N5pEY2JRhdn/sp6Q/Oaty3iuOWeW5sd4c4KKBkoq9s0dfa8ihLGIQkpSX5vINk91OaNAMT
J0Be3em8ByeDt2G0ki9lduuJR9CK/ohGSee6470Stqzvm8we6BU0WvkGlmvkI7Eh+3ShAhr8B4RO
ydi9Ut+GEq8k+d9LpQQ5kPGIhzZsJXVcOnGV7Ao9igMpq7wBNDA75vSWMyGnDdx9hG1H4D2SFcnn
aFxzNVsXkq7c3qZBki6tPybxXJ80THDsodmIHYbg7uy/jT9Ig3kdv41UqvnGAk7ggiibv8lQprco
6h1jVsHaDkGKJEW5RerBm+pAVoStHNO7d0XnGxhdG+QziUtAzugECrwW8T7vGhJdoZYxbOgND6Yj
jTewMCPmkprn0KzBtZKR55BrBwgIFKR2t1rRr+pTmzB0/C7KrwAp3J+YwhRJWIreIJMxVv0JqqTu
6fFxDQqY+d9/1j6f+DQ9x5xsMfAxnNHgxIY/pXu5HCQ19QQG0O1TjXsGCPvRqA5IIjBBMd6D71WL
JtpRBXYbm2vYIDvxVQ4SiU5YKqrAsdfmnL2ZlWl0MwMA3kd8u6Q/2Eb0BE/zI/3N4qEoUwpJ73bV
5lshG+Q1Bb5+fDCRZPdc6+dmA6affayw7Fy9KLXpTSqNquUhWXAPis2uclpaYPU3+rYrBm0kz9vk
A0mz/1pBIqTHHVcctfr9SnlWFJuaOb+VM6G5LhiQSDWfLZrWrEkqWgts5XL/hCerp395RH2V9vao
bPuUez/F4AUQyFHvtcAzJrSb5J1tQzxfAf4yMCZS0ejt09wp25hDbbN0x4BhH4Uduab1Qe3rnNqD
3+Ue8Xg05wM6Nb21jhr0+2EzhLt9nJ0VIriSAYBxwrdga+w8Dj1pG5H1cJ9s/GJaAzSQsps/aBvC
kCQi6oP4CeQvhMpAho87V94lqDZ4Tvcr5PHwlyZXPbutsIkCXObALhSy0Q0IWKM76y3q+qAEi19j
hzHT1guUuoVv6kNIouy8LysLdczKitoZpOJqEehapAdK3hihdSteMwyz5c53oqV42k4W3eAanPCT
+XyQZ6XBCjKBWMGxipsdholkyJyIYA1BiBZonSCL3oWJEgP54783ZYuINWKobaFdDIfXXQ20JNak
i9gbbEi/mnwxpPto5jR4KqVjgAmrFuW9xF3A0RHZrbXpKbRJzB/4n/UPB4QVBNYKxpsDwMPrVukr
Dh+h0xOxblYu3xm7oooCcJeQjsPXcXpGiHiBOWLNl+1dmcYDo2BPZs4iltWNaSzhRawfGjUuEzwA
QH9lolY33GOvXd/VuCDYVda95Na3p7OeCwc4RYfHhilWDBfr7dn5P/q4uWhy3V2zbemnauLiGh9B
uYzx9UYzBGPW+HmYHweW8GuVz8swo1NcVqGFTWA6fcI1X0sSgos+nGRtPniOFHI1veAQ0PAAOLgw
+aQ7minDKE1AmhMtv0hOx5w5p2zDzU4QDrdOhstsT5zi4wUPl2I6kJ2hPtx/pP6IeMEHiTSX1XGq
KbSAm27yu13LK9DKLUQnpmqa1WPSgnhf7VRoA6kb5ywDrZw4wihRoXcSWlwKKRxquyyXzfCRlwNb
qHWkUlDB+u1A19pAvNtOt4HTTcbuIdJsQIwQtuJR2hWAqHDOcSQ4Uocd30yeyESjRRAu3hkYyniP
kU5xssSRB8kPLDeIpVaO3rYOpF2+QCX6BLbNRJ4+k2R2NYl3lEt4UvgG9k6GlotDtwNFQJ8201GG
mdV23vV8SmXoRk2qG+HL6/oE8a2CRkd5W3SZ30gAA1xP+cnMvbzZQVchme5S/ku3MfUrsNYoISkq
0A0h2LdP/gb3w1X/Im3Y+3zwnoL14vwtXv6E3IvXvBxMmdRex0P8Rmv3ibIcuBk4cxyHCfwtlEfX
9dT8rHisM66ACWvs+QVZeGNp/JHlIA0m4g8XJEbjrRHsT/l+tEAACmsfwn4+Eqp8WwGXnh6GCWt7
U7061uIsKbYENM3iMivF/6hn+XXD2y7icrlOisffOoC+UwNE3TEKUNyB/pbkYjZWW2y89J5i9WfE
5ZP4FxjuJ1i0Bz0mI4czpjXs28iMeovaZeJWFRfzLt3ug6z1zkTHFBQeBy4apVzc1fS6hSY66Gv6
hoERmA8aGUg4O8QsC8Fyphx69ZJ2huydeGG3m6s2vK1s5kzX2k5GVgngVjXEM9wnDlQumflApPYK
mzHhoF/fdhCovJ0LCu2xEp119N3LwFVVFer5awHzqhD6DftjIxLy11I/owx+Q1+RoTN8VPVcqHhd
mdvgf6AKhz84rVRVGx2mz7AF1weRsJkSFFhEap5HZP/rpimS/pgsvGY9Loc7Irh9cgoKBLPZxCRA
VCAeJKsUoeJ9epqRH8BWBkuWXu8ZdZzwWFmaL0C2vTCwUamJi+dRJ129OmL3JoZ08raauD6mSLD5
slPd61jFqcSqcu6E3wzzzci7SYol1mw0w3QN7q2JhyNkLD+/caJOSqZcMWdGgM0BvhaHxSPeP74v
hHoyMWw0sL/8mAYhurUxMKoGNkyH85s1bCaXNIUP1vu7QyR+6pQ9v9dSKQSy5REBfiDiewGuNTxE
MjfEcFU2lZu0YdrGIrU0lsWt+BUS70NNdE5CfhY5qA6xet3xuOLRJnkRehofi7ofRpaJwyzb9hTB
dVsyzJ/0aNAm0blsyLsszjW9ahTAslKXnJ+QktINN9F1QJCurUzH0BlduW2h9dMbEg2FXNTZTaev
gD+ICUWFndkc7W/J3v7oVn0GzR2eGC0voOnMSXPTrU0gQ23Ap9uCtgagSp9cSy5NN6OOcAWZRq00
gZu3bebfwvr+KzCBcSgFx1lXr1wGy/MEguLC11fJwqyH3thCuzQkzsrl3CXotqr8/ElJnF7sxLT2
x9SjX68Z/YFbg79uzGK0keyGVuxOBsGaHSavpQfsNKYw882ol7ffwqHsMoc7X2CBF+Cv2ET34A9E
4mbB12QLp+u3TqA3gEySnJc9CaO4XBHeG4MBMepdOQvDb9FkFvULvrZg6WWWUjJjr4ZGx9QTL1VC
nnJ4JGj2/+l4uBueQ6ExcyXCGt5Mrkkb2mOlRNvN9U3kcLX8Mb7guGAEEGBQDGFobT1mb7r+ODGQ
TLOI1fhlzZkJY7EzuwPHNBlwYGXSu1hqNIKJvILGCF6AS8wjRxuOK0h31IXXhHrLsmv0Jd8ZpeE5
IiMSDfFIVSjeJptOGL4+U7DePdg7vt9T4ulXmS07AMBiLhSucYtOT4DiUlyo15jiZDPPw60OEBx+
ItbCzRI1qKNBB+uA7bd0m1NL5s3UPqvt0NHMyf7uA33jXL3eh+fwemJaXVS+h/enyOjibIS3b68X
uwaMszRQcfYyBVJN8hY41Jb+33ELwiVbt2CBk7mD8/wvoPPd4nHMbFZlGdejd5XlQ0Z5/kMTiF9m
TM2tNN82mM2WRJY4WmnTYAQtjJwqcVq7vSYQFS86XZ6lnYpFmVw0as9tPRyE0b64yBiJFWZwgMOS
ejTo3+Zfa5VO0kBToDL4607syovkHMWmEK8irrSLcSWVOVQnaQyyfqxDuiCKFVcgdbYVtMMbsz7X
ToNcApHnuTg/CnpWXo4StGNc+Wyzt4236BljjlJM7ha+XB+m/q/V9GbcQgRv9BSPO3/s1Yq2OTXq
VqW0kimp4ZFOn5f9K1aoJ8GrtuC+N9r7N30cGxNrOyVJs/uKd45O8q+YxrT3AAbpDtus93iCFmCo
/bGVPh+wTOlvCkfhWlJSYQYCEbyz7vompIOZS4HmOG0Z9eLN6AZuYId4K6MYUoN54SLdi40I2XVO
N/wO7KbvsvIF2c7oPWBKcp/GKMW86KSnVnMdpiZk+9nW2KgyJqHwHNDidQ5zVgoTX20nITJvaWpC
BkPtoydX0YbOFJkTnbKt4csgAJbZbPMbQv2KcXoBarsw2G+iY6X5betZEiry0jX2mUDjpsW2WeJ4
SdmT7+yndpnAFgKwAHb65is55/y6qv1fSGnj512rZ9SejvHxsRnI4IwDOkKTzUm5azW6pYJIGMro
Oof8MuXt8hLBh2NBpm43TOxqv+xhKIpAQNUTpkBLa7WfNEtZ+SgZDCYN1MfSzUDoJGL5bDH7UZhe
PUNy/Q4sUCyikLftarQCnYd99vlOUX3J//TaeaTpV3v5KR1CpuLCbjXjlE02rkFw8dfKr47FD+Ye
/w+wf38yEUTuXffi3zlwZ3sZZmApm1SKRV+nj8orufmmLo+9+NP0k/yUWwXTtDX8VCODuyi1KVWy
/25O7KvBBTihEQzmMWdBU9I5SRBWyPT3v6xHGWFkaRLijdLszi6MrH6kbm2U4E73ueKiiD+f8CeO
tQBepS6z13qCwNsc8okFKxCO7EjdBGQN2/k4cFHaH3CFvvJycrt5lryK4yrhY1+cLr3vkj7y4iJ9
5ZP/5BjfkFl1/MVl20r6bZwqzj0lQU3upcAgrV+h4m9G8ur0BULZDTzUitK7EbxnXFstRFlqVlEM
OTpfVyAKdLDlomqXgydVgYjo6XuiqelFItkbofHZJAgHdZUUdSGGBGoPM9O60SLG4B6pazTiMo9Z
JotMnU8bnO+ed8NX1W/JJJXH7XDYrsolfdaJP6sOTCizcuxnje+ZuWH7/4Vg4jn34SRZCDUFnkAx
w2gi1OEsHgjLbBIWPhRSzNjJzV/B4ttViRZCFtJ5NXn81Ze57YkaSHvXYG2R1bGWUmvOFofyz0yT
ec6FJPIwlBJU08RQzl4rOrkLRR+3BG+nYLfrS6kkWu1LNmkCufKOKWmetpEssyxp2LVuz5CCJXL7
B55ho6lbjoSbwZqNWVJ/n1VelqYlN3aWNBMi855z4KQNuyhx2aYIGi7AG4AoU3pvmvfOHsx8Ac1s
mZw/wvmCK4gTCFlXLDxM3EL5TJwcMBJeghDWf5LR0Vjzavn36bxlLLGBLVq6GmaOAHPKk07EWrx7
x2IV99CrC4j8zUkWdpJWa3RMXrU6VcSrsUpVaTNWD7t/K1GZQ01GQAh+0F3zxkpCzLV7rzC2YMT0
Cqy5G2tGAJS7l8exTuWPcDIoEKkl1sA+5xc3tOWLfqJzhEDwMo2n8yW9H4BRjU4nbh+tF0koZ4Jf
U4t5Zy5Z9YynY1/pgdJNJHd72zY2uHt8PJSc1wq9A1kp0CCU/nUydmNUs/n0R6RR+Hl42kqs7y4v
FHekjx5BXDlsoYPpzI15AVktwzziwF/B7GmdAEv8+mv9Xxf541Dr4YwJXdxg3JO1Tx/vW6sSwpcw
UnrDBdskRl1KreQmH2/N9P78ARLFVpVxhDaoWu7pnzDueyfOGx6qBaNoW0xXY8EGfsT3lslNoiqZ
NX4ubwiMM0+ettVsabvjAFkU+mC/ElgZR9sRbYCesuxxdZHjMXuQga+drXkOtpHfEKOXZWq105y4
zbg2CKKSafAxsOVc5RefbLkNQL9/XQCratoaRYDaILXOBfv1YsnR1BM19eInHRSFLrCymNXeQBZv
0Kil0V7NUi4YTrYyZG0UYAYqcrDS5xb8ys69ZBcvTxZ8aQP5qeol63yZA9lPMO+zmwZi3hUoQMmn
QrKgjxI/lbf4ATFdHxKuHRJ+HTMlRZTU1ZeGHTeEkDAq2+4zcSA3fCfK0XYhvyB01MiHZJnwW1Nw
IFXbWgHh1qGjaGS9BzGprPI5VXb2SjJ3AOoBdQfdH1ceGxX1t0ynH0Ix+lF6eP8p8is5j/82llEF
VdpCd9vx+yTkPvFPQsgf9BVSZ/TxEc7Viktnk6ZiDuT8KOO474RhEKKvFlKp0HyQB8aphMOKWoZm
mmGFO1lxTffjXGwLK2lKIwCoMi8BJ2vLPyLanV7pm+qdlA7ecLGmlKh/268CdALTYFoKuWd+5IjV
h+XBl1zV9lLw/wRUffo9ZlAiENjFnHu5YPWGAyyXB+0vNMLic4aZMIE8Xu3BoKAw9D7VuWLb51V0
lDlz+OZ2WN7faQG+iHynFIsQvY+3UX9PvgGJux+ncrh2Rgxirpil0xsH/gz2Q4kIp8gQRheqfYjV
LrN9VeqpqExba+HoK5ALIlEeYqq6k5/ATBDSrL3MxC1nW+yDyCJ7yqC6iLysmw3vAssxQUHPcL/i
7F5q7+O2/3M8TpYDXLmPfaKp4lMvhV7BFVyG9dYa9lmK9I04YAifOMLj5oEaFtJT4cpPG82BXR64
gEvqrFJ30jtM/exZVKUDkoxEcIlq8p87jeVbhmJKzd1V8GoryGBUwEIMgcw8ro8fg/mFThgOOepi
vTjbRPATIq5iWPhYNVhYp1ir5HAM+Q9n0lexmq3mbVstAZFAqa60qzYXHqhqqoC1Y9ZQicLax66x
aWG5kHY/5mmsPktpPFbkOzEUq2+gB/qyDxnN2+XbxKYpr+dKdols5/MEv2u+uUJ+PnYKXlDKgciN
jE2pvzmJ3weyKJ/Z+tl2Tr5zoI9Uvq6K0ub/KcwO6fVNp5sDl6lqicLSwVSoJoTbAuUVojBX7Y25
+6w4uU8BVl6uj7Y7ik9M5xeohu42fUmLwiLLUtikHVprlvj41Po7gOwiu5D39NCuNSIvQNoGqvkU
l5W6A0GaAIdy0lKnmAyU1pgTmgjhKWBCxg+2lfo+YgnW++k/0azmBvRIiPnwfzj2BN2G0xiEj7QH
avzHtqZV4yBkmFN+k9ITt85Q0cNVaet8jpiOEHMo/B3ABL0Lz35nFx0lyIuWIZOkzPhskhraFBze
M5rhM6V61CxysTOY0e3AA+mLhqXJMairEAVPdP/Ayx2Be3YwxcTJVF7yoK+FIScFixTeD66NEDmG
+YuJ6eVvQWUxYKvQDwcD9b7h1SkZHYhO1VP61+3rPB/lUIc/VumSHs3JTPx3BvKwlLvKq/rcId3G
E+Y3svLml6hV2ZbtiD6bWa3nfV9GU/1Grk+tAPEYj8dXVFTDXirvCgNSe7eg7WUB5/eRZMe0TkiC
fAB9zbS8IoRChR2X3V1RxrnNWzOci2rD0LwptVUO2GwUoHVlj93RQEJq9cWG7iZMPrsMnlIHuy8P
Opy33hFzkEcLs00dv2h3o0TQlCUzHdbPgQhuMjo9Ed87E84XsFReJnuHD9pljWWe3/TwHPBz2Jcq
CxyYtUnnpNJtnplilB4GL24Hscdt3Y13eKy7QQYOzKTQBjKIRccXB3dKZKVAL3tlqHjcEl4ETIua
w5/VS8GkBHUXAdhJMdVLb1ZLrObzaeYANTaPbsBccSiTgx+mQ8w99jwoW/4Ozb3H28qMP4jNJzIB
qJwBegwKVgd0O8h3qS/uCYGta8QhQn6wb7onnDi64fK3ef668GixM+tQU4PX9geCp+Za2XurONPI
QnKBIMud0Cfz/75SiJk6CIvNzD30Up+pT5d6sKlo7/B2ub4H2WdBlKkV/Ra37t4hj8nXDUGrgzez
o+qeDpiqGkWRCGjswhOl8qPKnnXaE6Qxu5k9l+tvFAvOjYYzIkrDQCVUKe3gold0TcXnPqCh3uFM
+dPDl456rTLp5CpUgnc7nVFcD2rJviQ46RxPE2Sn09qByXgxtc6dxBpGluHOz9Cqe79VXw9kWFqN
IxVAepheE39rBBikUQG1y1ITuIqS8MvcnWtoKbn4NvTWMVDEssM1IyIxVT5UEOpK/dfinY2VDS8s
a8aycR9RXxPCCBXOT6bqnKTW1Sc1eL+hgD/5z28iqstWEgDTNkzgfLt0HRvkQvofY9/r1E8ovacQ
GiPlrlDN5N/9m2bLn3Cbe0Khu/y12Hp29s9FFYfzSZ0p4mpyil8OReHOA81ELHftI/TQkiBBy76x
w07lUbuTRYLwE+H6h7sHyrbHdsmOhxEJRGbqo96MiHZu3xIDr9e+grbmBR9UQM9iFTXwNH01thbd
TP74ul6fOiCiCLYoLM7Ku0DqjmQQga5PJnAwRDgdcm8HKO+1HjROYTFG/QHiV7Np0FwozpDuvAhm
+FscsbMTgRDSVHRg6IXVGM7NynajO2L2Mx3DBr6bNGb+DJkaYsGm8XzZfQNkgZA6ArKOlhkqOcWm
V7pdM72Yv4zIisaZ2Nzo9ZtmL1nfqJHJqdBHOc8/HkKQiMtcQkhysfV1He1Yc2qlh3m11E8KEuhS
RxUjhQH6yo8pI6FCTlGoiMdOIwWjXBlQVS7TyE6xhVQCP4T9PDYF5dE9oEgcGwuEOTT4mgo8uiuU
U0ejEwAnZAv79Z7nEXFwayGZ/92WXlaofR8ksn4ao3oQoEiOdqdB77UgH8uxEdu5mbl8F6RKpJDc
hAnq2UfmkzSp1zc/8g0pxwvg3/OY/eAKbX69CZJ2W/oL3af+/8Av4+37xhSSvl0RntMFp00UPg+c
XvJ8PrgrbW9D1c8WYj4PtcNvhekOxN399NTbMWtZaletsW22TMGz8OMOCcFUDP2PKZ80v0labGsH
uQ1JiDYN1wOXc12Df8CjcLu+HM1/SpNXnsPxzqRgbXPMipXmiDG3iXwb0niGTmq7JDiuFHYH5DxV
dNu3D3K+vygBJXAumoJCYZzp//1YUElcakxl5eMvKPliBbpdtZKtxmB9mM38kmEY3Vm510hLqutw
t3gC8SC/vGzHM37Vr16/h/D4ZIJXQC9YUhlO+3uHAYhl19IncA/INyeVoihzhKnhe+rr0i8eTFW4
G6Pqed5u0Us1V2PjRu/6SvTj17OT1ME5VUlhPOUeklfuWYPGxmJ/mjOKB9XuSrlGz/xdLMV26HZ1
VHM3E/C2H69D81RknN9nzct9b2N+eDtoPKo0LotOfHUTk1WcTCWB2hkyXsy8a3h6KXJ+jysjiPgt
13tDKkwb3uaaI5BcO0nEBTaEaSNPo7kitQjLB24joHn9PzI8BHBnIGwOwYXBEwBgt0OkZ0X70gFk
lowm6cs67OgYV0wDT4iNoWCjmfx6D6jQq/zBmdGRbAlYSDaW5va8r1Jg32Cp8zh6+9pI6enkbiBK
HHnboiat035qbFqC5lM8CkodHKrGhEIwN+1JRX8uWB2yV+SnQwtf9xs+JDu6IRGe5Hjlg5D9BzjL
uZz9hX0BR8YkdDqNbi8987BuSgNuQs19lpwzFz7s9FM1b4zB/bBIkbddZNeoI8aK89BVT7XrdPSb
EuNB7EmK0bK5jppS7WVfP3tPqpKQuh1DPtWjIMh80rDF0YCSyhknYhBdhZwnjEl8gSSbDY0TnLkH
Vs9Fn/1hPULIb+Fa5kGLkTGH0mFpMJUhAUKk/SBuwnfHQvRyrY293h3oTTCclFlkBb91IOs91iQv
293T92w2RPJh4FLIXRU34euTDRQ3K87N0xbvSXgP2lQkOb7jG+2pEQvXcIjLxwjrwBgPruQl4GMt
Nl8JMsPuYzcZs7hdXm0F1iDBPs+HCFjLWlsP3A/KxHHZ12i7HWt18fC49tGcLKWsTS/eNOz9doRe
hyzH3kxirUc3iggXQAK8F5MTML3hKb3tnvfc06VhkO3d1DSVyq/FZB9J+U3n2Ei8WhRWFvycc5hg
D4Nz6FAnUj91ZImuJgzFCTTXPW7zAX5zUMn4L4MMNh6h0T00w/Dd5qPWrPagQoPwlRBZPIZTzMLW
LkPmImAoqe2ecwrZOMX+9egdHlng3SBP+A/x0qEZ+zvXeIzVS1Qe85GT6m14UdoXY4pI2I5ssavV
yyU0Ei9ZAHyNz98j/jOiueJAwBMklBft2esranTpEQBp7dSSWv7ccuLMdB7lgNVR9kifB6q4sM5l
HfnzA5aa5WZBgcpzE0T9pZgZaQnG9UGf7+c15NXdsjDCltc/LylnTkoGrX3nqgX1TIszUxkxRjAM
RLTWjEnKgt49mHyCHWrhu/pypTDJZ/sdf1UFHB6BT0ZDZQExLpTWCFxADg33Zw7oVN7HrOImM0cw
1Lx4sDBdEMuO2H8TOft+w9KoSTwnKuWn3TzylaoxKxIH6ZFG4jzkFGGkljhAOYrp9aiodiX18xuJ
haKg9es7vnDIXGbXzJsS6qIE7CElMvXhVwWR/kHi0CpY46qCiiw+NlitfqZgt/sexu+BVIZoLBJl
6VZsiSfmapp/WO0GAtslm5wqtzVhcI65tT6/kl/gqBxpFsOEHcmI61s1LxtBH/Ab0QFBhfhRHBhX
PdUNc9DmNWH+qLFjGGAWETEgaYVzmT3t0ZPZgeRBJ1pGQc4KYTM7GXh6eRcDlrMUYQC1fhq1J5YC
xAPYr8mKD8pHkFiNLIoBNKL9eRHLLTXVEInQYWv+o5DBAwxbJfDlFvCzB6Nodw9I3CtGsm0Uv5pV
uUeHFPFO5Q/2zopCZcB18RErTvXWon0yylJfw2LqlcUIClcpbtPdb4kD2uLI1bqeh466i4wFTAji
Wz/LutBkSr/gYbt6NbI7kJRUgdJ8apsVWn9qcgUCR64qKfnFSuxBbiTW+MRDb9WDT11mYo2fpn8g
7Jeno9ff81zzo3vMW0rSjGBFmuZnqwMYgV35iI0g5/sytQhQ/G+uSAJO4WjXhYJSQLW/+68L94v0
er4+y1FF8pmrSQoZOfDMwYZ4LScHgfEBcyV4Ld0wvSeD/P/YU+1Nl76cFDRyvN7/gs1iISzmljcC
NOqOlabqBPMm/BiB6SmhHFotiQkRy2jOX5dVXbah8uqEQeNvsvY4Qi/k+jTegz47ucoD0wQSaKeN
4+TYngIc211HcDohg4qijn+ofMR7CSoEMblNboCpIDWlUZxw3VAQvCIO+OABzy0quzHOTsYyTw9k
ySbz3pZW3utsfKlI3xWb+mYFlqQ9izgusBqrHG9GL2d945HEX2YClrqfKLCcbO24wMAgFwXCkohi
OhXDUcccx8mqdxIzzV0XBNKBre6xBAzmvCEvl0ZlyTvVDTo6q4ytVG29/p2mof92MmwfgH7/ARZ2
LNSRaTHM1VR3Xk4TCO+lpRRrlvXbv++HLlyZlpbdeiD3MjS9DA0r3nrH34YCKz1R0S40vNLv1yvB
4s/qoa2DxQOEmKku9MipMOl9+efoC6X6e8OJVzfWQIee6K1L0POPi5U1LDJKWUuDf+FxcRVlVtGq
65Y0uo6jYHAW2gM8LGkH2v3S6WqmPRE/THl75EZ4WCYeEAPOzA905iIgV48I0irRF0VkH9DVb9lO
tgWmJb9rNaloOg9ewvX5RjGbSpv6C68XaIdOuF0kvjYNDcdX3milHipXhSwNruOF1gaqQAaA2OQz
bOOYAr+2Tpqlry9sITBUmujJA9NrTKE8AjRyB5K2kC5jyJPwDP+L9yi9UO1fN1jno7TooMNctdbq
cAd2gvrsZWDEmqT8ubpXCK7eBMPRvW44UrUhAxXalRgn2MPnhqGiduwoPccbqDtgjp0xmJa2T0WM
0xDalI5KG8U+k8F3+08m7gGdOoCsfYeDWz+ovMZypDQxyE70fe/UEZfWfMu/JUJIafBNePD4qEgU
y3kdO/4SZrth1MYRIr9sS84tTZV96HpoVmsM4KG6XsQcezrszjve1YbbXMK91AUTlUfgPazafwvG
zNbcdrkDBmiG1oxaK+/YWGwEKVpwMVsLPGhvqXONnmjL2WGJI1JpFO312rg2lmdQ0IVMExmjWWOY
7PK/HQF7yLDxa3tDKLHQMd/wY4eh0xYxY7Btj0wANOC6NaakZJQEDKYYP+0WGsrT0qllxXjqnGTE
hs2TIFnWFBASb/Hgmms2V2aQcgc8rQ6PoZtcCjl/vd6y9AW96pIxila7vTZpoOSNIeDSWkK1Wi1f
pvDDe0oX1oNcvmbRPvXVppqHWdWhsN0rJ9CC2VeHF/E2ZxwBaYBwSspANZlENhiX78eD5V1p8cmY
6Iw1o9szqCgGr7k1aw0eGh9AD22if6DO4Aeu9vIxAbzJQa2LlzIeIwGVm5no0w4zJ+74RKFTwpni
/2WdKWuXoxnjhsQt5K1BOmJDnhBmy2lz12YLVNmN/EjEwIObENYNNR2Oo3t3rM429YIdgOJqsSXK
TrQTdhZszN8JCvKRwkQyTZi+d85GwssZnDdf0HLcRtGSVQVcifqXGDCd2T8Wv5d+hwLUO001n6aj
/v72+yWumJiuxicb0Iz/XcYR5Bh3+LI0EQ1S/9vcaNYosv8it6gMUWPKb/mJb+voXWMGYwo7ueUR
vFd4nPly5EmsExO5R2cxns4WvmSfeokIQfYQbtzlpjQgJ6RyBu+jwpfDmv1SsDuslgVOWDSTmfcR
k+SfX1RhZN78cIsCsbuytEKTlhL8owHoWYKhTZq8ioWNksjAVweRJNMVYP7pwwdngd8O+2GNzARP
/mZpRGyuCfn5+RgrIHPcARxQQtRYCKMph+WK+K2XvJPew10xPXjm0Am0GEi0d3rBfROnxBcb2CqV
GBdjwvd24v/tH5XNZCNmmZs8s4afXYfwYhUW3Mk3bA0tKTvEs4Krie6YoWfpR3n6hjhjERXFAAX/
YVh0zIKaWHvr/bgG2MSF9tCKthKD5MQ/03OZGJI1UkV7qNCmn/ABmN8Z1AyXwEqbFWHGdcXUTUmv
FPcur0mYE4Ylaf7hr3T8D46SfZWE/8sGONuj6MHNIfv2m90MwG+8bw1lRDL+6jH7hObueOi+raTR
lMOUIkSGC5O8cmZxwC0IsDxfAj4Uw3ct9yVTOsfAumJUkYagTyNhDPvv9xAwY3ydYeZhpqa6vQ89
XlLPQY08TiipvJume9YyZph0SIC6BFuOLAbNtLsNdBtrh3oka1xFbmJNKS12BvsHe+KqPgGuSb33
kgzto6PtIJYsDmrI+q4uFv8xYmQENdmBBmW5CzySSeqd8q3biTMyXUY7nya4mRyMnUZ784gO0Zm5
e48ObKb66MAFHORNG0HjLwFop0etOfF/mD0sINoY6AGw1eDgWLAcQ1fHlH7GcPxhDrnWeaywdIoB
rDJIYw7t8F0DFYEgDkYVRc1kC0EhITORM3bWhJ7QiOEHGrLKVrIkHg2bdgmyEeo1uISzua3HsTy/
TqoQaffisvIgpMOsp/1ZaCzxTP2YKp56tU/QD6pTadBxyEko1elvQYongAR1ZjnB2UYs7S9dWNqh
YsuvwesrVnhLBMIFIHtRoy4MHvBLkaTQQR+QQqDTkgPohRqnreYXtyvUIkVJXJokSWKXhYBp0vXh
tOQ6VqD+z2eiJrZhC0jvpefzs3i2DH5PQJEekjg9T08U1SBBX0Q2xS2SODmlsNjcKrW8CBqJdG2g
pURxvQRebUHLNxZ5q8FkWfd2XoFy+GtltVrwpGqKsIsXsfg4RoL2+Q2bbVmSBEkhhOe/6sPu773V
EdrF1QBzzPOTKdyvktXY0Lw1KFsUiby6D29u6bi7P1x9yigkRVaKmexPKC+9dX4aibF+eNv1/NT4
mExJuJedcqGf5YDkbHjM/UdLw9aJDaJzpSMcgr+uDLAAl/ItLRKzEw5gxv2ebDZRFXXxyLG4Ruaa
3PS8OqTJsGOvNmkHTeS9h65c1B3TW2jF+9dfYUMV3FzGduTrdFL9Uv4WWFfcu38LFUB8pjoDVfMA
cIAX/otph/YJV6WvJ8668anCwQS6bjFZU0NitQ7zZzzRQPMjkQNwhY9Xr4cgBHnZ5cz6BlgtothD
pjiHSj3Lzcmszm6C95YSkTPKvko1rUttK+7xrSPiIAoGCYKNQq/7G0cobCU2/FEuL6j0FvDDYOUZ
rVatDgpNPkTYLZlxX1KSUc38Av0t9qNcUeG/DsJnOX2m8kA4+nKeCMZZwuB74CadUovXDZiYbJK9
J8NrPMMmost1s0VIG4rZjpyRwJ80sWU6OATyDgXgcADszIiEaSgwdGMN0p8ofJ0ahTwQePe+3IpQ
rcta1pgCfiosve9Llt1JNWtf1HKfjDpD9gwFW3IsjpfPKARC0IjlbQGouzqnyhw1TOZOSTttY2WJ
sjYD/r02eh/FOPOYAiW2GnwZCg4RDvRKzLsbGJrbSWb6bFSLUdPKvosLF1LG8eaApudQXs39LD8o
ExJ/MpjmF3gAwXI2lk304lBTYf6GkATc7EDzVD2JT6oqV/10QIRQvHIWZdDw8VtgAYPj3Poh02mV
9VifwB605mYtvRL0FY2eQ38SdxkenZ6vyhqZ7YrnxKOmghRH+6Xa+Qr63ORSyyh07gE8e+bNPbw+
HZEpnFo4k08gfKw7v2PV2QF943huT/DtrKRZGHhcHRx/o9cXoDfUnLgwkaZsSZFvowIBeTPya54Q
xx4cYbAt/Za7SWg7LyWYvinPQa9QfHM0zB5Wwg9dqaGv4CGwcCJ1GuUVuiyBcX6IQnIfHIa4mtSv
RaGmkRtSzZnzzMSz70yFxTdKDBTNJR1t2yRAMEG3nJFrbf8c9/ia91w904G2u1fVTdmSc/zZbrPf
KQUi4VLON0K9a5AIJB1s//8nP4N+km6qk6X5Z+9NntKwa4SYa7441hiBRE3CGY+ePZgm4dPIQXDB
Wx62v2Rb7AjB4yRT21TnxN8qsEmGKXt3nTq2wH+5xbBLztleqze6q6iKRCSnT47EDBNfRYvDsxhb
gcvFfhlXbYMo71m2RkgAAoA0nDCFvE0xjzXk0hw7zZms6r9y7XGPis1Vt3lt5z5Ep7Et9hF9qjV4
PvtquYybiRkel7clZ2ffWnMCSmMUPrBwztoM2xTHtGoFhE89LyxEgJOv/8azHyviAVOIxpLI9kFZ
q5MuDopsi6lxkTFiF5WD0tBZsfYI9NjbJehZsD5OxpdFbqCQhLoyTdF/oDcYgvWW41etL/N9affq
01L5GSlk5UqVNuaGGsf01fq2kbeHooFANn0q1VDwloR1C1fvtLJ5bJq6UzqLNBLvKWBPn3ar6I6X
w+17el1AfktJpr4LRN1rpWUB04I58I4OkNSH4ZqPH0fvoT4ScRC3Jdb/4Cw1bRkWw/Ou19cSulcQ
FnPf0zUcU9qW6/oQmwqz+uMFdWwQVAfN6iHcd2t7NSJh9lYNNjC73XVdLncLwl8TdkbDmFBrFOE/
p8WC/Ctu7dc3EdmBlrfMYGeVpWvl+hiFgc2J9gi9MmshACBPScml1XGExsQjq+nEFL0Aq0xAEtGh
0RI4wkcdnukooZkLHSLtA0NdRTrI9xEfTPegjaY7DAUTGaQwbZ+GoXf9cDy6bosnlHEdDad98f+Y
wOdTcNPSmWrN6D+4hzt1vDYV0+kOd7Pcu0S1fLysfBmftQwfJZ8xsioaU3EgzBpvQR1ge/dsXykO
V9qH6wmXmuAOFnpa0N1sEbfdjCksfpMKKP8STQVXX/hPFcs36B/Fu6uMVXcWLBdI66cVvXo6cFWL
8shkqwU79LNEHwSe9rOTZyX6usyfbK50Whwn26m6Cbu29x+ooGfFGRs5OQ6j7Qu838qb/VV+PW9N
ypjyVgwBX6+IvaCORuBBYDp92B8ywptghSt/nEHlMA1zdNF29CzGwx3iZ7hq/Oks+6CX6k2Ok2NU
ZUu1Emh3zpKnn1A67wT4kyG/yWYb9S2JH7AvVpk4HrLDS6RfEkQos9weSUJ7eG0JnsxlZh7/JUuO
PWAgLikzFlh8GiNyKZWmOCVD38Mi/n2hVNySVMQA22uNs53FPMnA/LGCaRG+NwIwR6aLpqsJQR4R
dEESqfqqgwdkGLxN77xEa4LyVu7lIwttcCO6TUsOH6BN+uxPTTdJSovAhjvVLkt71n+XjS7ZLvrE
peMlzv4YJUXEBKVyHroLSFw23ABpfkzNa+vYHBI7U0pn+zhAEcpWFWSG8bmwTRov1c/9KyvDGENL
fxczNIbmqgqWqzT7xasOblM+Nr3c6Z4xOGfR5gSW96CA3Fad395Rlea+WbckoovRm4DH6WrC7tsZ
QywCGIs5EWdrNB09wxWhwqtiYpv8Ifi2IMxyIIdH6UWj23EhmxsKPFvurEC7AokWx5QJm7EGleTU
CqmMhiN2XUOUrynRkkFnH6mL/Fk4PC4XkQBLg8GOms/WQT4uyJkd37uxAmlUYr3ayr72q4Pm3iQ+
nqG9L02oX22xIRXr3ipJsGTIFEwKcq58b+MYDNXB5meA7vPXN63f6hWHM+baM4/7+3pfCOLgu5lu
viNtho2dbAK3WhCGgwwHLPEvK3NZT1tyCdScdtVCEpn7zU+vo9rQTlUSrneuJmsFTaVdj+o9r7TE
xxpHca8Le/eQo0s0YYbClmdbrsA5ZOUgFPozGt2IBVyWruavefy2KdxuOryXrEUJHYEboSyx9tUS
BWSFNvYqGD3LFAuLz0tluoiSMR+IpKFhdCM/JZJh+MeSwE/UHuQabZ8Rj+yHEuDIq2iFz1ddXVPU
dAw4sejFj8utRDRb7b1bupz1u6PA3wg5XEJZTB+eVF6IUIXPC0pCoYuNW6eOAHcwEZ4cD3RhlneS
wpMJUI1kmWbjBnwppAfNHNNDFarBc6MkJNFSga9vkLJWPINTgNO/rHMyCRfwRel2RsE6EJSbBlul
b96J22QPDNNg+a0/0SdfUYfZ9JcCtNUugSvew2QxqWtgj6IQkoLAorGujdTkq9JHQWpFYCLgM1aP
Er6XZ3Lz7faPvFP7r1TIF5Tlpv4fqqdvLwHjNfyExP9s8f0+LsHhjzkbnOXdOz0J3OoTMe6cBn7X
s3GONm8dh1gsUHnEZ8iRbR/MfWRSRKldt3OzqN16lePpCW4AVQcP5gdz0iHHI6TnKTsriiOM+bC9
hOYmXxG3kC/w1d/zcXWtDwYluhEQjCbCJtnxiL5/VGQtkRps8fkjcrDDxzqnBWh/qfbWNB2hyNfj
lYqbKrcXVcb05vchoSecEWtQEG0kV3zfW0dXHP29GRt7AsJQzN57kRmIQkscmafGt3UYki/4pngl
cvp7wj149F4F1kCK+mN5pokJH9Y5XVcGXTfOkO7iGj4lI6iRwRBn9ekCRp+WjJsZeC1hD5AndFhN
zCp8rbx6FrhWxN3L2RrLZk00WVF2nlBtADHQIIZaSY+R3mJM8EmVwNSAKtmLtODWFWvHHAUnN8VG
FYOfejVL4wHjafDqucnE1J8dDy/pRf07YpazQeouD4FZ2Y29OyBOOTIqyrF/PM/U4a3g1G4+Pxdr
OHks521vpYrLIJvb7yqHywrw732zH4OJHs/COW2iVfYDXqMqQl0jwd9G2AdvPhh+q9wx9A1Ja2vj
3Sm3wd58S8lYRmy06IntISK7ncwAL8pkovvYsMdz2xmyXzEEmI+MzjvAFZ8NNQqJcu/+ZE1jYq3e
kIzSv5WfoPRU9xAFASTN1ew7HOCoKI0KHCna9zeUbIp5KS6wHi56UlAFZXkSOk5QpjgVwGmWnKoU
E+qm/RJm+TkPS7gyToc0Q4O+ESJtJOAfV3c5mb0a8rTzZfQEurktLlHar49Ejy4pAG6VEF3mEP7p
B79nlqAlyaHUuwKPMa08aPv0VC4eUbYCjLkCP6ZB6iJV34JRGSBqbCU8R/5XBIUd1UxlvzieSok9
lwaVg/v9vBzoXiaog6L3xcweXdyfOeA4DWPzyY7HdVB7prO0fEG+OtFNivMz/0ETcnooBN0zSM9R
WG1ALywhJkBVYnWfcVfwjibD18E/9DVJhKMcCiYt4Fk4l+wzoLuCStMA2hw5LeyPQAWNGmyHVreo
489wWkGchGs6kVSUQ4qkMkWJi/29TgQ7zrPp3jOdynkVA4jMkhysQvcvBElIg3uUes7rE+rNyaU9
rLFOfVj44TX3sILrkxHCOoKgG3/itHoCBgG0tE0SH3ipamt9ZqugVryJ0PctNG4uo0U8SsL7bvxW
UgcGIhTuZz/iL+G8g5z3chZvs4LOqK5uNIViYwuQYGWtqvwUENR0yljS4ZUn85Cr+7Ni1iPpQiUO
8ssIbvuT1xqPwfW45knW1K0fbpe+zCjFNEx4LaEU7Fy5NGmTUAlnNCRvJsZohzORv3+qikqskSvB
QikEOG/gMoTKHLf3Ket/YH5YQM3nf3fF5yW/MxOMS6d9lCm2FjMPy/WyFFrpKPZurCGRTmhy27yE
p9rFotz+izg89gXepD75fofsEouCJicSv+6H9LInvf47vIH0D+qdv4XWMmxbYgm990iHNUEJK/lD
T5/MA5tJJxxRWupzfsXo5cwhb0dkJ8U+be2Iw8d/kLaVDYV02tyyszRUKnYm4FuejJSTgLPNB/Yy
HUt7hENIKsYvrbbEBRgt39OxUWozRJ0i3dc1prhqo1w3ebNHDl0fe3pGDWWUqTwDkBntKsuxiwFx
DWLILonysBJXhkw2IbMM0bArJV6MWaB0PD4PZX6kajaCYaPqD5njdc+0UmHmTuQIdJYrcawKYgcl
s3iHg9Bvrz0tg7mQ8AOI1AsoBDbGxsZ1nELojm1pD7ERwM1JSn4xJy1dnPNScMvZzhm61bxQYLGc
mLAvUC7NB2ZBS/IoTdetcraKIGP0JBjwpfOdbI3Cz7ichju6zNSrQWg73kOngFLskvPcwIBTxhl0
jnacnMmzZOfVyd672Cw9Ggk/wQJVQXNu3f8uTxNnV+GefBxU/56ub3PrM0iiq5xP7/Hcl5oNfaIw
xkOxKi5blP2iTnqsc1kV4cVMeAxSl40XMYkt8LOeTyHCv6YTd1/XWUFR0yy60mOLpHnYPp4hka5B
LA0703KnCpTcin9vPqAAw1mvc9I08++xtiXD+w5ojk3LT2QhaaJgjTAady3SDvah6HIKnka5lYWg
PggknRfmaf6IgO4WLa27nVPYGtHZ+pC3w5TNgoXt+/lwlkZ2qVjFIxCv1El5nh2URbFF4OX4gJb6
2i0QYn5mGUkR/rIReOZ68DtNRP1fG+tKNx7epRy0hZXaKjItMYDGQVLf3oPwlTRcG512OalFs4Ai
gketadI2y0XgeO59qR/fdxCWvwd9ezAc3uUliVEmf65YqHrdno6VIyNy3Abk8lX/3VWZjGXVD0qv
0xU87rDzMbftDtyFTadwxiwKkkHEW8hQZIiV47ruQBqyT2QDcyCkcULLNCShO5KNCMlmi5EclM+S
XUDp2siO8m65USg53A9XjENdD+phpK3dOwgLsgAskpwZR8e2AjwOCQWzWv9r7s3WeUMyjEHNHREi
cozaxjewfhw7QoOKuKY/J4IogMpDcSmsYgsO2rCrXWjw51Q1ncDBroP/+d/LBz8/MgFMN+Y2Hrur
RjJ+YapGMB6Nvy/oNORurYMYfTcz82/M8rX7q9xN1CRE3QWeH3Ds9uIFveoT9T0zPU+JOJe51Csc
bTvoOj2wx8W48VbwnK3x/d8T1CPGrBxfp/sZ8tN/WnueYq3D/nwwtGrmG0OrVnl4uo5SLX5LRsZU
mja3Da66S62I/SILe1Bl90buisNfnH9osWNMA1zFN2Wkf61Xh1GhsrKOFFnzX1u3dYTxMslxS6lF
Nr7PYSTIuLR+5LXCYZBELC1LJ6oonQ5vBZlsRdktS1Q9t+B7c/GvQZYB9Q1OYFeykvbfKlOnm/Wv
Zww0jXywVrw4vOpEBh0IKU91AlEJ2iZahs0ViPvOsNnTnt2A9+woddYpcbE1hFQKBdREb0Y/U4SK
a3gsn3av4Va7f36xOabUesgq203rCDnZ2vR+Z0vsZu3xSqLIQ56hrR92ENL3KAfzs69oJm/TqC/v
IkTQWfg+pz7cSQR9gXFEsul3wOLSrDqVR7TurQM9csGxAx6fAQFOwbMREGsL70nFfNXBHLcDz925
VAhMQqakzS1Vw+3oqa613vTskMJJwziQJ0UVZIGlNuG+jJyruVF+CfIlcE1zrnj9grjmazwiUMSd
hhj+J46YOeHWnzIO+42Sz6t2ECuuLKMavsn5fp/XZACPcSM1Jne3GOPEDLpWczVMdESf0x8xXU8O
TYZ/CmRkiFCXJ7a0V/1JS3SezkzVvt0vGQ46jAIZbaXMi/ov5oulImYZxZZnW2PHKGcvLZArBOs1
zANnHSSuSO5RE1RKrIEQpy9ZJSBrcgvl56C0kHsSQS3V/qvAHpibohtFD7ihmwJwJy4CHdLxsyTP
twBLiJWBOxqh3Kawz4MnI06oA1taRMalgiDej712ZTPrAPoCkJroi74ZFVvKxc4Tesjn8QRw1okw
g6kFvglhER3Fvppfqj6jio6ya4yx5Wp85n39BRcbpt0Nyzru5mjXXodFWpcArfSNAVOwS1EWvBeH
km0Z+fe7Ifsaxcw/l1CAiayPf+SFyPOEtKY5XJCZRc7zTwCCbo4S+cj9kR4b+GEN39FfVjoTgzM+
VOgFvLxh4XJDHLeOhCbJJgvSeY2Dar23OpbBzMkJp2OHwTFEZIzLwmKtsuhR/ecwqzxKcAzs+zE/
72elwVvXfOJG23zHVJtWJLzmDPACNwlmI84loetcc3/6eFb4tBt/TC7TzhIMYF2zJFpqYxJBGzZZ
YOYYSOsw3kk2sDDNVAk/9xNmwULUihJHyEvVUEM3k7uOTEFaG3aNCCF57rZ9ocQCtvwt2Vji9Xhm
pn6qb/wceevrMeDBcZV/Tm/jVGYVyrwLSlqhLUideAhg5k/Dqe/G3CCaj8ta7TQqLnabRqXVt2Tm
pOsMXnnPJuTY7f4+RQWBAH7uSheXgZinyb7BtbqJGA3okNMCZeqDNyZ4d7MGnarvFXALBM6bubse
KOTmuMNR6ZHhkUHwtWUyVJqNOmO8TI+TfMb8dudEdhzcxTCqO/ZiSeoD/BPnaXyh1AIF89a7ZjAI
07vwF218bUCZnmYybI0MTAd36WVA4yGUcyMU2jj0E9pwH9jk5L0djIa4mwqyMEvpqwSNjjLJloZM
k0w8tX3ZjOFS++WHujb1FL/z7+3iEEnCRPDBlGSxhAz4Z3XnymHKeFNzbDTthREoVapC+JhwVp2Z
1b92DJxPBi5s+CSyZMCTkrxE6CK+i92y+YQd2UdFEfDC8kiVOF2aF5N+rHvYtxfRntrIzW84LdNu
e5WCo0F8nRbATdUTo860ZwoIaoeQOzWK3LKd4EGRHHIWa+3Pi0rDh8rCrGqi8rkpveypcVLVyzX6
fRnH1irrRkwpuiBsdcxfZs1+M7C2pZpLqbY6a4QJ5mCAphjB43v3kFRQ3I5zHqOXCr7gnoft1FNv
4Y+hdestaNUykFrA/UySPiX7h2AJN5OYAWAcxZf/QAv730KEqcJ6+sxTxbKrC4qthlDLLl4EOcQX
i9u4GQeAu+392YYNrF1kYIB3jFb8QRqkd7m4EapEtE5+x5cusnkftcpnPTei036e7g2iWRGEQila
OlX0Dp2Ia8LVtPLxxCO5NPrArFbRxdF8jS+q6yHxf3O3zXvwD6CqrT9eoZPtCIFJ28jk1FXBDQLV
T4fP+V4vsuUtMmEuwYtxniG33TvlTWPyS9swMFxYYNOK+1ys0imJfr0DzSBu2RkaFtkh0FNxKZob
coGFukod4GmdPUyqw6U9XQXQbAxB2OBYSn8/QXs1SJI+cSUw0KwsVY8MDrOjvY80PsGwSsW/WIRb
QzEGGnHfvnPXXtUgzN9vzMvKwIzKDpDNtm606x+WwRMTmz5/grlFmsiXzNGa8x7VGM2lT52pa5gR
TESX1Q1J2WmszVLN392/xwLgsBEErd2h3nWKpoO10amzlZWBPYhbZL9gsLv8jnJ0JVQQs1X7Gr9J
a4KpCh2+Xyu80rTAQkOy15zLIJBL4j0/fVDdK2Hzkc9QnQasRVTGisEzPUaIq+LtaI1c+m++ftFy
tCRMcs5U3RwklrLCfSmdupexFxd8ZmAssfInweVWyfzQVMsdlMgqM/TCNU2oW+ZvcTMAcyMyPGQI
yHZcY1QzgFyixuLsOSvnD68O93E5R0foqAi33IJIhGfkgBFvC9tCIjbv1xyB3054KRfqJbcI7jhQ
OQ2wbZ7RNXks9CeBTm5YxoAz/1fg50163yvhms/ZVaTt4xGh6XvoCX5FM9IuiNo7TOdwEAarO4/c
6lE0ISw1Za6Np479kIXRlTjVchDpbSb5WcBgNlFC3FjhTKKxv1vPvX4zLS7HXR06CzLXDpTl679Y
bTM6Wy+Q0vznpTp7sn3rXYyZuiFf5uff4eUtlKNX2AD6R+fUqlLPv/clUxuZkLaXTwilC2FscUJM
AbdMY4TAMss0ZEGeQcDZ4AW4qqRXhII3mSNgYJ0LQWfOa8zmdaRftJXXuIrbY/K1SIHKMZ2AvCCR
INGsLkHY1DM4hBmSENBHvR2Rtfg2oO/uIJOYLWuQLR2bb7Ctf19DaSW2wsp3w07pJLAigpIyUiCG
ziTSDYs1r7sTS/Hu1/c5Qh3v9OUBsUQUqZHI5+4XSW9Jvbfx1mnx4eDpJCiZgYnH1/FLXKeEsVpv
IQbWbwMhJ5LSEf2pP+rlv/oBb1KaaAE5LaIEI0ZdIQrRgtqr3GeDDv1d9HuMdxbjVySY5Ehxd4pF
L+mTxyoEp/x1PQEvsyA5fI6Yd/uyErcrA7+B24dONNUFtuWjGwe5plhMdxqLPzJQb5lRMVj8QCmB
w/L3PxsDpVDOmoI1D1lCS+EkuHHaThxoITT9sCBHxRbuLqgrm8PTCWmfVIXPKOYirQ9Wx6vxJ7vR
TX8p9wZyRpM3+LoC5dia/3FYLuVml39Hvk4HJPqHGYrAwvkMVMAggghMDpvyG0/FnfVTDnTIrZb3
qq5dfWGgAVwM654AmEXq8TrYLErOB7I2Jq1cV6Uz5bW6SgoW/MhuF0Yue+hTIrxvMHWerOp0qlFI
i6BGF0ulKPmPIGQGIXokQgDuLdxtRoIJZyV0O90RhEuRCQnviEThgZINqjdny/8rlvycEHZEHbcm
hBISmLbB0Kwy10wg46wnsjPvM2Plt/rTsVDOQaItqIw1eawpo4hOCQG6EuUtqP225gGn8JBs3kok
dKKUQET+VolNFd6Cagn++hXXPhmnlOnsX/ytQFRWcUuW1dCLdL8CBBA6Y8cxbzk2xvDycuZ4umCB
KEoEOX7lxeRod3LoHRvXms3vWwz3i9f0hlJNLO1DATBYdnCM/3zagVVAokrqjhlDD8aHsgYMKj55
WpLpXOg+U8ThW3zreJ6ddEazU4ULbTD3iJHCuYETcyPas1bU9Iep39pUZmMgwhRWlZce7RaMmUQp
TBk4PMK4IIp33zk66ysClUmaPJUfgVjxCmys81j0YWSACEqTmR4ABaXhSTLMNpx8/SbZ1l5mmEFE
eRvnq7+sVvu0uEdSo7eAew3LZlinFw+A+l8f3YS+SX1t4KyhZ2DM4twjjI1arXFY2JgVg7triPpQ
Zlxp6LBHwKUvVyRLtKFXnxp2mrncZJAv2z6CKFwn3q7cY/HSMJHafC7+Z/dV3EXiqKD7TuhJctxP
rWjFAMolW+4EsQu+jJwW+nYcxGyxxa05hvkgeb5W4WxyDOiKWZnTgxNE8tWiXWjyRvZa0ZoMu5U1
JCDCKotlcgysyLz/5P1RtsUKTSFzcvOMr/QMdtMwxsehOl021GHOpwyKRFOGhF22cDi73N4Vw+I/
6RBdUfFFOCfisUpe/y9XGNZ4FIdsWl3diLKzc/h+a4ZNKeSR4SVPCWi+2WySTP9+2fB50gLvrJaT
9pXV4d+fsoN/gQGs6nF8lLiP9L2T7RdPAohnTmz7JM2q6fqjcMRW6FtSdEIELFi+P9JR9xPJDJn5
xueNju6xhWqwCCiSsjc2Ze6DtqLgkTX5WkKRfGWTIEdo9QmosmcY2Y9peD896Zjy4Cke8AdMfVHl
avrRdIIR6kI7WVUMEQZTXlpX50YNIIqjp5zc33JJrVhyFveWXzObjkMawfEIM1dQRx+AE2lD+mIz
r2AY8R0LzUdVA4RMUnJOE50qjTZQJMkPvwBXikdRcG+8pSq93GGukMZlSPZ7SZmMAh9RDEM7U3P8
F9+6I8qpWxYYfJ8ysQ/3eo70Ej6nMh7jehWBbar15k8x1H19mZjQjLM3+DgqKft0/8UsGjSfa0OA
xEgzao1r3PFjaITn32x4szvDBkl/mR2AdFav/yGyVO5hn0A1v5bSP7Emprdlq/mLRMRVePRJTOIU
Ex9+sXyiUkreAsDX7vWPxJu1kdIn3ZdsuXwGLV+FVvw09ziXo9ebT9kg6zEln/pTLTIgtRZiGTwG
Dh3+hn46ff69167PlhXd8fZN7UiD6hJzpUseh3OoyO8mNKbhu7jJI3v0obzXO6uzcrQPniKPbViH
3y69JvX7jl/9KKjpgGsNufvmG66+dyK/TkDeqJZruIdqP6MLPADCIpl6uraeUymRgr0Y1J7d2scn
2XeKiBi/Mz2k6hi5vjZhxOVJdyKH1HMkDzkvD59EcsCYWzyv7MSgSa0Gt4ZdpQHjPBXwZT5+BLLE
/dATHFOIDeGfJn5u1F5K1zzTC1CoKtiU3relJuyXz4L8QldrUMCmJMKEVEgsovWsa8Hauz0xTrLx
ujnDCpyb8G5bsDt+ypFhVnkN30rb2Gy6+PV0cz4XdgHzLxpEYEUdw9kL5F8tD+M1pD0iAvTxZBXR
WRTBUezh2rS4ucZf+3Ba9pqGRFnnKh1LVRY0rPqxeY/TqB0DYvvDOFQVqAdhPos+5aun03SKgkQ/
luHZqA1Sg9fB08dY+Du3JL7LoukgvIPP/gfDMt8gP/QUvrcw8Wo078dmwekUlP7uqzTu7lW5Tzd5
epEOi6M97yqxNLR6kHVPGcb8hFy/IeXRgN1qetHOmM/F7JiLlmrXgZwlOfbSWFql6Ji9Kt+pQ0fC
UkxIbjOSDk/9bR7TdWKRs3VYdjx0V69KE09ZOESdsJ+nmFQ2qNgEQ6BC4vVjqPG36ROmLZCeU3IU
iD+MdUp7UkFW9zj4sbiJac6Wd8tTC9iIG4F1GgrM39zkeXj6W4Z0ryPC2WpH+2YB5oOb3xKLtupi
fhVjFXsxOu0QARkzI5BbRy08KN5SXf7HuCJDDwjOvJNBBZYSYeU7XeapibNbOM2m450sNzWbtwtk
QabglWhhLU+eeDByFiv52w4yCSeEoUdD4jatK6WoRcKLrRsymroCHHr1YfY27NZQQJxOej9gLiZG
klKShvW8pbrWy2urA8fb7BVCpx7qfrGyiCPeoLtBf08cEF8ig3LnfO2/p8R2DNTJZogqDpw9QQuG
2V8eG0Ud9QJXu9cQ68hygVdhPRbBAvrRv2jMmOlJyE66AAjejLiKPyxcyGcC7C0zLL/ofqRYot+D
0EqT42puuBLELvg39ykHNSzUbS8CtPjz2yQtBqvAKjLYNUmCnX0uhbSmU6TnZsS1mK/FhxlpFMui
zy+KCioM+HbET6Z2o+906BxygqjO2asIwto/MIH1LJeH/H6Om6ih+XOAViKoEI2lN015SVjCZY3k
JHXHPz4JsdC1sT4hOX6dPTpB/BGc5S5+sx9VSDQB1ZSeUqTumnj/Pv9lzwKhI1/fzaFTlPMR8t7q
Eagv6oZ4ZfMdt2TOermYVozWpiux7cwZDSPgAkqmYIe8DE6jqqywKGb3kbRNfEmYX89bE6Pmf7S8
X4PWnDqvl70Rw/MI44IzbufkJu5QbetDUD2J4wNZ3drwoFv7ycKrG2rmey1F1fImEdFXy/WDLgd3
XHGWgguzZdRG17d5zg7gbXZfBwH7oozq/bjA37h+kqFOtOGG3LP79YcJSFreex+0EmH3vjdkUHtV
H/sAR3oAakQHufcJ0m+dKZKmV+4QbVo6QpgCibw+10f4zqOiZN6oURC+XAl/iFnZ+dBl8tjnDiHT
h0JKKQ9Ah6REFRZMyJcq7/5m4EiZayvuaVIM3ubNfq6PQuMWA75en0/ujyuESpjt/vtwmzmphEP4
MDYpTLBxEGdkU58a4Vy9krKgZyj0banjym982BlnDLfAU0PViRHqhgObgHyC3K9toyeUQB0QAiKO
9nteZa3lHmd6qAuW2CI5coI406a5m9abmgXJEITzPlnme4YyiG0jMpkacEecCDKzqwdmcpKfwJQI
STYo85LTsm88ZMVs5L1GGW1JFPShrfLEJ4O4fSHDyOmxz6h+AD25Gk7upMp9OlBNQmgHen/KO74b
JpVsizrJ9gg+Dl/v2goh9dy12KFP2l55eZ+ezBQ2Ea0sYqntcijN+nU44bAlBgJTwuFT2jk9mZ0O
Nd5dKvvpnsBIIbtd6V4omPwj8FgGRdT6GlkdF6JoNIRhpIgEeY405doAojdVMaf8Xf+XZVC1KiiL
dV9slY3PwyCDZuXOrK3dtDb9zcNl7caosumddOsv7nnCW33/G7iFst3nm0pMVao2qUIHcic33C0i
HBMI2KHnUYtz7GEPGeR7AZYcY+y2CgGO5Q680TCXtCEo6qDubfYbDhtl8SwGltrcB/lrOf5gK7M0
+TrZGugEMm6USvbT0DHpoth4CIoZDuRdzFlDTbscb1xGrhhNmbGDK5oZJhvcxQaGXoI7dOwOkku5
3vH+upgBLmE3G3Ld4KI/SxQqK2Fc7qjK+aoiznI+pravYBwx78P+fKRczWr5P4l12cuk2TDUIR/o
5rN1ARtMXLMYDznxrqws23ZFG8d7v0pyVMCZbZkSt/BoFysSfvK5srJ7OdFRBYRgGgR5zHxOGCQg
pAADjz/XMt3tzkaEOwEYjB/JdiTmmZTjKOWTmBYYS/wtYVvxxurqR8qhBfWDithZPZxpn+b822FI
r10Of7z8+9C64whlmISsGJf/cNcj5ep4485s2ST72H/fxXrmj8atSreSsY6lL7utU/nzhowvLrvX
2xGZw9iE2aoK6AE6l4WmAUPv4jSWfz8rZvNtIj2a9odY8401nYpERIjjzdQkbwoVBQM3Z5+73YxV
I6aCyNBm8n3bKo506kQ5BTW+AG6+m+Y7ztUn1JoqbRxxJPmHtu/o1WJeCOzkeguNSy5NR0LuTX/T
HU3FWVjgKPN+2YUS+GjaGQlz/w5JEevH5El1NABCasvsX4izO25CxUZCph+A+V6YEScMkLUY7WNB
OVNIivBfFiVvFsQjWVpWxYug2HyALEJthgbUrEL6Urk7MeLzCNxrCeIrxky1aDZi5YlC24CHz5s2
Vv0vbQjD0tx/aEHxDOXXE7NjuV5NECDDgaYQ8poefXYwhhnDepND2/O30JEY1AiRDKJ/hZHT4Qr8
09ma+rRhHkTxz+NdU/QzGvrl6zv51QYLz+zpg02TKS8yBkz5yU47Y1Vm8gYoaRVu7Wne3XJaOIuA
CtlDCAMn1oPEALGU7hYrnsAP+208kttay+oodfTnSs5Kc0Tps4iziSG/E/xlY8qlmc/OeTQP6BKg
KVDtpjevFwGQvcQCLWPY+FLgy7DRUHnuRJJjKIMd097zp1DrwUsIZtqgDlOTiGq/iZ4n9dlb9jIm
WPCxW2gkZ77ZdadMy7f2t/HpMhjjjZWiryssnm8QHFlq6cyC0TQCKtOmkfDc3BNmcJypt9W7wG5K
hBokMAVEa41bb3lCvGYwbN8VDKdgIokOMGJ/KJv9r8uC4suRpuhqWZRcEnPUqeumYn+4Z729Orqq
kgwHaXFdquxchFFoBsR4KoMiwKIDe2o7+6jHDlEUAkvQnC4IyWzQlgvtvF1kQ/RWGXFGcGOJZm9o
rdst+aEJEW/kb2jHxMtnfcy80TXuAt5XnEmfuf14V7TsCLO7bKU3Iu0keDnJBzj5KZoaDIVBMrF5
kLzMqXKrvZtpXgfWh7KHC7mkYZfCGAJf9XrtaOj7zlSDr5y81MxgP59/jonePXCvbYccpB1p1QNR
vDO5ZMkkzbTrkvEpouzNosJk1WX6AYKWa5V49SG/+idz8Bmo2QDXHEctTavGn1VPvEgWS7rrSIeN
ldX3MvCWK3lPmiztvOOYdF9WBurxdbFeZih70sB7M9d7w2nZ9uWO/5YoZ4ealW2JQdG8KEeu/NBO
8dMUvaX2uj/4RWudXjBsUrnZ4ugTnZTqrKw0Vxh5Z5OiSbUD7yKSkMh+WCa5kfeMSV6HV09CSZgt
W5zSSYz53WNc/abJATTRjBlYNfZ7eV74/93a72EI3vElJfJOS//d3VXjvlW7zb+Y5zgQDI+eUNNn
ico9qzkwlp06tWHyoA/iIRI4flZjy14c7/ak2nWWAa40Kw3tAN/hzkEWfnv4tiFihKnpSQeKm98B
wwQyYpGHq7Hv/84ZVjk9GB0oEefs/n+viR977SY17luXkLDbVVGpZnTfe9QZcb9d8wTMXw/tXKns
scYwNGzVs3SLL/mTejZoaP+jolQubNZv117KMRmirBIMH3gj8666T1qZdanRvPWThhq6BkXk1omK
mnLsD9pLEmM6/SNth9OEY135ah5Jf09h2wRE3teJ7UhimOClYynoO8wnNou7xtEalUUR5iFw3tsr
kbRTN7wLN02R++Lc7W2sp0hkE1N5qih/W74IF4tgf+LoOp5vB1O5TpRVr2rPmLAHnBMFpuHuh9gK
IArAMcjKjPf1MJdUdQW9pZ5YaM3wNN5L48MqC0xLG6Qzdq1W0GX9Tqr6B1IKrUqaMn4n6f70kQRF
0qsEOGQ/0o2dNNJaBWgthQYJ7eyCJFktWSEqXsxYf0Vo1ecY+Gf7rDca1l99qROwUjD49Td9EWUu
dC9FcXUrr/scBh/hnHGtXXj33ppU+pJlINmoQBnPF2CNaPuPhcW13c2xck8Ljqa/rEPbHmMADMc7
c/ZwechyJBld5oxuWJjImezvtr8ON+5sx8EL0hpe/DPA/eD6f8pIwnmo32uTDsNitsyx+7Z9a+Lm
AtkyScPp6gK0yi6GM0qqUFlsiX3IhxfhXEERMNp7qGpjjxxi3vNsRMIinEL8Om+ITyRwzAKtXg4u
iu3BscSE+o7/jBFIpvZ+exEILVdNtfGQef9WPd1Go3lH2uMBCkIy2GZS4vgkO0Q+c7aN6yEtjTIa
NrazySk9qx9aBj5kpKrQlSIRFxmr4w3kluvDDAyxCaAbr2ocoolCj6iK8ni8g1gPvnPbb4bOeENZ
Ppqz4vR64KFSfsZg1usvYIg1zGWL6gfknNsxA/yZYi05dibYfBeREQ7onFxsveOmNx3mlguaavde
GOSX3NX8vNx+Ee0OKmYS3RYRcx6FhJrmgMW70dvY9mhb15bIq8shaXoxssuqBX7K+gimqHpYPLwR
j+cPVjVauqe8dWlja9smFGBHKpZN/vJ36mWd+OWfSe0oUcYAnn+rBRkmUg0dSOl0CkCTcgJS82lF
3Yd4u1zYJMQjV4/A3WbzjmeSv9qEZZCHwVNvQt451BpyELEOrJd/gSKZehzZbkQ+kdb9Pw8ezST+
AwIXr+GF9PQ4+wTI8Gkw+kMiFfNhv2El4mPq02XzHL37OtP2cjpCuwspaf4hKM9XWy2++7EoTv3r
o9zYT3ombcPswpJa1J5iUmbm6Fgi4We63DuDH5BNiydwwKicRyywGzlE0xJxfnuq7YS7tf9xGJkC
er56zuKdcY+xO7SlibSqgNRpgYoVL2vgsRBbp26wNxX8n5PudZBxWRe+dEJImPq0PjsdzgIyfAvj
1RLmWrc1NKBgWCkYGlnsgNgIiAvShTiYz1Ry6GSsPyRF1krXv5hRHX9vxhPWbk0E1psL6mDTNHrq
1WicQbOyOudNujQ/AHyZJWZ4sBf77Lk5g1LHpvH7BGEoZr/5BlZrUK22yafmG3PFw02tox/XiNN/
mvd/JH4seoB6OGb3qPyMgh2UgnWUoJUF3iAI//O8AZpxOJ6NzPX+ULi65J4R2Sxd0f7oQgFtuvKq
Ga3o4reqllM26svgBzuwMLbgSbJrYvClGRzSUQQ1BV7OoTRYwNkRjDfHpbHDaMnLzBgpEt0TputF
uBYx0vsQnu0HVIE5CaTVk+YuuIkmFMddReupItYxyIDJy9SWUe+wqRpZpnvIT8FgV2rnnooH8LgH
7WVI/ddhE6lJ/lfwzxGRV7nU999LkXpQp0EqINkq1sFbzeJsw/9dDeAtldzVafkcJvzIJbUR51wf
TmgHli0fQWyv5XJtyvB0BZDV4QTOJmcUZC5NE+KbueQ4iB7ub+WBNw4sQ91Pw8X+akLS9UTZAr2s
1pe42H7Z1VOTXmkyY5DpOIh+ycc+PjB4QsUh//Rl9gHtZWLgalqzGaI6LODM2HvImwG3ruyLFP3G
szrrX13aAJVANYaUSLR1clixPo9V7A94kVynspdebjvpaQXmPejfnPqxe5ko/iELHjnx81ykgl0z
dKpgbadSGWRFuz8Ax2ijxSOzmpRlrM3TZuYJ+zyp08D1YXHl8lq2niymITgWF8bBk8EH9dSAV0un
8t63gEpwKN17yHeTNGiykWdIeTQSO0QzgourzXlJteZwwAQa1bNUJfBjx6zG8oZwbutlzt6buYUQ
35NxL3pSoBe6xLhDselzrE/LvDHluJuwNnD/zhuuM4YCpghaGGgNZ2v/p4mGVFYPoqx9wsSQCmwY
qoLrXgOO+XNV3DBM+QPZGGw0yFlXYRmLtcSS5S69QXOQh4Ga2hA9g3KR7THFpL/i61qOu7b/+UsA
cMMCw/C7pwPRqHrlgmZjvXwe3njK9KkEws0GpNxSo3zWz930lJoiMu8p/SolqS8BliFZFtX7u1Lf
J2vHYL6LEYHMwHpGw+13BMYvHHVqCBZj6ZJCh5ce5tDgt6RPpPU45ZvzfXP0dKdWsjuIj0oWJpZ3
crssz9jACCyH3n4CindX4dzjDi+I6LDNs5oR7ssYHkfNu3xDTmEXbkOHztrBv9fhs/xomkVUZHlI
9h1C3RNr/iIEB0PToBDYiPEPrzqPS8DZMB98agc37G1v/bU53J3rw/70Bd9CvR13icoyInd/el/M
r7Au2ORtdrAGWLJV6TA0JQRI4w2azJ1uYYS8UZ0LG6075GGNnB/O4nSMJhA0lGPtdZ1wP2bea3YQ
KT+VGT0C8aW8qTaDsjKXjuLnPVKCgfEDGrqesAm31DqNFgF+EeDwyiV+ByM6e5MWaS221TmhBNxe
jpf8eie0VOLksEyW7m61X12qitosXzXwrNuIJV6cYSIl68xtn1Ly9GKEZZaPkXB8mzQnwar6U8Os
9DpcAdApwTiWiPqYLpytc7f+NAfNzrsBSqPzaLLTW3WD0Pif1wuNL3jtGvHP+W6EiwilYQ9rRecO
RFaZHz+f8uzBL5co7YN7wmqi8fX2DSPn5Czc1MNl/JoIITqqYpj2PUE6JLvNOvTnBkFeanxKflZ+
iEVLFG7icU+HA3VPjhb7EjsOtpFijKElRSYYkJiCDNyaOp+l8KKTYeYR3OYI12B4gGMyDrGmrtOl
v09zt3HRd0ylWXQm6SHl+Wzg3T1Bv5JBQnKdzya9fE4ijjrdubrk7JnDMKWW59BKSSljlVpkHUE2
mSxpw/C9r/sEHbOuWfMD+bXKwoSHhndP4WhgiQ4AvwjaYkZjZeR1yjEPB+zkcP0ll3OiQkMv95uu
oiwZNvQzcfkZMljix2DlDtFifzclyLycHBJrESicfHR9fIu4XJ7Ggj4POB2g7DKYgo/K/aFveilX
e2S+34skacBjQYtuXrmhsvw4S8NjuqtB2LyOREquXm+BNQkFg741aNQG+pCYBPxyv/4LgBI00bgH
YFt9DddJpUJW3PKBGlYywdYWpFunnJ76ZxVgzrm43SmjU2ELdc92SOUZeRf652PI270xr08MYRUq
kJ3Kx5XgwAg3dg8kgsJ5yWOsRObzaLPU+o7bv+CFT0ekRwWVtT11r9caTUV8qU671LwQWAUe9O8j
efnGkDz8FUTq+0yHLSe+55lonUjJf7vOFFfhXcCzdKg3+8yGDqBh+3aWyMNPpYoB3OCTt+VENSmk
x0hod64sQFQ9RFhA0Mx15m43EpUwyIzar229CtoXlmd8Kx8/BhLKyaPBJCqBxDnhsLx/nWfVVYja
lDhAa53X3B/S+MR5k0O/5s6t3zzwLiUNBUmAbgvhFWTRdm2qH+AF5sKFWec0d5WoJ/9KEWJCKaW9
6yTcw+sn+DIYfzT6o0b2rKqRVtF69W1LX6hQD+f2yh9kfjUBy13S9C3brVIwy7PNVBxehlZ7HbAx
3fR5QUgpV0//eUBiz51e+vb49wULv63ljTg8DnWVEHpvp6+rZx7+caoemRvMxw7kKoxVrbqt5Lar
TvEiACMYeyiB8Yl+W/1MNi336ji2VlkTc0znZlHvYmBezGoNb/AK0a6/UxXq/+a0KFC9fTG3lM5Y
eW2P77VivpM2pGQqqJr6e1SNxSfP5wE6saeD3ukfDhpR8/BuhUuvplzIdppbhbuIAQj4UL11LflO
moG8AV6F6N/XvwsxlDlipsDf6s+FCsxergCMztlDC9Nehfu62pVo9EBiZN4Iyk0BmKXMQ5vhHM3l
6dmdgYwtJgRTHOV30XTmxYEh6EFeQys2FQ7/NUe0ckPQWxPX+DgX6xlAjWToCH7URbNRcx4tuOcl
NDALOPAMnSh+1vjtM1Grwkpz0aLjrMxqhfDKX2j1oMIECDWAnP9IJHbWymg5+zeH6FABitIpSs4H
/aI/IlGL4ZdVq8AuslzOtWFzZokeh3ocayFd7bWjnqczsAkXhl5YHh5mJ4jyg6Hz5X+LJv3MRYu5
2Q/8Tzapa3hjv9p7+YKcG1lailkI91jcV67F/2sWruYKCNekZasvavE6WuMqIvzmyyb6KL28sTGY
3QTgUhuPT5BjzHE66JYOaJXoOeerOyxvR1cAsYuWZNSH6AjwgVma8hEROrXXrwh1n0kkBbULEh9P
VVQeoR2VBKFPPxjY9T95CpoAZBgxMzyr67P+xkSIA4MZmQvMIKzejVoYtsj6eXDYYhueqnXXQ60r
WCLApufJNm0zE81s0HCIQJpD6yK9l01vp5ChokyP1RYtp8Nh25j9weTYi50G8ZoXmdWGFz4HIaMu
3m3grpM016rG6fsIetCFOS1tCLUBF6UnyT4b/2ZKVYn9sv7VgipHOz6F0BtlKFHlCKrLBMPCMcQN
fBHH8BsoYW38gMgiSt4AXw8dD+qIxHFNSM1arp35vvH+nlyFq1uYLjPWDulnjj2kYOo+kJtn5tv8
lT0KL6eIZyrwc3Wd5/suU/lLTfXhpd8MqZiwaywJgcmvtm0RoSxG7YTr8sy75TIoulwEotgPAKBr
J76VplJ/hhtSMqybZ/cJGzdZjBUGMbfqUf/bnE3VuYo0Zdnmj26zzmzhItZ5ruvky15KYGKEhzgW
cZB4uMMCT6q7ZtzIg9vs+o4A44LcmIipsigT0Qw01qHFhKehCa8rc4z9skTWXCGEoWtBR/CWz17u
9vdo/xU+2ciyJ5e0suuxrOyn0ACWwIMSU5dVAxa/lnFCA+NTwAfbXyvRn0qUYvJLE37Z14YqbcFt
Cmgdm7eCN69IwmGWHsGb6v4eazlX5f+u/d3jSLVcnSAuL4SO2ZuZ5Re8Ol7m4ACiaLIXsy68LNPO
vPRd2uUU5AY5gYjn9ooPAcC0jVuDMmxU5x5fFGuQ34T29KOg9v1CZqEEegCRp2Bm84POGYVH2aLy
wM+evQaFqAeg/w4aikcf/fYdZx7lBOBIzcLCHdZoVBJMUQUzgUVP5mm1ARx0iz7dKlPInvUk/Enc
W+80c5+T++Xnkqi8WZCxEPvG/KT9U9hO3336djzFKRPEXHEIg/tpmAZkXDSfurG5exCeUmeB9VM9
OANn8JGHaDSDOAN+gE/fK9goZIFXDrjMW3YAlHddssn9i+ZMKfO23penJzdQeBj9w+1yvGPCCNrk
NgrzMi7f4ZwOb32prG8T4F8ojkLBfNpi+mO/HkpqW5KvzwF/aXu6gRrIib775W2ie1dHkz10BfgU
0lWCpcC07NxUacfF8yjUmUzxkDXbeZuQ0JdHsIx/0UDyCMHoEEMl9B87tJp18Ri9OzbDCik4T9y6
ghRjtj984uEZ2xeq3gePiZ5aXGXyWQ3gIkcSvM6TQTUqRKLRbrzXGEWKbfK/0AG5WO7MbPvghHso
LTCvGZB+p3rxQQ22s8TkP9Zsb9Cet4pFwZL51sL8kYVPCWj3PK4yToj1gGv9adh3EOxzFcN/VCDf
/orcESN2sqxb3u1Yr/TDL2LkH0cneK/ASSSILBARHCCyLvapwrkmAVnlQvqtfnHfortccjYGJvmG
zIpOBjddyhvfm/uxLGGD6mZ1TOjH+WyQ4X1YIJSairHAcMOV9615V6/d6SIGQfpcPcGXy9BxKZLp
HowLnQW8cgFC0M/B4cDqnbtHoIcV0UK246RInb8Os1+thkU56BVpuV02k9jGd5I5oxvreBQzZ0JJ
+giN0JUcvl+V9I168QanQIw7XfiCs5cKCmnpQZUPLD1XqbSbkluyaHUe/ZBRhkUKLs7WdbU2xPsG
oQ6hk1zjTa7t0i1YEipaHjCpgHC5bUYJ1zhn59DTMek+JGOEgQfPgx97e9UL0Kl1cZPFqK5EM7KP
sr/SuxVvkHYWO0vi3rl3PFZwV9nF7njlVRD6JROsismC2hdhH971843AqBNf/6JMy4Md0qp/1Hgz
YbESSBKEiR3byeT5C+zwhgNkgsQJhwW/mllH12bykSpLD12gbqjUKX1bZhvdD/spT3nEBu3EjGui
ho/FzDt+mabuQOHYxYh+LAab2rv3x8fE0qvsqA6LdIKosyfyq+svjukvx3CGzuwRfuPM2JGVUQVz
GZOtSmqdxGqHGQElGxvCdFJvgb2tESazDiw6W5Rnbm7wq/9fOpZUBzlLGAgdEFAkaqDDURNz3yCG
pnMaUhPeJeh+UWCFYqf24nOpuQI8j2q9mpVpMEAfFxkNZcco3Uci2wi+8CIsBY5QtYG0wffpbA+U
/vhHoGW0lDtidoq0dPuvZH1sJIofSjAuUInFICzwP8P/SbaVvgO93WMlKx8IzsQaKZ6fbQlu7N3J
PM5xbP2wKy/qoDgnsbZ896mk2mHq3H8BUVutckUrQGHtZ9J9woXYE1dvR3vHhf1mc6LzjK/w9SQn
w46uFM2ZNuXaiHeKDvbURuzivARxdUCXTW67lymynJZXGni7+7wcMXysJ6ESF0UAAr7usKRQz4nU
HMQMduKHvc2S/FfGDrzCFhI4MMXLdJOIGfzk+JTkcLg7R0iSNMxmzB4aZFv46RrpOq4aSKSZJ9bU
zXyB9ONONLbGj6VNwD6Oc2hcBGYQi3ezhSMTMLTSa/imKyfXZeNpsybY4j9N43NFLdFbh7f9lSYe
qn8HNBLg+zEPswek9aKVFvOTBOSvP/gaydeLqpuX3sdeGteo/mNOi25rho0Mehti2ExE+cUR4h9z
5mhkmovDewMfDalsu6EGWA0fiXrrR5MIVQsHgnHnM0wpOoCqHIC8/cvy0n4iCzwAkoehakB0IUFI
sA7ty2Um3f3UZ2ntSioTw4kE47UHztReeb30/qWU/9oVSMRF1nJ0qutodnr5x5HfRf/EFGDRqZZC
r1XCv38UxNtvsoxHYn27nCpVyRUvqLSaGqRKbBNWspEaaxsWzfxL3AF3AjRWuzRiooMiqNhqD3i8
AkKtUHtpVRK6uPVGrerdRU32csB+ULcboGYW6yT184YtDtfGtUGRRXeVTTKnPZnl3ddB2PkG7+GA
Ef+N4xGdAskG+5lvO/EWyik2N2qKIlDxHvJSciy/7YcUCNjY+nMgeYLhIeW8aSnHZQRBJ/RqIERP
sJhJ5OkUeniFSTZHNBzWSaIwuE/lVl7adX0c5D/t4i2aOmJ1VXfRW78zXVTnn50T5VbqJ20Ag5qr
0VY+sf8utiWcSCUEGOgZ+9OJXXFOfIlAwrHk53kNGqcXyv6ZIW8N7d5/EydJjiXB2oCVm2i/862A
PbUK1PaH6cS/E+2XMpS+1WCGabcisd35J9IoNNdsrWlE/PmD1OFVZAV/q8ZCrM6s+Xd7bpi8SIZT
HfOZUagezseD5pSCHRBMZp8ovQxLaodaCiOG+nsAEqu/NIj0UkEoEi/CVjRuO6tB7//0k/p2grw+
09esl5IZnZIt9J/KicTIm8mzYO+xS6mG7/+7qtw+D10oPWvFZVDbgL7JxqHvrq7SZn8/meORvU5L
V6B10ULPSdkT6MA8pwH9hF9c21vP3rVtGzemo3o37YIfTIcg7TKMOODzrmYHo6HPZkFZ8mS0nBxs
iZnPjqJfHqNJx9w6mr0tWTjyBKe0bKgfDx82vWVmncbfXymPXY63rT9Ju6p/WVXV2dpAoHgzYigL
8vxssXBDt+8D+jRgA73u63uEP2hgeBoldH74o8wiDm2nR3Z1DRCKGpbT2p8pTPnB4DpgLDl9uovu
TN95XE7IBCgrT7Hd/lacuXO67lBNfTYhKp4J+VMKKHSvcODx0q+PxCUoNYuKgV5nWF0rEdw4Qcq7
usAF7z7rzp6zXUIXAgTvKJeb9VFbCGv4bPPBOGFBNRebVPA4Iayr2PPG7aGGDu8QH5i9I+enOdfF
Kq1oAzmOFaSlrUKdzG2yTX72bu5x8HkzDLpZS5Wmldte81xFhwfFptStiHh/UUZuIoTc9sLc8dDE
zsev3inu0Hvd+ZyoZFKECP38qvQ4qOs0sdxmfGc8D2ydWIV1p7Q/ykGYQcYp3912OQ0K4rFtHcxx
rC0muJW4Q+FKo42DJ+SiDaWmuh1O/ACWJmZR/jVf3tCzFZaHgFiIB1Y10p5tBMG0FoxQaoEhc4Kd
jdJK2+woHdth+UweQUV9n+fHQPmZe9CzObQ6TkTqdu4iUQTpAs5xjrVp1HIP+VZxQ2bT6mlDYQMP
v40BhAgQTWwXFlMksRFOCezTmWhAIP+24ttFABMJuSoUgTHoL8zzDlj7VzycxwyyN/HE6914gFfT
l158iG1MCEzsTFncQux9tHl/3sLYhpY3FAeFLMpUqsWkaUK9O0idgpI2v9z5nEuKoMkjUoh5C8GD
yxmI7i+4mNHPsrMyerD+ASxnN0d2x2w/R42gT3aHRaJX4BxF9uP1IFtp+dMLiaBGdxNuBqLRgL74
NrYmJwuol/K+1dVQWt4otDGuBn6ClCQvVqCPX037JmOVgS3AdhN2lgQsS0aInR6qckjBwkVUIbQn
c3wurCEQCF/K6E9bxjKppH0yEVzYuxKF+qhlIQ7td4MATPC/A/eK2Gi/dg88Uidvogj+JvdLvJHf
D2/bi0jkCsHdFpXheROBY4YdnjvXybVA2x+Xa7cI6tEaRuwQ4DhI/0KRjhSMp3VfjiHF6gkF6Yx6
7harCoHxeLdh4M76tVg1SG9aJk6U+RKETICT3c3uO+GTtLaXtxs+UQk5XHdZuHvbs1eu02IBm7c5
suI9V+DFH9XhaD/KV88kL/SNfBIkJTlpDtPZuwuT0r0glEX0+PxfxmB2ECC64yOBvRkwf9riz7fs
dwIcalDVQco98a2K7p6Yz1LeVflBFi3dZFX8XFCcdmqZwohkvUped0JmfcVQI3GxgVXC8UcqPJki
hBFEP72DL8ZsZ9r2HUcrVddkYLzXRlXA4rVi4CSxFw4a/PYmrGhVND6GhxFYWIKTRxJVTCh8+z8U
WqObMwf8gaIfGqcXn3Qr0Zhm7ctp9pyxrtUkxQalcGz25VtgnPhgQ2mQzMkHBA8vPoLNQY8y4PhA
HNtif8payRuQdFO0hIg+iAFXnJifzu4rfQsuAl0SuLS8EEf/xZNDqVf249MiN16thDGITIxtCNEd
EZYWj/Gz2ddHGfqyCrZzmgTH7pcjzvo9lVB8cGes3NUjlnNB55Q3yVjHqLTsE8So0VoN+AcDo/fh
53lYbm+KiLLNl6DXKqNbVi+XOs8f8dvt5K53oOvhBoq6WG/t2E6v6/0kAFS2rDcSnCd4ffG9OrUk
2DxlgjFFWFPDdMoFZtPRTuTdYHgchNAYjtT6AnSUcnetprfn3xaDLUZ5yQAe9/P2CsGdd+bglVk6
Nl0g4nCZ2tWyDhxpLNc5c/rRN+LV3sqQhvOLwk1sjsDYqDAS+QEh/Cj1AdnwJ6OAAraR7SC3p/RQ
6er+gh+YkLahi0aY/tnjAn0zJ3xRmWLIkknyj8YAqGEv9gwJlVVF0YlKVxjUu+XhkGLybfp38kAa
HfH8T3WV7Gmb7yvkpIoV+YjaezD4MnAnIQUe6rV/+A2agFKh1mOClkyroQD+hthlI31mPr+z395O
Su+cNn2gs2M1JnOlwioqA54ta9KMA4VnbTEF9RkV8E1VgohmCdl6QZQdAbE4utdTjhRUFKCi63La
mOu4QAkjv2QHt33moJk+73bUwyTV+cL9JT8F3NrJ1BUGJI8QAbzawPTuLRPkvBXsddryV7QrJFuF
EZiVkLqhmH6BwYwxPrsJc9k5oNUGdhzBz5f/RKPcbgDft3lnxOX5YADF1wjS5PMR/m+K/NJCvK7W
25sEdJ0ZK7LLdwsPoBmNdZ/5AIPt9D8LjeQhY7CJ6j+nqyg7Uvw2yB00IpVzysD6z1lNsS2o3x2a
Ptg9uU/4SsT0KSqQpajuNp1wSV4bjJaBgu+xvSl22PRDOc8Vr1RpfuCkeu9u/cNZAHV+tESebKBd
YNhicn07Fq1A2EZOHycAHy53OiSJzoMALUQugBm7fQAFWCoahsPtjLb87mmvRJ1MSv1UOJBgX2mT
TfOka4U3KqdpxLkeJC7vhZpa+E647PqtXu/CA8U341m+vbYfFkgR4eW3YafZXkL64YWZt0pFLQp9
S5JpmhtI8bSFINqCbizOe0uikh2EaPEwkyiMquNnLcNuUDjSygQxHyP4g7Gm1iYdx0I2qUHL7pDl
BLau70qm+1fxgpR36aqXjhx48XKceYPrq4aZtoXZG07h7n++ZOIMVUNylCEklc/IZ0+cqs6/P2P2
/7XwH9o1ZAuEwLN82WDQEt+rtqCtZFWi8SaqkCSFR0BT/rexssalbSwudJpfZ2lsRIqpBniZht0e
E9Rn+xbHjBccbVo0VCUjyeHsulGxKUjARmRUPG61jBnpveIuftRkCzdJjWpUtxV143NOXOf/BAVk
AX19YgOtmbhHRMhGdRpuL3AjOGFEBfr5kYo61o1/3OVazdFLZvfVUrWQp6hN2bWFsgUuzw4D8TTy
t4kAW/FaisbL+JtfiSN+dL6lB/+XXSYhUJjkvudlAo9t6UrLE5Gftdf7tE6T7oazUJEdwQHcjlCa
9/gwuR5R74XvizwBBYEej7Z0AAq9fcwVzUoTeZtnB+WXa1sLZ0rE6w7lItN9amw9AIiK58VYK1V1
qRa+yGbfKwAwIvMKYzjxu7kD6GtOB2sDJsKel2ujpfTojgN8z/miLfyN/ssvdE2s+nFpTXySDBsG
nQ/bX+Nj+7B9wEbj67kIXwBJ2CHT2VNB9OnZSNt0EeJHf8QidvvE5JFds3s2Mpos6eKEPzX8cUv/
tZYEG23cZrYjKr1Endx+aLll0sM6TOdkNYTe7zXabWOYw7QuIsOvWpcesj8tI+BmRkquH1+Km+dT
pZt+BJxOuYCYIdn99FbY+/wI87rHVIEPYhTHsSTrNRlBh4cgRRP4WA9nK8jcipF4FusfiLTJq/n8
Xk0izpROXG7eLJ593sUR8AJmkU1q5Y4PXVSzBcA+9skwWAqpZNU4fiLQzJ3TF8QZLFe8kueKF5/s
rp0Z2unJn+s3w8a9khfPpqAnVgXJktigVgl+FeATR6HTimIQdDKSFotZlC3zcRRY+lX3h/AljdDk
kuT5YJmqTtCOJysS/8d1B3y8WoSnFZynejiCyhfGa7xhYhlnwjOp0cMKKbhqWiS8uyXFh9BBjbGQ
UkjgDyx/lYNRRn8rJBtVuBia8tgVc5rhNq0xVLTp1cmXswyPQ5Z4SBvhmwZHscjq73Eems9F22mA
QbwbddiFt+AI9cYR0xHBGIj6TXQmZ9BsnK5VDz2sf6Nn6ZVZypnFaXwsq+EShM8qME8CWw3da8De
9V3EqtJLHJFP9leQ0OXabZt+cd+CEF8u5dCqLL4TeCI8E5P70FDzWR5OtDRbjnB3loxcyS4ZDo6m
UE5bOHdNAjPW1fR6TxA1ZUWjYSDLkSRaPFkMIic1v8jAhzPwZqqy0Hzw8ylH1Dez6mba08YBQ5c/
KHcMP8NL9FgvDgpSGSxezS3gMdK4hqpNFdsOe605pN+OgMv3hcjRDaPduBbsGOo50qgX92ElX2zy
mRiTOkLIM1lHKhO7QMXoNpY3+PTXLgmTIk+qBTW5k5TgAsa0GtbvcciYu78bIG+IYv0KDhWPgUMX
qUMLl96a23HsEz/2q9hnD/vV33eHaiG77+qpYE19l6srdPyXDhPI30PTbzsRVsaYN8WdVmUNV5R7
TAV83sb60yqukJxabS/equAPUbxSoPvljkWpZXH7pQhy7jlJRewrxWn/tOxbVvsApi4x/t6peNYv
YsDpTG23VxIhjUdnXm0MO+kYYVj/eWa/tptzZCXhlhdJQW5zEq5/LcWkoxE1ZGwAVgdhxNP550u7
qTt5AA+h9LmI+ISB25oHDME5rL6K8pQzycILpM9z9qh2UNQlA44e+4zj9zd0COYN17qIxGYglQ5O
oPdIl4+E9khlTARN0sJiloCMwBF0OAZrYTF3FVIGeJAjPxgmPRrVy70Fw+MWz5yOsOblcEsdk024
+UvBB6fM24QmxHbwaSEt2QKwnm0DJPiVCXtZ/cSf2VBoD5n7ttOEb68ighBw4DIQ1h3+oAFHppEy
DVYfTsnhkmrlPRJRbs8dAK8sSnEYYKWBCMR+LvR2DKcBG4vsFW7F1PKxdCUks/wP0vphafpCSqWh
AKm98nLD+2tNk952FtstLInkJw5P4QyCJgtyLJZeIBYMw02v3jnBjPF4viI0yP+cHSrFySYaG1lB
FXX1156biIa5+yzqouKJmSQObAUCVHoMsktwdvPfEiNz9PMRrQotlbksDC+TPnj9m9hBD4HXxDi2
Ruxet6AbcWiZg/YqLwSQUOCej9NPUREjwawsNFWNA08J01YlSSPcncLdfECu7b/EyvO46/UIs5/C
m5ecUlZbtY0DomFywXb12D3jKZFgGIHUwKkfhB7jDpov2RvTmuQpAfGg7O6+AW2z5IUgAHAVSzkZ
q3VWJkF9TYQ3tRM2M3Utj6nw0LdRZDhU13ObmrY5dteUN/mqE/gFZqCRTkr4nIrlILhRjTTpCC00
27wJtghqrMDyMBx62uo9nMRoyfDPbr67zSXIl6KGo/MUG1u5pWhSWb7XoscnfWw8qlwyGMOAQrXo
wtl3Akj66c57EPxs43J3p8K0FEDgG4xbeQ40yyRkX1uEiORZ2RMLJf/L/wfbhXcozwqzo2QiftpB
Y/PalMe/0g8OIeG63q1nbgaS4DEkPcw1wqcFHK1jwAo48qFmDDFWATHROWzBsfZ7HV537pxalw/p
hguQ4mWw+XL+Dd/B9aJn2/cR3eOksZy1OCQZSIklmYG0LNXvMkhsHObitYBJim6FKgv8kJZjzzPo
MGBICYF0Z60yKFAI5R6+1Y+5Guiv42lJkdyCoeB2Wqx4bjvfipXHnbt9O9zAF/x5Etv1Y7/NLDwK
/5SsR7zmdHdx6YqkIMPTvS2bxgs3ofMsFDmF9fSm4/jtBr9ArOAg2q9X+UZPhSr9Hh1db3n1wlXJ
b6aVwW7P3WWYRaJ+1x4LHbA9nTs/kdnh4rx+ySHNCNULsS5YpSAeQmZK6aoITa4hBd+WMqYGp3ET
9kiSKH9qyLtHH50cwF18KegXfd1d7+4cZ7syl+ZuR8/4oxq4uSAvF7iY4yU3+3xBeTNN/gRMm72B
gQA1B8B8DK5CZyR9N7PDcVhBnTSqA8FaODsAJL6FvYDLknCaZVC3NFlPfAdMfhLFA290seao4xOF
bg0krHvdTzIeIkmeN3f2l6kQgbweY3wmHKdcq4STE3rtS5zuMfnyqeL/5PHaO4ttR/PwuOElFoUB
G6pds2J45/0gasyPnJQ40bvSpb/+wgqw8+/AcXWP/b6HI+5GwdgZtyXkeesCArf0tPoyZkAuMRWo
1sKwi7VSRAqt/FdsUrbT94igIeLX791bN3KyUnLjFR4Hmz/amYlu8VjyTKXyNk7lgbim1y/W8mWE
YngPD0gIwgZgH7H5Uy2yRWmGyr7Q+e8kHIWpUs3MAGhekzjy1qHZvQ+x4c7VJEdLXtritNerSCnt
XNEL62AgClgseuLzCHwPxpBOb0yA+7rXvhMebeMhT9OXIpcKzMMivsuHfE/+9PmqBaLNGWJ9pcbc
1ee9bze96evnUu3lPqYF//BRWubPQBiK7QL8rUyBGu+yvTni8QQdqAdgX3lPt6zJy6Qor1t4XS4o
DhYwa9egc4eRSMEJ3yf12+loH1TDzWTLT66VXlb7dK9UIjAb3bAu4h82eyjDPjUMCnqZURyJoI3c
gPbQbNwxoByU6vxAaz/BtG2soDaR9bnPpV/DIsHy34DyBdzKwTAObg+Tiy+19vLnc9OHFxdyTxm5
uOV28/JfbjtYUuDV4G84JzergKoLfhlDseP2eqDhSj361sEuInz5FEjvkfbqglXF6ejL/q3KhjQ5
lE/D5b7njFY8/evEZFrLGbWoa2H7ood5mkwK4Dnua+zWw8vKVv6XEDMzR0veKjk2Fw/UKpLqVxq/
nZcTqLwUnlnctGVRZ75YSXpJKDnxXnY1Y+NHc2GXy+lY9bC8hGA7M3A1pz5liMQX6mGvi9g7tHZz
v3fWDlcCVF8mykC+/25fu0CSMy+we2LSWxySaHHP0J6i2QqAehPleKyQJhw6LSD+8NPoSwSBGQSJ
UrM0dknXqJDsqXehV+DhhpSB3IOKuM74L/k+S7Yx/ZfjLHL1wbZOsnGRrswBj0IzceCBkVZJC8qv
RU7bkNd9oa/uWV95N4NJ3BUutLeQ3EcvXyesjdM0KVszJwPr1nl8Es98kxAlqxnhn/I98tkg0ZxJ
Xo1xB6PEM1qCje3yjwzBD1k3f1ArH07GO5o0tITl8rBfDf5V1Tr5A+62TKcswkBeuBCTFm01ifMM
6aUlb1tkZCRw7N6hX3FncGtzfsen5YpKANF/UO9K/vfSqwIjLiH463cTxMqw1B8gWMMZwOm3uwrO
AKlLGsW9QE3eUVzuLESVxAhKHhp+ChFS7N0behLBqpohzAwQ1yoQ7JX6b2tnWlTPoTcXGPirbqMC
o2BGpaS1yssqg47vqPB14hQHRVzd9v46U0+CiNjJPe+XgQu3C0l3ayDrWONjM1euo76OUJDoDjr0
YSsi1xesi2A8Av0hR6Z7jkAsFq0TCotQEsIYSxV2cHXiVW/qcmX6VkTjQaduNdDC9x9zAI2R4xjB
jycXPv+V+z59+ohE4S0hOfVNe6Tk3K5S+oEjkeUXFDhNnVVz1lx3tu2/6V+k7vCFZX86zmT3VH5Y
diEUR6Fv5Ys5KQVYoCBHEVt22gPLSJncfFupJQJkxRPlX1gKvkr4kFc0YDY3BEVqdvKnlzWNKgqj
1nMH4orGS1462mteWyMQ5nD6342OxcQvGQ9xqbgAl34K6Bm842djv6tDxxjfCViniyYk+EsU3SWw
70dngV8giYJhaskrwcr72qnHnIUZZrX0LFbyRCUqti9Kj6ll671TykqvbotL/7mmZLwaf1KYlxF7
CWCxz9ZFRm7PODAROc7+84pyoFEVrxeePThDNLirEo5qkHLr5ME/jJQ8IpNUzALmRBqfyfUzgW2m
F2G7F4q7zwvmiF5pyMm93vJdFL52qMOMCJ7Djt2AWEwNxK+Xf4h1Mnh7AHrqjkVZkKLSo6SI6pPb
Ti6d6h8/XfqvrllFPrSDo65Fs+l0h7C9q7I6xqetiX6kjjfZfh2a34gFg+NcI/gx3g17yXcTQUcv
HTp1kHU1ydiOT1fXPhOo04AnyIWf5eYlqSvLj/72skC0dFwEaFCbBvMRgfQ5i5SWE+vS1Y87XsRr
2GZMcqvye+I2T5YpGVgcAdfdAsVDuSgBsoGp6OTLLepsd4P1hCx3nOfeDnm/G9z3dn3FczwP9xev
HiRCj9bweH454I04Z812ooqJpOYOIPUW5lv/AV3rLOD3adGnPX9pKJygnturMfIpEiKI4iAOsNUS
lPfECsvEjnmMIaIE4yjIKznd2wTsafc0Q3UfA9ECLQHCPS53S9V0/IneZ6lUCj7Dm/US0xJPpOci
syW7N1wZCYBmjNoSRybDL5HdY63H6GyvEaEjqLR/mfF0zD52tzSYa7DgPXP5KOKCQavHczQQvKL9
Xh0EN6Ge36P04YzzsyjouzlOh+8NrhiisxAbCJMJFhWTU1cb/Tm8vGtjsV1OAVQxTOGi3DFNt7TA
k5e0CnfEZkryix1DA0evuyZIsolb0pgQ7GX8cHWHhbTwcllfTmfBBROumKjzHwFC9/Zius6wiIv2
lUg6fYFFtgQpbQSFOl93PJf8lSbMjAgTjxL//AIO1KrD+XGU3LfJhnrDcNXAurLdAhOz8zdhvx4C
7s284h7R7C4tgA9gpP9fMHBPDPim039gQxT/gR4s77MsrMpMiG9QKEE4a5RQLQzkJfwB9GPfRY/C
Wn2zDR332bKPwZpDmkGPMTUkT8bGYFxo7n7Wp+fooatTgb60vhOX3qlC1YKS1JIU42lkCX00FZv1
EhMXzEG7qaGH7lxdwX68cxPnsSjSRQ2aJhrGhgGNoK5qA7iAXZd3HoDL/qMdmUjPuu1Xc+sdc4CC
Hpbx9jPuBzKsub35CjhMIXASi1vSLnLqVpL/nU+4mzJdJE2X8Ra156DJCj/fmgxgfA1GLTal2NiZ
rOBInIuTWo12utlE+P7rnmXl6v/NSTja0oL2fJJl8gnt+gGQ/aUSdaxKCHdA2r46EUGjrlTDs2et
xkaCGu1nYxfvDyZdh1m9sn8PP8n4efY4G2r6FtvmgLbgR6T9ojGcIIACL7cAXs07CeLhm3Rog9/N
/emyBvTZpGAZLx89ZSGZtZbvSG0LvrCyd8X+tG8UwqKPWPZ2BsThigP4maZFnyJdre7B6T+5vWCn
+eXuHuJjaEuBFNWHayF1/9xS1fYYfbv/0fqbZMf6AaT7wCiku/uxNzSwXReMouh2dbLxXUIsfRET
3wdJHiJomhSgIAlh4ZNFJag18zYAHQ7OtTXORb0rH2erGOrJ4Ca6JQ6kRWmCkQqzBxZ/0pQ5BEzY
MSTrRtpUILNxHdkrhQmYYhBP4O3OnRgXJe91wVMbwRdWgAUe0t2EuvQ4bOoFRm1ojZCodeBx1gLk
9krra79WsfiqBPFSI1KO9BAMxUdf0QMPz+0xpe3t3YXG+47cwzMDZbDtHtoy4jSQE2nsi0Gkeijq
VTz/LtF8CZhP9sU+SsDkPYGGQKvw5r5JxHahcKUCfITmipwqav86kgqGhH9d0iqKr05g/X8SLhGq
QLWRfxzbOWmiGu6JKbO354QAGiJivYDjWzWCoxF04xzcNPCjRwJKhviRfDdxEy4YY3YJtI7dF33N
xF5Z/n/PMGbuwtWD3llQyV7gv4v6lpyDeF8v/DmcWt6Q5Ksi55i4pSR1ZS+Z6vWT4u9qOSi4nak3
LrJtnNoVtZYJ6MdJO6NxDzHKAnC+nbt1sUNrHlbCTBe5QYwFRDboonVhou7O0Oi9aGTY1WZXETaU
hTHubqOE5+czoiY9WlKvmIBOiQkfHzebh+kh54iRjZOS0z+sdr//MtZIAfARAfa0KkUenm0YfaVH
2gbg1J5rsDlPNvvTS6RBP9vtF95Wwn6VyVbZY5W1FtIdYgGvDB4e+Sc0183sydAqJ1QD5je624D+
6Q87VTth9O7/DE81AQmpHXcMDApziOjoJZ+w1zKFiGDOxzRHHlPe3GPQmm7VwakIoMJ+z+xkueIh
DGJxL2pJRPDxIyFQ2+fFP00d8omy3nfu9TYB6DW0h/R+VrsrU9Xfq+4qLopB6j7YWjBfLAELsvUq
0IqfF8cOwTAHZKknSfy6G3rqvs9uKXP5uiK6F2KmudRiP7jMVn+6SztFAMe6FMc7Dwd5ftvUkHxY
PCtA1PEgiB+VFyTa0k7Sq7jspc8vsz8QgNRrGDIxQjyClEoxqZMG7Wz97jcO/ex7pAHWb0LzbP56
j66RCaOQFoKJQLmCIm6ZbKkDQhJ1EQib0fGfqPq4VQ6zP7dg3iaPcT1n54HTadyh8Wrqw3e3vEXv
K8uk8xA0qR7Yotd1t5TmkMn4FZ1F0paHsA4HUSQy5KNjHovLzZUPWNW1GnX9nA/0FAvxdH17YfKt
r28UmBrkXfE0cIGkCATlP0aGzXIOBciYt1cWxB7HOqLmgzbcYpkCJrpH6goVpTelZ+IYFCfaGdhT
NhAmH6tfU+jktXGshtMoSTHaG+Xe4EKTTHtbiY5oXu9D1M0u6BG/fLF5lJULGT02nuERk1exp9uD
jhQVs3CkosOXFysOqblQ+dDBcsesG0Wiud4zCYN8oNETVtmfrqeh4jboIPxiulV2kStItQh+pILE
jEpYr5KXWVj4TqCDYCNK8GpTHtHgGQcP+kobRjihuVPO4my76hU8RCGTSwQWACsn5MUNLujdtwD3
DvcBEsaiixg+hSdqcnPkuNmNcwy6N9OAzFk4K9NgIK+0DtHy2aBUVmorBt9ImHLLA4Mtp/0JTlRd
jREWqSvRskxl0zjgD6+SlI/gwNHOQ/cgiJT655m8yjTXWqWOfXCMY5ywBHGy/80uClXlFq54b8zV
aX7/3nonJnsqt680i2F7caUnWU19kZ763PyJfty1q2JuT7zNCyimfzJC0cq3Mb24POp6POrELZmI
5EqQxWpRZOhOKV5etqjS/c5fxyRcdtR++DbfKJ39mhKnbdxdhfFS/oUBU9ELBISHT8Ay+PVAw7Vs
xloHiEK2p+l60R8NsuxofpFzGysZWdEsfI4ZUS7IwgMZJaMWsQek2Wb2PAUW9iP4Zf7D+DKGs+Lp
u0XG6L2ZrUYm9rqKgn3n9tWf9VSpvgonKKgAxzBhpp96Jg92P+hWMs6WfSsYDnnq1irquEjMO0Em
yHXGHKLxpKmISX0ScQrDf5Z9FI/RGuxp8M3bz6TS1lPlQ0uWYl1BBRlUM1l89sCKzA1CDoTOd4Dd
mHvPzmnsG3KD04klzJBsUb6rIyDLPJo3qPHX9HEOQWkwRfhvYHwO7Zt+N7798ahTcUz4mvSoRD09
8PnKws5KxdNPksVXcVKBD1FcYvqkFCKcvsunzeMx2bBGsV+IW0wW4MAL2qeph9R9NcFUzs0qfxY0
eXZcheNBVlrjRyq5Nt4FH3RPvnZHX4IDXTWehLci0tmANwaTt4KYbdmGLgJLcS9Km4xH54aqQ2e1
9XtPXMpdw3yIj27TJLLgc9nYTKOQ1zKX/iVlGXLX+TYDuZP3s6HrkOLOBru63xDAmC9JU1qfIpxv
GnpqxdwclEtkFUxaCTphv0IZBAZf4i46vqcCuknqmszva4VinFep2ouv91jFq07+oPjbbYki/ott
IAVL9MCB02jbJHTLiKGAkQAJh0JHO81buRXt0Unjss1HmapQ8cy1TjxpWJsHO6uAeUxH8xwO8aA9
IT0bkAUQD9gX6pKbk/kJqSF/NRL4xMSAn95W0iFQCT9nvdmIG27SH6BU91up+F7xOTCO0TSms1Ei
lldhmCLLtQ1xwLeu7rhLvuaGYgp5XkYnF6+TnDCGwYYDsqsfL9KI/V2X8Q+FtlIgDVG1/UkAaowN
ZA7QH0MdHUwO6l+NJwx3vu++SSOmDHmyHSYEWKTGov8YL/MoaAaxAUAsTwanJ3nrCagJxoVBXLYs
Gt1G6MqnUxD9SBeBEveF83EOUpcrHyr7vVJDosZOb+aarfI5+M4X7vg3TO3Ucsy/0YB67NwztQe2
S1rUZX+s6GcChadnPo1zBDNInrVNOdpcJi2XneANUxT0H2Pui2Wejd3mg+l62rAVPPTY615sZsJV
99Z2O9h0qmBBCEY0pwb4MRNoaiC5xZV5r0ADxHQOGirYFKYYpB9OfNazuIkAakb29+E7LhGbGtvC
mXZDI4+KCuFLxxB2aK8fcXLJJfDdrE6qltCW72zmLMAUR3mfAV/MfGJ9Sp23Isic0W8+1mA7O92B
p1Mq0hQiOMc8e8aLOo26xQzi7mZt1ZtDdgPm8kwnkeflrNlJK8MVwEy+sdh2PD3zgIjtkRc4ZJBN
3JuqFw4NBd0uT4VEK1nJKlRXKojfA+ZHOFvdR6DynddpLaPJ9pjEsjNe34TV+SR2ME5xFJXhW4Ct
pwk7Yde4wK7zAluPQEThaPmb+3nkUu7bWAxnlTBEQeBFTSJYguoQpklHEZlpWWB8c6u0CAt+I6p2
KKGkxIjJ2PlhgkpfWshfrE1wakrUwa+KXQhtbjv7M0zHlSg42b4ChNrSMpy2h7R79PUFVKLbWEky
E+4U6U51QT5CsxwaI0QCbedh8ZAdOp5Q8A9WW1aEMjVlOxVcMEyR5+wH/LxDXZrdnytb4E0or/iC
51Ls9ZoptGm476Ynu7hQv362BpmrdmkoIk05/qPxkRBuBOGXBYhkQvAtreeVVYee8jxFCkUB67/p
+e2Oy5XJSbf/9HHE2lsJylBePhThD7mfQP+tjoRS394u0T5a3HZKuIvwgUdO8ppOWmpGMsotlC9O
rP12IN5nNzVOXs+kg90PYtKwnD5F75RRr8uu0Fc0B4lwY+brYvWr6NGc3RshuLxgsN3clBw0oxC+
fNdMWk3eRKh9GyO9in0ag17o2lF7Uq72lEvyLbsHZMllmIrmFgLM0z3igF7RB1QhwQQ/Os7qZHX7
+Ez3VQXP0rRiGVCq7Jkxpocf0qxrMnfj1FTSXMstSwOcLbi7lnSbws/aGu76AEdtKfmw9nsnsakB
dfm/gbQqPdIyVzDjrUZxuGgp1QgX6Tcjl3zkGY16ENlieKpBUQB1EOEpAMtgEqXUKUV94+nSRil3
Oxw26TEmIbrYRyNVWAufGw1DhlPG2EOIL59AQ45aRTxqi6g8n1s0fgc/r8r81o3JjhvoqrBtI9Mt
p8n9GBp3No+9qBi5oVYcqo0SXjJECPKqM4+Ngt9PNLbNG5yL5u5Z2qoML194+/T3/7n08I+vc0J/
xu3lZVZUhudeQk8sr4Vf0BeQMjFTeDXW9aioYkmnzydieu6ei6Dyf7gwdOLi5Y2ensrhriky0T/9
68S+Kzkh4IeS/5qNWsuUu9iJeIk3CLzOYCnwOHT/dZgltZe2lV33bSO7a29Rtx/KCXe1svg0/Efh
IB/CZysMS3HL0fNDyTz5aNUxPPrCe0JkUIU1GJqsq3GvXkZafWnAATKIs0mOGvHZF6gyh5cACGNM
i3btbq7W68O/ygdoPiTPU//4OdqknBcCYkQvtNqsDuviPLFj6nj6EGMG3OdcTl7Ct4H1feNxVGYw
WXq6bqGHX2I1yzB3B2unmKYE+3CMs+/HdL9ni+eH28HwLKjOHIgmpyLkyLMP/rqlZRIlfIGBM/ww
zeF8UblRPnzG59+n07fx4wvegCiVXcCC6g/6AHdImHEVNTEacVNMp87/8IRd5K+nhv2GGiiqhhnl
cNm4KqYmFBeZoNHtrfsQXqod4Lvquu4SKEVfYhRJ+1x3Pnc5OtPGuJCb+yBhOLSnkOU7iIuuqvnm
/2DxuqFHlFI0JQNyukHDRckgj4MVRVaur1MEIM3eo3k0CwTN7aC0gqyMTJ+iCZXXKAz6gj8AR1kP
diVkv7zV2syt2hnxZQB+M0zJDa3SPnvdF0vBkNJ/7rrKK4nm8v4SsrivGsXeuMtihGJq7X4hrFDA
J7ezWkL5IjE1quJQJRaqYOIInrMCKMF19LoX7/hLnqThOiefDUwBdkMscE1oyJScjRcpyp314fPG
6XbLj9ExliUw2O9TzcYTnrS2n7rgnOGDUlYybRgWhB5ngILfHQVuOVBdbYBY6Km//3+El7PVyYIp
2bH65b0FhGBu/J7AC2MqwT49vImspDYmCqUD96xgtPuP20yijEY0IkOPXc2RlMWA27pmNvX85Hfc
RiTJ7fWfRpHt41HSWBBHO0jICH/ULg5AFixzdwUt23C/M5GJONf6hMHeUjt7sAgVkeea0Ld4sD/k
yLUOUbBmmGbLfmV5rrrn5HtedjLhl0+We4iX5x0ad6fHxAshZcD314ReUvmRviM2w2+Y1/SGCO1C
cd/63T4dGGh6H4Lo8b9Wbup+sCc7Davl6xd+QbFUodKJaexXLX8jKfbwuZoY1tkIev7g6ql7xLrv
Dfc2m7yMSm7NuhXVeAiddEidwN9OTBC0/l6FP/69sG/oXydoW1iXhtUbuFjER+cttUN0Q/Ais7uC
+lY3/Pi9TSJlPds3jSjta0aIPaXnShS/sp4+14UqwHnP/fCiracpmxBeLR3bMwalhSiwdic5luiL
t+PfWuE6cZ/xh4DVqeMIm2cp0MK54D5YkOy8Dm2HQTzRXR/FmxpEkBObsaUJivCxhxnhlzed2/nb
i89UgTT/mCDgjQPYg7i8JtmBlmwOCg099P9LTACIOvKtQCwSVytGN+qGR+HeeGNlhwZXT3NaqG+i
DvTVo4ulVzmIP81fVUrkIj+4O/Gax+CAr/ENThvmboQwxwbNKnQ9QvVBj485REms4D1pADIBdbQw
tRZjyyHIPfVdUChvC9UCKk1VXgwVaJouc+zQJiXXFuHCYT0NNVMffmn/SPmAuWHeWW8W2MHq0I98
9o6AwM295rsLb0VjOKn6zMwLWlmEt0M6WCoQfWx3O/pZmwz72Dw84WV85qSG/XnoPe5ZpJgvR34E
2HTpDRcJuGLCiXS+FY5HcEvqEi3jKgZfJKSiVgBrPedSP5QbKa1hcrszD8Rakq+2/NEyRLpl7KVF
l8R7R2IAAKMX4eso8mZ1S7/iJdmS5ZhDuwkoJoVi8rfGugHJmM4gZB8t868+Op8bHsrsGKYr6Rgg
8Mljrn59q394lbh2vSvBnc4RNbYCD8M8Ku6sLMiI2+oIvTwC+9HYJjgYLExOM2Xy9pa875+T931x
+fkvv7XA26p12NLZuuAl3MJ/ZeWrk86BpIbL3Awcq+Js9LZhaEVPRSY9wyFTkUAM7NBq6lOOHloZ
uXdtjyINR2PpaGSDBgC2kefsgBkh0PjEWJ4MAztepuEBsJ1uWgwZhO52novpgmXSw8Cb+vUfQ1vd
uLAPYee6d75XdYqQptx8R0tznNxkY65QFNptWJadaHgMhE3RKEQVV9mZl6I82hjUopeKDU+gJuc7
GNLKcKypm+/Q7VUN6cd2xGQmD5ILDX3kddI//MmTkXEoe7MKbF3r7msP4u6sYZ6VRyPufb5QTGmT
VlIcg7JRE10F1FLhexfxoYZQgiKXGkDW/rFxpF5UvjpnbIQNbNYlxxG7W4MDeSAZIv3jyPF7F2ve
dwqbEi/qdvdbnSpjroHhQfrnXOJqPcsX/bfXCn9P8kdvsDeO7z6FPjns3SmAxasPKgHJvO0wlfsD
g0kjPWa2pd/MvUGCLKiJVjnMEL6lWy9zR+9NIOyhNI7m7rumwPnIRyHjhaxVWvyJCZdKPE1IQ8eU
7fvdpzak5+RnshyhgmyMZIzp3uAAZgQO1/qD80fj9vK7n4HAzBCCRPCnT7uEsY0eyiQdpA/LAGQZ
xPYihdTeHyUK63bRnho741hLXeTbMBTZE1og0EMQxvICDdOBwP9L0AvDPutbTPIqefdbsQVsM7uq
ZPGqzA1YJ3USP3nVKEE6byPOyBxcIbjC8sNmD91Pn0dGjqV/+4Rkl1INl8VWT4bBZgto9H+mkC3q
7cFc0MauIT1KkCrxQaMSeWoC+PXzqOCYOKz7+zY+DMtlU9txfgpZzC9hQEAmJtsBxf3bbwOrjeqM
KAjHZ9n0IFIEOvznsM+dycJgxo803Lq2dQ8d9hRknwOkv+edQ5eW4AFfTppI4PwD4JMIdvPseSla
TonZvaHkX54kgDK/TEKsBn1/Stn70u9TFzdCdtuIBqh26mhirfWv6ugVuaFXMWWUNkIJP7EV6cTm
JMs+GvyRWURznT+I9LowjRuUMCyoTc91hWw8kMM5nPLwjLHK6u+QKlKintt/VlpZlSaQJDuR+JRK
tVrKbkMWuc9ZMMPaX2vrE2V/Y24DveT2EYA3ni6AUeA/QTnSBySr+Wz1CQV1LhLGlwg/2TBAQSa0
xH6UXbIXs3kpCpf56uDEgSjwlm/B/GVU6f/ZSPUMkD2FQwu3lfo7vQCcjlmr8OsbPHv2Wc/s/xnP
Fld6MzhoRL+lf0LcWIg8/EqNmshgPypuWettnHOKKY45R6VlWIYJ5untXg0BZxCEe5HEGXOu4OqN
zPGuLZQm+THDYe8GUjUvJft51TD8Oh6v2vYisPSwAImFY96R3JNzZ18VXPo8rqOga1IRiWIJzWrV
JTXURayY0L6qX5WuFWLAmD8p88pF0gozp2gu9uEMStm9TRPgoNVhlIgPcdudRLk2S1rWtikAXSig
ZkH65tF5Bl3ACb68uNj6EZ0r/YhtexXvk/ipf74ab0RjBfwDkheBkvMYHXgWtf9LVWpcdNaMwhnR
WBML+O1MZgUu0vQyzC5NcSFhOa3QPTiUoOISZ4PYdkVZ/flrtUW1CLzMxuvP5LlTcua3SqUr7DQp
/SPZayYMjoJoYCLbQTvqcvjw3wnEtde/4SdDOwek7bHlpBs+ZHuf1FEB9rEvS2BsDGqhhIqVlTxc
1dktltH+OXe5PQA8UrOFx4l3+ck1SJVVx7/3/RmCO6I256LKZgBLZtfalBvEOumGXtOSl0TNy/J2
rgP/185JEjhVDck/xaaN/L631fTIY1zibGIFIB7IYK5Fdhzq2t/zWG31n4SSewbrv7rDMJ7+sFUL
w3yM9M9yI+T2K1ZkqPqph1CSrFr/QDsvhcg6v2MvymP06qRxmLOve5OX2PfStbecYm8QsjF1ZZkY
YkjlcjVfHdpSwrkTDWHRqtIN2mzvm/i/hl+4FEJCnoAkvk13AoTIIPNK0vEgqtm9A90I7iUeGmwz
jIooTlMxFQa9JcQyp6TXt9oKNG1aqvGMWkAYj9lVqcckMNNehlTaI18btt5cFEhmiuRQrsVI6MLv
50Jh5zhB8U78NewyNftrkJLG1w3nfCQSolgE5SPsIWHlKChH1rqahZ4ifTFM60kLApnAA/d3HatD
EL/9c7ykVH19gviVcxIYUOzXBihnOZxzG8pyZXNEgqh3Nv0h859GLY5m8XeAh48Ngf2JYXAA7lUV
h2n/1zAKijVJZ4XTWHCGIzl59Ac7Y01rYpzd/Z9A/wXDjt+ey0SsyZJuu2hFXrhwqxeeVYZ1y4tz
dZhw6cxeAFLadojnlMoWBj9q/b2kGeYhG+Td0rrZ1D88PCgUj/XSVkBptf4/JKBgxCRbzWxw5Wzt
B/BA/LD/FmSIhhZmaCZQnipdye89B+NH3W5gdc5YaNFnPDdSS8F133Xucoazw50I15A8ouYZ/K0r
eOq79468PncpPwrkwhuoNRK/M57nIZgtSc09VqeD2jVHclbrf3iYZpRQhpl8wwxVIUTsGzkab9GG
vp2Tsy3oSGlem6nO5/sFYrcPc82B4B9dGhZp13eyoEEWzQoJ6ZoKhu+QLxhI17YWy9qJXgmet8fI
tD62D1ugUPOLSYIpTzXxZxg/tvQKv4mQ3ydnnXubEEHFTb92SSFpX6G6i9uUrginO4n31x8E5hhb
zQpMbiznn3s5R640prNJSIbOZLDH1SfzWN7co1iSNpF2I3ujWD1O4Zq+Q+fbtketZNAGx0bninzx
gr1Bhob7oKbvfseTNdtSN4LF1h3t/86HHLLNKbc7ik0ZVmmMWfCl2tVMQfcilNWJRPiztocmcei6
PBXbZtA0cYHwVl7lwZ8mEdgzk5hgLg7TSGtHuhkezgDtzEZpoMudwYPJHiK8w2G4zG0VEVdOcP1C
bkk0+vV1HlugG+bqknZkTwyljTQvgabEQcOwFwSSaSe5RSMr6YVonYZmkO1I/oYSiQGYjsGgPreN
vJw1x7MAeNn9F/n1XCdI74ywnKZBvqnc3UzeaRjgj3w+FRl0sG7VYg3CEO+JwnxaHS3wZ9N/wyl/
A3hqoBP+Q2EOxpeptHxrdrMvEV1FSQQfYTifutyKfzJI0Kipe0YSzYImG39xbMxDeTahN000cQ3v
kl6huIlmeK7dRwQJI5ZG+rN4eVEeSMxHJ7t4pOu7THaAukM2sRCw7axvN7hSzkopeKqoUrIWr3iO
s3w9IcPAgMlD+k2oBUXRNgh5NzbPIk2lkY9UzDwIamDII9eGpYiK63rDCD2TEPMdl4fm84zA/i7k
Q9k14eF3JgNXxZMY+QA4zDAAXco3t8zo+AgE7QopoXt/Q6OuwAIoOUgo/ngLqzU2N50Pyk7nP6y5
D+fkjoPFEkImPsk/MT/POZVj+rGDE8X4VmwvxdjGSXZV9MS6lV9V4LAl6cp2xdYiYjHq3/IjKXae
sSIB71cc0GBR2BFQKWehKum0vI8RYo1DAwlNgF910Y1UCsUNjVzxvDialrsP7WRn5MA27SRsDiUn
qdPe0RAU0A2dA8aflTm/hRozuL5Q0/G4JghJdPSlJnoxAO+yBHh1jEA0CnsG24wiARhVvEDvCDsG
GSVVFTd+YbTl2v7JSqr6+lniJGALP0BhH2GoBeXGXU9e/9Gifgyl6+9eTxdCLAJVi7/Y1DU8YSkb
2e5ssBdNPEYmW0dnUSurzk/iA7rNJDSgwISME+AOxHl8dwYvdPAzMc8YMmAsR1zroW3rwYAo6oL+
UKPoA8USNxFvgvOF4VmEvkHsjkfIXiFGZbwQghbET3wqiRe/Rr/VDhlfZ8Fh0wcGaefOhkYAX1Ew
Pby4BLSzuqhjgrvxxnlO3biHRTlJk8WfeKHi9d/b+7pvXijy0y6zWZ2ME4HP7kgB0MSvNqXmahpr
x/STN9hZse4BmS6IICUjY7KQ3yfk4wCp8j1wvokaWr9trRrcBb+bIkbXHmYcsLoqQglifHDGJ+AY
xPQ+7mxD0OmoH9HufR2xk/E0sPykJsTuZWbQVEeqpuFd2TvVOMKbZoRXyaG5cbC64GXyWYH39IQh
NgHyxj6reQrhtxtUKhp9DJz3rE+zAy4iEq9OBluBLzbuZfDg9Q0QcdZAN33plJj0vAFvYwsWeUor
xsFo85RIwX9nIzIAdczY9xS6VqDmq8BoOjx5J/5DzJIbHdr7J+rqC8eBVzm3uvAE7mXk/jN20tZY
QhaEM06K6FOkRgZv65HEpuoUY8h5D50Hnk5KRIXaTH2AJxA344jdGtyewQ7uDiELsBt5NWeRJpCa
Zkr5kqgv0CPtzsP4UJVvm9upZmMuQeh4CQYICCu2elpzHB1x5MAsAaeIXJWjwHzLq2OsKci8+WzU
Td0DcsReKdLBmJEQmPKNp4HxOVxUwBuYijuo8016EiOh+Qfv2GKjAAPPYrONFyTM7I+IDDN23ChA
b6/d5AakLQqRLGxq7muLSBl5a6+ib+P4zCyhKKd/2GwBr3QYEuPphF1Gjq92Te2H/lUaV16FkclH
0HpM4MTApi2K+vy6V53AauhlqvVSan79DIlF+czsZ2D5qjil4Kjrbgqgj2hpH6gGqzZTjuYFWvRN
rapB/jDx3OCr5m/Q95CE2TNUyRKWLkhiFrvDHA64X4/9QXzJl2diNqsLoM+MidhNUcjH/JSzKfVW
CiLMoFND5tZ9dKW+hJrITcxnbagFP7ffkpI1bwqqByVdgqdMybNnDxS8E7WYBCGh/Jic/es+V+Cm
ofxmFeh4WGwY7tU0wmVHkpqj+Bwj3cvs72IwuOyaqrUgIh2zWlLu204vaV12FuE48kr2LyB2M+vO
A/Jjz2OrNJJwd72PPPDMpCdNyJSihkfshsgecrK/cTrh3UyHajZMYvyrbE9gQK1qoQF0tV/3Va3q
DoIYB9KndoquslyB4DCTn0UFRZQmlMLuepS3tM/PtjQo+wLsaJfsi0sb4cOUGkFOVx85zCX89gPE
kuXeJVy+sQzSvZ8NlE/mw0Nig6Cw5e5f9pKc2exQCDNT9PakyWdyKR63pkeSNR02NPSeJmup+nHA
OqSWxpBUDL+awVFZC6nDRH8qb6fTy+spNzof6E4n/byX0bf5+KQNJywL5u7l2SoB9MtKWLC8ySpQ
AhQePE9Tn7YoXHv5t8uDxE1Pj62Hcf5/EqyNoqiXx2HuHVuTaFE/2bBJJ/wQgWZf9X1wsdUjTJUf
uEifo4Y3h+zo5pvPef+CIVyON4JUQKd2orWKAlSz27bYr81KkanYXIQ7JGwfRe4TZ4+29uMCtBPw
fr/E1MKOzpgh1mqKQeiyRatMEJYlbfC+ppMrn/QGkQtLSf8TwSKgikrQDmXwQbKCg84al/rf/Csw
8miafivz7LWyZU16CJuoGMqQ0dai/X3VOMBt+xwNYwsBfdVITXAiCEB3B1Uuo0trHcuS92EwNrCY
YZFqj3Tyq4TWUgFKZmHcH3VwMIUDmp4wVxTvyUSwyfLtut1eod7Qm3rjcKGyNtP9HufRZrvjIwj/
DyGwL8w8oG2w86vQAy2NInTOOzBFxFymQOxKcLgS2qOEAqgF7dxKaibVcfyFu9NSvonioKR0YJyr
gzB7n184ERpUFgseSQ9Ej+TP/3ZM5uFkoCaB7bh9ywWOSUESkp2JJ/A+iGRKMj7Vy+InV1DQDi1X
Zd8jOtlxc4+G1uj/75jl5FtBrJ0MZabiw4FzzgZLxDEgbmA1mh00jEviyp1dNF7vxSzzy5bQ/veT
m3dgQposq6cwkkQBegfHsDlQAf6v9h2c6cxWzXaalBpBa/FHuu3uJaQ/gBUKfrnPEtudPaKqjzyM
vIPsY9Vh/ujGbWPaOMaCvbY3D5Vb95W8hOMex1EBzSNDJqjvk0eX2YmDCkUR4XGvS9Vgd6zxLnOo
32ARgDb9nKfxiXtRUbCEHlE/T9M/+V68UI6Jn9ximJIGPl8QbkCHa0Z1d61Qmy3lCGqbz6qyDFOn
090PxJB35ozUqbvGzXI/TT3NTs9ZjsjJn1rIwwl++DPGATRSsOf3mHAlfEuzG+GmgEr/OqBNkorK
74JJGR4Aj+AjHxltR3eRl5P6QOvzOaTpYh24DI4h5Of9g0GRAs3qvoLrSvR5MGySekb918h9kw9J
q2UAunORxUcBom/Zxbn3haAo6ZtUMyqfVsXgHZEtHpMAR+4v9l/3Tve6aa947Zg0dk5t1ya+fBZa
x+/Ze6kK+eibRjXLdBNdvNUDsONYAvFEToxu17xenmzKpwhfXUUTlN4oVASoJT0PpEHWVIX+y3PK
BKLHbawIt7hwRDsNenodICQlBtVeCRRl9KKPH15iVJBts5K60pEmbBRT4MR7JlE1JMowIIAcC+/Q
iWMOBsWRqL6phebPIbj87BUYaFKBlI7Lg5JDAccvJARCqNy1ZSRJ/gJR4SeUHPjiBCHdGhjMDFfL
P36CcN4eIAY92xvqRl7KzZEibLalf0vZmZhtxOCW8gxikJEDliVDSmX+rG/WKMCnMVw7NvJWGIbG
Kny/+E6ntUxHdYFFVSRVukstiBsg06nwTd1fVDbw3J85AfXSKxqbZ2RWIvyggEw7ZwaaD0UHj4Yg
4JUDwWwJtbpJwW1ZjK7iM3a6jm9+Od6RP+0f8h7GAci36BMZVmklS5tV9xjJ2+5OHvQqBF/x79B8
RH8+BoEjIs2fXI7NzRpphAfAj04X0eLr5nl6N6a2esUXFpeRg4F59d5FiXCT6L1i4es2F0yuntxH
AnVT5aNEYBUecqraPODDNbLyz7xsZG33LDdprRvQ6Aj+pLP647HfzMAFhPpvKlYTJ0c3sxeNoAHE
x1PZayp1Bq2l1Z8PZ4JBO/o1rIaJmX/F8Cc1mDytYy/LXVgs84WXEvKWjt9MuFzA747UtpTSK/zR
m1pVhtm/UJViraUS0+XGcBWOncKLBoZOb7lE3b6abnMpauT8aIxORk5dFPryVhk7Y1gdeb3xG17b
xdytcPTKLRGxDMZ1vvY/pAbDiRbYDEKacovmGM2dlWEA0IFkf8LSJCggG+Lyd0uWvowGlvc3aUBg
ewmm+ye7IHwYYdqDgsKyqmzdVzpiQCI3Lo8P2AUIz/kUvWV3uSnDz5yU6cSP10jh1m7apoOagZ6s
VrLVBfEK7v8KIiKuqskkfutNc0vvZr/HKJPXPds4+9emUBFV6o1DBi+FmHY47fMi/3bBt8DSz58Z
+Y8E9OD1nD+ZTO2y3O8I2VJUAu9FmehhQU//qRyLqGRkeu5KZUT70zRtDbldbyGlDvYX0q5+9Vwg
8j9nkW6Iiqxz5EiWGOrXWOWnsqaDF0+m5CBw5I7lzdV0fXOW0F0XI6Ac85wiLwC2EKkjRo7zCtzI
UXo9EHDDRQOGIgfesG2404DJD59c3fADvsrFoM9euK1C7ISE3fnpd4IF3F5aRel3F1c4WzibcZhZ
UWeRDcVSNi9Bk2oJzUtHZ4EQuPGeIpn4Fdw+BUzU/UuGyUw86QHXmD6srqORpj8HA+Ecp/s1xJab
0YhyVk9iT+h6OVRlg3hFBi7GfPl9q3TYUJFKHnoZK8j/YcKMQFAd0wAzADzxffKXIijxaQKppmtI
VwK1l6w3y8pfMP5dkqdLZmHE1Nqb015HD0R5a6qdV7Wxh2Lyd3S4tz+Kg1IgKI4Bx5h8hYsMWhb1
fCl4UNRuXArJViZCd+LdnzNYAvaALaOSp+Y+xrdoW99geKbYv0nx7Bo7ds7OjUORTquKbE81M30U
Mo1yGjutIwjzZtugNTvh2nWBSA6lXMZt6R+rZ7hZsKD1NMiYS3jyGZNpUr/qSBBQquKk7BrdmF2u
yKrifdYyGlB89Lq7i3pbmmHz0rV0wz6nkStT4gAN6TSUf0iHQOs4OmledLlg7ojvplGceQTLAjMh
oJ6MAftMj9ZKoBqCZX0KSWZBdOJn78U9xPInpngTxxvyVYo8XU4s/fr6hEJnhFO0e5m9AtY/uKjz
LphTrDHOZtmupB6T8KyjWWLxlGqOkQ7aR3JQcEYQURn8eaHkmV65eaDjmpGqOJdS3e4FniLuiT0O
olU20gJpHVXL/3Y9GaoVWNElzdKCRL6Yo6nevcVNgMt0y7d2oMDa1q6quBZNgN24nduKqgB3zsP8
gWWinguKhU5R0Ik/xDtw/GTXTNuBLtNrFLgvSACgQ0m/IsxrIQG+xbroY9tAnJhaIcHg2RLD4j5g
l/22mfgHgwMxQejbuKegXPbQrE02LClpyYL3NxGaPFPGH/3+ytOuYvtxpG68IfRgfTHMgUG12OX7
ZNVMdnY35tN1vhzpjMlCRrrJHAhHNWxQFGFL7tal9pV3vHhARhk9grrUdBzuPFG90e26f+BmTxSQ
JCg99tDXFmRLjAOGEq5ohts261AsJVJ8mNrU2NPz7atxhnBFWrBIfch+MNVv8adYPYCcObc9iNnP
JFf15N7X2nOzbTLc/GfKE4ueDCRx1jX8ME25gwaPSuTL7o2tbx9+iYarvFV6u8vHSsqXLEryGF44
WtS3XfPhGSc1EfwRFEHH/5uTOUqLhLe3M+ztodo5vdwKzwr592Q6s+R6eYJ8nIFjjD44zcCbromE
4/fi48xhUaw/9jGRfjj1Rc1vJsO2I3j8I+TkNaz9YfvM2TOJc1ML0jW0cFq66EIm+JAjI8pjTUDE
PvX5s9gGVMZ20VkjHpn6tSGJCqwB7tWw8JHgdFpz81Fx0lfFi4j4QpMzv2/10svQtw0hHHH0IE4Z
w+CE/wxrrd3AsnAqgaQojXJAXILFmVUwTB0lcnEzQ4I2Bce0zvqExiTktAHV3RFEqNc2khXrhanU
GHpnPavpq3CMmCxx3QtFQD0VRrznoIT7RarWOs4mkV/3O55Y9mJbRMaSav8PMIc0YsIDc+DkKHjd
MNLcs8PPwpv79TTBqx8R8KohGT5CNhSj8JA/oTWpsBd1j5Zp6h0pZbpU59CXk0h5fSI9EIZD8VDG
wK7cgIeTrs58E2zMbvqiRcLn+Pn+zJZIPtAHcqHgZvk2q4T9hBDFt5yAdwLM9TBggnS3AAOL6n3j
pjG1MF761z/p1eh3HV8WsWmiZdxkQKGQ0c/s7BmRC0eTX9WQlR9WFFZqkNDleZikRpV5xQqmDPJD
8Hmx7xgg2dPzyWg5RxRpTJz5/2khHNawHPOpsYYa7Cx6KkeETZuSY0qGCNdMIo3YGkn5APK36rOm
vK28H2DJutH45GNVx/BbCsT1rJB1dzZUoraAGYW71qgvkqPzABxIn9WCUWkh8Od/Gn62GYN6hleK
gS8CL7ssu/MpMmG018YqdeQoJViiX3KDOpAKO4TP4kIDaDHruZCPr3ow0RpiguJzNnLJP4XexOTB
JT5YKOfkLxptw/pGhYRK/H2zpeoFqFodkNdg5bOAd3R1IDCNsJHiEwfEF17yju4vFWGrzHVa+I0Y
w8LfU0ItAQuwlvjANbcFDNujMsyp03IaSSwWIWpXXzY3zlP3KjZMclMZ4K/++3QbVNp+4kdV1eHs
gejoZxQZX76TyP74WGiMBfVrMl5FP1lUVdWt+1AzBvdHPWy6uH7st++iDCYAXzlcX5bWvaZO21zi
RYt+tayqDlQH6HcbSIDotN3OkVKgXmcfdIH+0viX6BdTpmM58+oadi+ep4UDWfuUMUKDOH3vlS8v
yRkuG5S19PWucPCvnj+0W2oSXY0TWhm72J3eT/b8QdSMsCMGifUuzKjsZsAw0x/vJWp8Tfi0oPVF
QcOPxb42/2N6nRL1zVZg+dSAaNtXcEmq+Q8xJjzsrTUx/w9EKLe/iciqVA5VvfMitJ/oriY9UUlw
uNEUWeRQyjLFXO1hATckHT8UHyTC1kb5xfn42QcQQUwW+MOHHmEFdRPLUSSyGdPqUIkczK/nHHeN
qLX0Lf/CuLNA92BCUkF6hbQNANMSK7ixpvymiZCgS/EDU5RFnd4nHusF9zn9FcoTEbg7HryafG+2
IO3vy0oetlGoMMypkocYRyIkOY2LrdaH7GWS8dsQ7qoNrHpvws/4r1wNBcmPRLXs5dTG8P65DyWu
t+u7MF13IddDpRmD0Fpbnh5azQ8TIQwXvFY5GupVU2FfeyQhM1/AePGcwZFOWN+XO0WvmQpOD+7L
u43nIUK8WWEGYDMUxzdUoEhz70QPqmBleC64SqKVnyXgLfN1vAHu6tIRLN9zjmFtSHWKI/i4xqeV
qfBtKy7S87Ictu/kjSyJHzSwb4OKP+xYAaQjVFZs4tP6KGJbj15Mgph2e19jx+n3P9gbec6f6GwN
xl2YztRbS3dhEY1jUzEEia53/4jK1P+kR7Lo5b7TOh5Wp/lR0FZRW3VohSmujZdgIrojU4jMXJjg
EkXUxUshAm2pm4bprjWQA4aNVzLh2IGfAIZ/1UXB0qkjKNziJrxgLci+ehAl2t2nS6YDIjRohijO
+Psc7c1lgjXPagp6ewmQc3LsCOcWMXezPR/rc4l+eVx16Kqti3lDmolGjlQJitXZPw0CPXHRFv4A
lhS5opwydoTRVQ1AkF5zsBeuS39Mq9w1bw9yenDMLrgeGkgIv8wjpG55MkSpFbD1Omgxh5LoK6zZ
MrTE9dCCM4V/Wlcac+A1JF1AJ6kUvxrWvCDHp64HhWVzxhtY61yahaFUBBlL7Ddv33bhJbZbFQCM
nPamhQYsp+8bPYD1Ucf33V2gZCMHEoQB3RV0/7oHwI/yp2q5lmzQWX2sbQKIb7brxpZ2a/CAeCz3
ZfuUrCoIFLVkV0TdoJZ+gsqKlt60PvfB5150lMTNB43EgL98bjgil+tcA/MVl5Set682EMnggCU9
4BD3Zm/sbTpRgRRvPMsGJGhM9nSCoVgBA2lXUtciYbh3Nhj1nmsvlgnIOi35CCYTE30Y+lkKBxDn
m8oArfKYvEDY2FzxVInnLqi8azlIH+3qdWngammV/2yU1PP7u9jp3CdjCzMieY93yjnFlgJ9Hjmd
FKFFWBaudGEW4SgZMJCJbH57B6BOdQ8/dLDc/VqqVyu14nsR0Zx6QOTMQ55Ivk1EmC24vYZFAXSF
3Aqq7kpYDscEJjkmS8o0nPBN4yc8zSRsedzR424aEkrM995tr61TGbnvWVfK4//R0mWm+MSDJNt2
SwbnSxgr3MoXxJdLIxwzzJVGCE2Y8Zk1sI8Ed7Y7lZIDmT8aOG+7bpVU6XeoI9vJ5hCAaDzznA+a
5IFy7vrK3IimWS5c7Zrxhhc+0Cuscd34D910Xy/xhZEfnJlW1eHZAwnGjSGW2dT2/WtbyQprbE7R
y7pe6XQ+JYjCPK72wAhohdUTXN34oncbC+doopPb7YjthVQ1/B5vI2ynO7aeSfijyinLqy13AWIA
EJG1BclA1TwuRjgwe2Gh3qDsfLZJuGmDsVUWPVvECWwcbgzlHmxngY5Bhch4ZWR65/4lrGBW+boC
JdKXhgaQLNVSsEm3o5W6p6n+bWuOZaZw/p3HtvAmjlgqGSyolJ1DdS8Vxc6YKbzV9cIIw0zVUBAw
EdIdI6Ll8r4L5wlO+Zk1LHmkyEQmtJLR3zk6AMRiqu61LBnTwuclUdRYAPgYtWKuxuBfWi68R781
Amev3iMuaeA0Z9wtuwM8Bgq4M2LGr/SdBJtI8MT7bfpTjMEy8CHMBtKm0trzsJx29NSWccZ7XMff
xKH94bLcxlpMGxJAt8tp0Hwb7EpNVTrOP4UGDQtqmrN/Rz1BklzH5HP5IMSQMJcpl0tDHAQrHaF0
02SUdtn6Ml5DNcgCQN/7cR/21Gf+ZZtNnDFd4k8+lK+GEf8tDxieBFZ0Q9yiY+J3f4jimAPUYeC9
49lfZ4sQ89aWt+bICjhU/apJFoedoiITGuLGU1nOK8gVk5lNgBvSdHgJw2WjdLHmwbafQgdwiFys
S5JrFNoaM53bY5CqxpcHZLRC5EUwOW50UX1ysguRaaYYO9MNhRLMSgc5wChjl9UC7FLPP4YNizqB
fnXDYQXWCBZ1VACAc4a58XA7YekYkRrYo3KAP1iUBwLYT6V7j4OaC7f/bkzJrEFVhq/7qxYrAJc8
zuDZNU6ftsMd3rVmpzS/Fx+POYHZuOJly1KvnWJJZGJIw0oxbmfqSbS8JDEVBOfYNk162HsjmHXi
INArZbQMFL3PINh4dmQEFKHfrJI7GToLZteqjAoKfSyCWO/pitEDs4JRbNZ6DkukVPLA2XJpQkNM
cuI1NRbKpzmEVTQUHpDfBj2Z/+SCKMJQGyFZHTTcDdWZPmVapHEmrUOvU3DpQ5CRXKf2occtsAUC
jPKLLUArVo/gTUzB7uul3WcirJ1CkXXlc9esToxm8UF4sXxB7ck9MqFlQpnlzmZXtu6haCjHOH8Y
jUkpEdfWNraT3jEdAxkqKXsus/UUXQEnNOUkiVAKVgritgpX2rGW9PyIxA8OSRXdtvVz1olQdS4T
QE59OJNW8tuaol93HsSly8d1MBm803a4Z6lay94L+TPhGgnzdcVfiG7xtaBHpTGLMqS0IrA9zizr
IkNqarHylnlC+3Ud3AdaLV5AjlUbMftwUMiOlFQABDWub5QN85oQt6l3L/gxL13KYy3yu7WMXY1g
5D8aYaWgi/3EMu1mZw/XZwzU6S8Ci+/TgNVevli+FF/9trPJEDx+EmChYyhEm+WhtkkfXz6GTkZK
zqcWBgNyIW+u3aeDUPYX1wY3nuZ/CIa6x4VO56yyAUuLKLNZbOqZHepMVreTzGFUQ8h70kSRYZK5
mD0DwmR82U4P649cP6eBL5HQ9W2azXrmbq9j1LA9A6vzLRlwTXx8/J6g13HrJ+iMBUXDrfHQKReA
U7L6szQvVbAorR9RFlTEcH8uNWP2gIpYglCR4GOKI2h+zRaqQa+vXHTUMDeDiMo4z+NKVFDSV24v
igZvi3FyaWCngYr1fNcx3fSlhHdn5/MeNhJc+Xr2vKW4qJfoITvIFY9t/Hb8/bAHwBXD4hLBhTBJ
ICrnIGAvNHGocd5xer7cyAY6w1+R2VdIqaVZld9800+TAO20lBSzB3+ph5lKOs+iYSLPR/WCtMmm
hOjLXxFe2cCCqZcjO1x4kWl3RaOcnzguoqNhxvjGwBlrhKp7/NfvSHHltXzDIJyj/V3guJfJfm7C
xu9j88iTDBS13Otiwqgm+mwCvphLLzERs0ygDdGjJSzAyX6sZQ/uI3ac0d2iK4TYUJ1dCPSLGRYx
QJVVg1A41uHTg4tTOir0r/0wS/l1Emj6TKPO/MvgfbYx9OFtg6Hs62RT7oAyPmDv9D+z0VzrUQZg
BJw53G4nm0QWZDWaU0/pg45i4wkDc0wj13gza22CsoEf5lpbQRkQSLwnL8iZiHtAGHFBevzqIRiS
yE44oYSt/SeoCqhnZo4zbXffvAj8tpUNq7BIdN8fWBGTqTjy2XTmWvtcUJqMaEEDY56OcJcFHUQk
iGJJpOJocbrEgQCWYQSNrh4hm/vTZB9Xw1DmBcIuyzg8hRk1E1uXo4iakqytP7nY0XThMmVPIRKT
TfvC58FPUxSxmeMlqk5Lrtzw9wB+aUSIo1aPwOfsq+hBtgTJmTY7qY4b05v6wguGDc1UkxrH10Lg
/4GZto3GzkQu0a6rFg2hqaAgmPDZio9BHjiMHFZTrRYQm46POYhP1CNmNCm4rjKVLPPp+dCDEB+X
99i/vNh9T0c6rRme7yFLx0+LBHdex8rtWxKVb+NnMWgYlPhkZH9Vn4dyVRixqw5wq5mx8izE0SjL
M4lyMgd/QTioIdW5B3Eko+ZoqjotXIqZpfMccE8HtIMFRGpmC3RfuG6jFvp6GKG8bShVboTVSpuT
42iOdD62zEvm3wrMf1NhZ6tYHDBUHkLCr4bQK5GrTSmD+GyhEE2rgsBkHKASS29S2t9aSm+79+Ve
rLEC4CejTTojLXANW3SZIOneaFQK0oLUYAxsyKqMY7StUSBLkS6eojISTkhruIuDqrdqFu+dySd0
ypghJbV7bkp4Rq+uozltnh3VHePT8Ghrxl3AIaS7pe7LUdXOfp0PEUlBxGRJz3qM58bXooPKgHjj
n6KdwUTg5xaMHMVQt7yL8E3R92JPUlQ1F9SunRlVpu8iyDk5Qubg5DGVoeEJOR6+owNwXvGCqmRg
3VInnvANgQqepMtyLb8XYyou+m/7YzG0Lqvdqf00GIFCPJDWf9q1dVENiPBhUERmdeHKnjWMRlsW
Qzx68rqgtvzixtZcjPJIys68yLRT4Bjhu4INh3OYjartZux0MLTgAfi9OO45r1Jq3jov4zUOQtNi
JdplV2kDTzoDpQ2DFL/6pXkrPLO8/qeplVsRLfNsKqfbkzRYUyYq8v03Ag9foaoKwjFZprHrlJwb
X/X0iKUJzNwpEzx7IE8my0gZvsYlmRUMtmNX43HYKzDQ5Cq3Ku498Br76CtZUPI5cA0GS+6BCXB7
/KbEbjtJCFanSn16oJb6gXXppAraBXMHHeqnOu1rX0IYukCrDvPyzc9E+85lBTAGSyApAAhaXAKE
5fU3psfUE07zwA4nDjAk9uI55tzP7+NAX0Vg7LMqa8L9f7vdMFlJcZFjby1fDt5qsnZxwdWmS+vg
RKUn5yzYN8CiK1avOHDd7xb9GYWqQXPnGhwSgz1p1nHq1YDH1mHiYQj71uBKw7ta33zSfJOIpeX3
+k010wjtlzseu2mAO5q5+xgerkfzGGmAEv5FdjRSA1jAgxQU1WdAQVcqjozyyAMVBz3H28WlV0Og
czNIKjLeaW1MT4zGahrSsY1ZjAbR1+0coSE0zxvonw4qa4LDg5Wjf6oU2jV/GYgQFyQA38TZ2A2+
pryNDfMQtorVB/C1DHbJmO2TTDC9HiCKM8FTYqLGsACDiZtGuRSGEIiLAC1l85kicwxke27Yhn3a
BjQqVVgY34kJIwLb4A8e4n4XzD/0irLgxIuCjz5mc3uk/zL8vhfrq4HnirEJ+EUNz9kMdGmIokGL
c/S22eDWfKU5JlMswo+AYFznYMKq0vU0EjF2d99tbIdX5CcMG+EnqFBaROled1o1A5f7A3I2c4Cx
hFS56jgcgsUOnVW15vtH+fh+IeWIK45itcfPvv+iM2XwKavskCYObY5OrRyQUnqhPZhx8tqsxp3K
qfy8PRUqmkihj+J6eEtoes6RFMNscrqymzSbNzPv4xmOMrKxtgM4/EuDSmAR4ootDz+iIpSl0FDz
HZKd6HfEDsB67AMn/S0y+3qi0gTNULbrulSQcTopGIKkhqdxsGzApRr6rwKPIVylQCH1AvkQoOYB
oZa/rv+/Mo5HcbxiZV6QAm8VaK92fFJBAJ7tEI3xzzvCE926EyNDlYMyTqOXWL6DMne9DyrbWqG+
b6LDcx/h/vHMvPKyNOMe2Bm7WOaFL6ZBPNDW/3tmNe/7aT7ou3rpBOcT4bScgMpcsia3/UGmcxC2
rUaOBVoqkuaap7F3UmE3ctO6UV4WiDDpj8fDP2/ZAZfvhy9cVn/BcvPO/RBEPERXorwqQQMfyZ3w
aihTorPZf20u+HoR6uxGkhO9cne6ypfK3VUIntz3Bodd6cAEkvUuzS95vYb0zXGhTx5nHS8+Wcm+
UzlfkbO352lXWYjn/yO5VXRf8Kv4Gap19lOmNjjRR4l8zZg659T1vAiGSaJ5pQMzfvvYjbuozgM0
qWOwUsMBTlvbYBaZTuSVCKmyO/BfBzV+G9t3Y8AIBjfG/KwL77rYZg34s85gszMSR01yH54GLIvV
qWM3A0925puXAJGvzWpEmR3oX3pPMSOa0MQKLaDj0JosZm8N/5lbg2anjzkIjGcuIJPHDxuavgp8
Fy9NQ5YR5Bkc6O7h6gFsaImWJo8ClvB6XbWldE/NqnivJLSRX6/cKRaJbJwHTGvbWGQpb4W9GAYK
q/iRdA/654H6p0yGJLDVMCIUgAxR4xjFLLkrgR1abVMckXSjVn5GwDU9PmnYMTXeukuwT1gdeSBU
H+ItopheqziuODz/hp9vlZRmaxsvU2Vu56yXqHFlMNuiYGjAlWwYVcTO+pmXyKcbHqi9SjGhck3S
KLSF+14FlILuUMDLkJg1ob7tkxQn+uMpCh9Jjb8rCPeqt/THxR4CCGma6rvILZHWMRk5tUtGq21A
23fUf1vym1U/y9nQtQxNGy6uAcIKWC0ohgwvCJeLzmdipamBuGq/Ggxe0iNOGQmVvlTGTTpZnDOY
a57gJWigsLSObDEMY7Srg1sSHKkwSDulskfD/lBm44WHLZMOiPYQkH94oHwEKU0UE7wepg+217w0
wZdBDUyJI3KyBmVpDU1BRwQpGWChELfwxsXtpwTb+N5OKB5XBfO3P5p9i/j5+1ei+3DGiL0Ublyf
RVuqpqDq4l1Y75tpb9BBiiGQzQ+9gJQbdq9j+3n6/64CViTQQa9is8e+mvcKt+whh0bO68QHFQuV
gO4ydHcgRb0K6TnPXKZD8fO6PC8wwCb+aZceOzU12UvPVUHUkdNuX/qQscWoW48g/cwrrhi40HhA
EU7RMjIUMABPKpQK83U77y7/QbMGVTm9h18S14lIg49F6s7K0s2aj8ELgIkR3+tnlXIaoD0P2v0C
AanslTLhZCQcVy9/dgrNhRG6fT3bQ3D5BsvIfQ28FRqIodZUpbRfnKaNXPTPVqlWzIeWL0z51/Fh
T68z6b3EfGSsJXVb6Cxs4RT0QFUFFXXcXNDc4YpWeGoHI4yyOYY1k3FS/ibqq+BkfVqqUsTmrrZF
8zud+FBk269ybN1VDSVBQ6Z6DZbu+voBd1dGUsQGdy9XRXmxvrkfAfo7dzgehxAJj27q+8VODuBv
vwgWLu/bdSyBbPplP9pyy/KdDkDoIOMTgR6DTBO8c1TD9WdkTCnoWGXepK6gtHbXL+odVH1SrU8X
AwPrveUAbEUuzHxtjIZuy8FyDNUcON2HTIqeUlePvjbP2Ues5J8GJOSIu+B5LrIBcqWchCV6fu+m
06C45yHZwfs7lkfvcBL0+lkWW1h1BnmHcRRw6Yaw5Nits1pRSL3+cXZEbf5NcJAOb5GbJkdSy4TY
8SiIdJ/5zMqY/edd+GnceJsgKDVCIvZaSkbQ5L2EgFVQl1IQUTUz4Rg2dVnpGKu36WgR2tVfgeea
mBVHbwJP04Wymmtr0YSLDsz0nBaiF5G31wPr9L1NzEshYdf7OZ0yFU3tkkSmHNfjzLUmPLAU/Df6
Fm6O2zYQiEmpLdinp8gQ3e9SUirzbl+Sh4sIAqboUk0R00OvGWhoQR8J8OUe7JO5LhMBMxvCHfBF
8yHafWDxfTh40EkyjwI9sYLDt8bCzJq4/XmBE8oq0dRxJglIWrD4UZYtwSy3p9omfjakLi2GQONl
z5WcKDv4IXxLrorl/9GwgkT8mT7z3SdzvT38Al1Jrjxzd/3TzFukfwTTr+23bsosk2VoIXa5XcRc
Z/9bTJvavGEJGMYW3MdnZ0TEF5huRmzdg+CCFBp9fSFgPQgKxC/zCBH43g1ENCD/uT0NlpG4CEB/
iqjD8pX/tsVE2QJMKCX2NGyd5BCHM/4xz4FWX3ZnygFYvKroArvnnSOwO2VkV0awP3cfFcbvjtK0
bhmZfTl0+KRsvTWJux3zQrOMLRxSRttICQW2CZRKuWaVQR5oIXS/DHYszrmeJMpb/6B16Ir2f2NH
DVQNF7cG2QlhnVlMvsSqPh516cuDhaiLpaucFnHMGeEpHkcKxf/g48KX2R6llwmYtqXQGLXq3p7Z
+aOyaBt64sMcP0mzGscyxk2zxtwZM1tpXjqPH8pyOMyvW7ak8XnsSI7l2kfO9B9h+j2KiDjhyh7z
jDAElnTL7JeQARa55IrDzPRNtdmPG/DU5zAr70MfQijgvIUvruDmRA0d76ISq9M2qypmXKMYJ2FI
Ptr5/TQhAvi6uTcI6/t3HoTqV8qJWDa2gpj2UcoTk5KCXJhugYl0+cRAhUD651OxoTx7RS4ecQt8
1bYXT4DgSZGFsGFQ2+4qqAhYOOdTOraI0IYttDNvyp++s2Cv4UMHLOR1Q2K9rig+LQS3xguHhK4r
tSQxOY76VeWo/BcZFWREndP20lOoPZGPUULR0ELBBPQ2bed0zFIiiyu2Oh+Fvl2HjSe09sICJoBS
4rtDtJGyVpqw5FHp6PqohN6Wozbe1lGUD1N/m/cRY5GuNeh65PsRvO3a6zVhdC5EGjpeudQLFAFg
i36unRajDtIF2WnFhCp23GL89H4Nt0vOpo3BbxtePkSBZ8/oIU/MeuVhRCxxrheDaVujIdC7b53Z
LZp10lE0kRyZczx/t+b6jImC5kEqdfkEC3h1gVZavw4L1V5izJmmrpiFQPAdvoPr1quOxDMdEEaY
fSFOHZQemxtWoPu9wi/6Mr/ViD2AvhRoOQMuDK+i3F4H4B8KAWgw/mlCV2c+7aGzZjZSG+IVqjql
WdjIV8eiv5HAKudB7YMy/zGKl04UI4aCt50dr8y0Z7ydikDIwZEJ62x3bjNkc2yqESo7PXqqbqae
lklRoKuyCFYtrB8D3b/CGHwNOu0q+fIW7GnHva6moIVRnUNK6b71mAAdT+qqz6zg/aQqeXOOOAnp
u9knyckVlwtvB/j+ukK2r8R+QGBUf6+fUrtVB2+cDxUI50JGyM5uHQqdBIK3Z0crcccThRMxKUrf
WJ0s6NUZCiifAjGE9CkZjNR/LlsuVEE6aZYLmD082sTqRcfVrmJhPc/XykA3KJb5/DjSfgvtTvqD
Wh4Znu6ossL0GunJGbbO2Vb6WjOJV46wBpE2CdvYVu97QExaqIjBs9Ynld24ZLrIX/joy9lYCki9
T12eWnB26rOf/yJb+uygNY+r3JUtvtQyKbW6vCEiISuk1Qw8/X0gyfqHQI8IFhV0uJEBJkny4E3e
33iG0mT7pp3nduPPTn6klVYS73f9EOT6ZcMFZHus33dIrLlhVBCgKMVhdenJwgCXiWV87doWqGAK
9TEtplRR/Msjr6cP+zrIlWkQ//20L7DBO0bpG6Qihi+nN3O6+zhmypgkdpjozZ7PqJaqaizloVXS
LiqbWUY5bM+E3VU3ML5zADHYB7wNAcXeyhulYYKPYqSWlO8vHpzAt1DhZE8e/ka5CcKhzhM+NZbO
SNeFe6wkbyiDBCYeKVf22EkEdCoHPgpvarG74C2/71swBDD9jpWg1j3oWch20OUaI70OWdXkQ+Vf
aCnMhN4kpQmdIruRhoyi9QL8MtfEMNCAH4MTPVF6n67szOlDgzu5xwTmhQtG9I0L4tgtTshkXljl
fHZosfnCePJ3Osn7LONbh4rh3xWQmUHr5KQiGalWOzi7fxIKdMlKOE0QrysOANOzMaTLnaEvGnko
Dp6XZALaaaYfFcptJgBplEVUxgK9t1D+aE2iNxb0U00p9DTObC5Z3EeIQAdQdQDdcFINHR+eliDx
JkQB2HoG4fOsFOjuK7km2PQnqYN1WEwFKDnEmKaleiHIL8H3KSGpr/weE4q0jtAZDfCbCYnPWhTe
bANSghRncjR1gfC0aykoTLLO78Q2rBWjr8gjLJqgKcU557A4osEQucVmBfDhOTOt/S27gSVQbT3/
9QPuRze200YAqW3cUhFOsN/ggIjbSqLYHVyEBi2mDBnDFJy9uwpHc6Lh7SG5Jq8Qv/wZLpSnvPyz
BnQXTVxAig9o4OOKhlYegU6tkafZnVZ8WJU71KDxpFD/DUFWJbc0y+5lW15IjKIhs/ozcFPQYzZh
P2xV34+EiwN3vpNxXp2evMdUE75b2JOdBH8D25jRViYzEBHFWFpNkLBU9eb+Kswy/8/UOZ77+PhR
Z4wCQWaZdvV2wf8EoCQ55xm4oPGgNB4Kpp9Wk6yLuKcKSq88YOatFCMHfB+hOnznrD2qku+X34mn
tlmwlO7nkycFePozchjLDKaaELgAWAHLwWZoautUbYmjbpRBuAq95iHAlZI2VbSLNNlELzfTLEOd
212gkwpotM0EvyFX8I2i0OvtNAKbJBnhawMmiBPoLDirQ8h+ca5Twbe8An9DRnLO2CbTnJEKRIee
5qZeGh/wGUSPiezGKLe3gF7DccnlLTZm8i5jCDO22SxOCxUqHpMRhXuzVFO5Ki9saYuCfzpHVUBY
JNf0zXtXFCn4t/0TN+4KN9vPDO59M8ck0Rz8esfIuZbRbWlN2WZL6ARp6EhcdgTpWsyv7omFDbkN
CDUGfgxLIoxQXCcXk3bMkfColRS7ZHGktrzAbN1kestQ+8E2bv+P0ahVJQI80rYG6N7tgTB7Dhr7
g/IT4QM8PuuSJV1YXw0IghQYp5KnrSTp21aMSfN4xQzqO0H+cYFJIu0LXJUuW8IKfinOUsvkPK37
u4Z3WwBAoukTscrND2nxLXk2LNfKRg/+eniJI/uPmxGV6RA0XWl7lMyEf799NxlYkexQDhTfquSk
NhwVLpFPtvuC3h8CdnTJjImHI/YrdSF1gZ/90A2jtCfPMgWblLPB+cnsaV1v82PJJ/xSsZ29n9Bl
WMkISZPZxyQDFJWrWZ0WT2j9Xwt6b3pWkiLC4Xa0CzZAtaziztc62fgOjKwxZklr0HREyr5WWRt2
+hHlIgZdFjMu0VK0epzjA/JQX9o2ryaIXA3Tnh93qUa42veIvpBuhgdbPrH/08tdX/x3WuA+kIBk
B5gCJaMQ8owrqX0qNLP7woXDLT+t0lftoP3UKpVt3QOnlwam9hkLf6Z04oFO7mJ6bJcUTvBKqEpe
nGRoYlwjn9sUAjEjQQEd0R6LIboJibHpGoVJuM+7JJDOrk2H6+5JP8JJvjF5gl1ppXAXZGQIBlRB
PG3GbVVNYN09xI/cU0raZyJo6g9vHocTck0lURiHIEgj7l0kLUelIBa76Z/ZCzJBbSoMCReAd96u
Fi8vXNYvXIUnAumU7nPj7KwC9+p0ETbg/yVVj8FoDDl5vrp8lZM7cxNM7SV+Alsl01Zy3PMMDpGr
v1k0vJ7U8nHAzCrv3xEFcWmxqFdSz8yHfx23BvCpkgfzuaBXnv5k5+4PKcuktdUFq2xrCaGbktnP
iK0Xn1Qj8sIOB/6gEL4amasrdloJbR4ApefEm02aL0UWhlc1hNJSE/h5Oh/5xvxMrGm+AWFkK/uK
u0O5W9fNgvZkOK93jxavoJDfqbf0oe20x9HXXbiub8x0lfPKRSu3xhFliFH5u3PKLkcA3/+opcHJ
74ndyqKS969ievoT12QEMfZE47MdGqWNpg1U/kDH9RO1kvxIPidiWNpY3OCF6egg534k/OT0E1Q7
cF6ObdrWEdUD9UdGYJbxj/ciegsw68/VHVF3YkDN6HNUVK6BkrL6Qz8g9Rpz9HwbEZ4/BtI0zind
J7yaiLW+V1oLVM0NfOOzB5O8BL0ROLuEAN4xY1RMUAcj7KYtVbpzTpfWD4hz23TtGknXhAIFLnt/
poRou/myR8exjbrmJj/f0h9IwYd02Qff6/dNn4U2TBQNrDmFkse3rE6WP+mSkYQab9+HfwO76jOC
olMcpwO2h3j38fakAzxljPtAQVNAX3bc7LWoPtbJZdQGzuL/k3xiroe5ejqLq8c5qrVfpxf+3Hck
WMgysOX6ltFiejontTwksBeIGGRf4mWOvg8DTktkoRSwrzA7xFGm99XkMSyyxIFW7cSUBysASFPM
MXvR7SaK933VrbjMWHeMO9uYcwGU7AJnGXQjfYNZQNYi/2QjsMcUor4M3MpLyBeQA8eAjxpacL42
nJzOJopWW1gIrkdad4S1FJJfxEcx2QnBD3OOp5NkPlxPDvEQd45XefgH5YGXtUCvUt9BWWuDIsHF
i4ccyghyiM8hSBd2+OXE323Ab2t/0fCabBPikXqxohWqs2od0fjyeTvQphaT/ahulaRzQONgkd5F
tAkaiHhQNqQkDMkQdJ3IwKpScK0yqaBP4gN9euw/BL3wFGlYO3mjOrEJ/wL+1WURnDfCf7NwAGnI
H7YQntGK+IjOO/N32IyKUwJhTCetgir5zB9n0o768p+4SVM++bTO3BKJsWcuXIYQewnq1R5WQoYY
Vyez5eevIfyybjOjldtvgb8ADIW79B64bjpq33vubgSpS2IqZbbLndP0NMoNAm52kvTpICnzwsUG
LeyijrIeVUrrQAKiB6VQ+hen/3raSc5R8fPIPQ5swdjaxvWiKnHb8CHV3aiVJQNJaxw3i/Bnz50c
6S0R0pqnfDmuXCc5SV/soDkzeFMihNzxpiydiYWOz0yQVJNg9Fr8DJ5AO2Snypm0ZVeQ7IU/x6ie
06qJ4+lYeM49HIvnbU6pAQtIrehJrprO5/A/8dFqRlPgmKFRYWegQCecIGojmWuk+b8mEHxhsrOc
lQU/pkB4ks3pjg4Gwda0BMuGrt9vKpEHAkmgMatRGgM0XiGo9H7YoSqlqMonwnqL72dGlbo15dse
On2douCrKkaSr/F7pNA2CPaMcibRH8ex+QBNtPpdbpEavkBFCUTuhmGqn+DriGufr6ESyVTHR6G5
qYkEF5XqLYKp3uDvAaKBzuh3RCA7v4uynHQyF1N/q0SNJ6HoXR7g5w+bbXVuUZRCbWCbfzcAxzvH
VA+UUJI5j3FOUGpSocTybVXyEznGJXSzuQ1I2HSz0EbGq8KxWgrfUz3JK4qUBKwUCyUl6zP2jV17
dS92+/clOPameQcyLGB7G/e6xjs8QkwDqqasoz5b5oHWjAqOlp3C6wPpQ5ashAABoRwwNPZSagRq
27y1m3r3MPnnBQa8TTfL84Dr58SHxpivBNwP7RGwQQnu68haFOXpcqD7+3DFDwkHJOV41HioUaWg
JRxgxICk22YHl+H6KuF6JnDwJVMCgHM+Vwi7sP3QH/Lemg2nl5grBtFEhxjvRcNfholpblsqKOgu
mOZ6fGP8Wm08xWrul1HC3CxQ8q8nP9D3LC+JdrWSXW6AqlaKlfwwmPTHvDHfEhY6K8VQ8xcmL6Y1
p9gt3TwlboZL1JuazLohkQVX0VjJ7cRt5onicmUnyDy8XD/AKQVK3UH5CCF3phS1dfYt9sENAUvE
GQpbNXutbznNxCcdZJlRgV/GyXrwI77myusfsrXAju9/LHXJ2siubMv/CitdYzFKPw2KoCAn5VHO
gbJxA9Z+BsIw3IKc8XOl7tf1Zuz5SRosWa0NHdeFLkLyaGinWo1o39knYW5fKRHuZBTPJJPNHMXt
Z8FLk6ui33dSSVrweulvlrvHydU/3xDoVADBnnc58957+SqpBwec6bRYaqj96udm7q9O6AGD7g5a
0rp6BSmaqcEXXiijAhBCzpjdDv9WujJ/7p646Yf94Q/YhQGhNdl/0kFiiJQPyU9AO7z73T9NNYIG
srs36wXs9LeywkuNGL/KHKPZosGhc+ZbcPOEWFJrZdNC0T47+CiCLi5qapgMa3YgQE86KUCJAxrl
pd1oK3SkUVBmHwrr70T7ALO47yqM9ZP8oZLTFzfWMyLEDJqKbm840rQZP7MK18oEvBspHnUIJ9N7
NFfGt6YLEN0GHW2trVVMcCFOpGJeO3LCGyHSjhkhFqU81yQyGYy/Bod2PMPOOJhfZFa3PWzdcREs
EmRGMQtDtvXR9xRsNb6UE1RkPMMwEFAZZjxeMhtbsQQVbjhUfFZN9/RAcrSO4FyNOsLRCFVO/kUX
sPtZBI6V8fhEYoLXlGiguEYdWiqg4QkeDO1nPcHOpSUEgCrI0r5hXiukmJ0P/MgEpWDDOkZmJjHH
0F+QxBTX6PoNhuZD5Ih5TZ5T9XZAnm4yPePFfHG5x/4bySQ3NboTJyCi/pISTpY6NvUJ35QGpEEj
GGurPFi+vEuyn4Ft4WEA6lAc6vNS1o1bWuLaoy8b9TthJD7W/kqhkavQUmVmHQd57US82yZKwxON
NbdTpwbYoXYx90hxAETLIN4ZpR9nL8OI/mnODQBuANm9weK4R1vFy9juhI/wYbK9XVJk6FUiPvqs
6XeV8NnxD58E5vZyvvgJaOLplOO1OBageJRJHzy3ABs3ujzwV1MDO6CPpb78rLPpSD10XseZs47k
RpDWHVbUIKyRNddkWUA7NcRneZdtTgb57AdG3fwNCTNOgpyLbzAszru1t3ivAnSKrQ/21SPtfggc
+GzjGnIaaSKFZtpWW2T+6Pms2v2shfiEAmWYZ+PHFMY7Oyy6LvBzGBPmdrTPiar2z/ZO+xt8J4RW
9OqrJsHPcTyDo7N+RF2oxOwFoxlchNfIzPUcjgNnkY7Hjbcu0fZiGFUthSb7Kc0o6pjsn+mlrpGB
LjNCXJeaGPsNQgNNYB5/sE85djuhyr691uPnQ+b2CBlPh/B0mtgrscqDonRtSTlk4XkNPg5AqUQE
1p8mlOi/ipOjcsc4CUi7SnKsAmX8THF+7+fHV/AMLdQTgOk/0pUZpAQkG1P4P4MixI/Oz50bOeq4
VlI23W5BejFquaVOY8TgNhdk2Ri8ioHEXzw3Om5MTTRqF33ERNRyArfO2/WysBCs4Y7XJIgXuQJB
cBNoRVastdPUVS2PYZrb0nXPYV1ZksNtvMDKyvZ8UYjv7On4sxrQx+2DGMCiD0mI3u9nPGj21I7N
lvZf9OM3FrIBMv1oLBbxe9pQclWLJDn79A4R2oFmY9rlFgZbFvhHPvpY0aOFjfufxqw2PVd1SeTj
oPd3F247dIIQox1bm+dUT6Y27gBSG9yfmWPuVDHTi3QmlU790YH9wiyg88WiRC0Aq2GuNyipxJrL
I3W6e6kOvQOsnzQNOLIrv+tzakV/IRrucSCcDZkuTLrBcS16EfRedrBs+lOn49vx06ay4rOT3vbC
8URlRFa/TLYXy+RlOVYUGQLehWesZUB5rvMBjbw8pLf3RRP2LptmW8P9tTr+WRsOeo89lsulsOKU
ciPt+E/3nTP01j2Hohu3pru8ccR8Dwxn3o9SXOZmKjIYM+XfBemJT2zTeXST3Gy4m6Hcd8mLEgbt
Fj7iilISLW1p2jVFlYh+FpaqD+ZQeuiNHo0mGzVEZ7V2sZg1WpT5Myf3AurM3XaMnc9a887ZNqQC
QlBKlQ9gVtYf1UmrLAan0Gxb6m0ZmCD58GzkArpFuVYicYA7/XDS9RqVe8iutNGgDAKsgQbmS8FL
xpIetA+ewLd3ZnB9y0D4h/VgpPS8SOxqGi7ZelvkYhjRZp85tvjXGqwUsNJWY7IFWgnbmwjvVJtP
1l6DjA7T4a7qIaA3I5RGbf4wvvAPDUtTDudVUaHPecvwuBq2BXtvfjhdQ8Dm5nU/T4UjPZWKHUFb
4iEGObZq19SkIF+s6VOhVELyknvIPMBC9MsGwAsI3ijwWiymJrM8xXzfxaa6YujVXd5jKDdsSvDx
VPhaHMTQyg8vGBoY6BQNyqGS/af1ALqBMO5ACLm/m/k99F7FN6rr5ZuSCCKHoH7TuwMmbqFYBzDw
Y8bBYe1f32rG+NMfoHnt3USeG5v1Ux7ZQUHbNwXSUzMOHcXg4gxoUCTiiLxCw80GaWtUb8eFcUoy
8z+F0IqJ/pkgfkt2f06ovVpplmNVx7EGpbpQz3dJ9Rkv2IYSV4MeB7VYSmzA1zP9meCDMhu3CF7N
Co+yuqEQL8Ft29CRPK/T3xEe6cR4dEvwDncJJ1COOmvQSCJHdlEMS/wKhrn7656XV6dyHLnl4AF2
NMHyOUWxO/WliHfYAPt8fDi7uonOSnLX6Nb5XZkIiQSeQBFxtICll9mAddlpjrz71Ryh+3MKSz0s
lcD2CjlPD/697hGZ3dYFIF8Jw6bbmUObtoI17/fjKdgYTfMwTRkVrAc5HKSQpW5Hlz2Qdzl7tTcD
rbkiSBmkGRVcB5H83QVp1zEoexaJgn9AHyhctDS6L0uKJA5N6Gg5Nx2VIFyfFof+Tk/qgpDCIsXQ
FskkdLVxULFGDUisP6CNMxwO1okl5l46SnhZhHpak3LWqiWkiRjEuH3+8ep1tB/ngUa6EaAjyG3Y
5EPt/wvf3r2m6nmxxTRbeJkEvTMjjHP1+rfkFApPKfp+rzkyyirEAb/JInbpAmbWDsFrzmiPaKzH
H/G17yuTG1Y6Hfr022GWSMCx42xgIxStwNepQRjvlXMKUkSE4aSA6yTabaGdeviliOQntqhja/65
WpQa8+oKFvqd4rDlVGdK7wbFR7dPLPj4Z9EpIn1vdnLjx6PWzheREmMw8W300sFBWo4TG+QMzGln
NA9SG1T7o2svvdztnDhXZq+rlr8QfaY0mr6QSX9j9DYMRjwX1uRZh8grl/k0gJn+fWgJF4Hc4S0y
3/JfFjCEAyhPKj42C0mVBdCrZvn2SLsfcrw3Z9EuXelhdxqCAvbTEMLbpTy/Bl59wYSTOiHMTYYm
97RPyQAwfv3wgnfXbyRb8oNm7fDQyMBrAsh91sH258WNGwUlXUrw1pThAlPJKYTTvJLVqcB8HY5B
NQoa/b5/pEzf8OTYRrNIpecfpxcAZtL2yf/0PWFNJccvHHNnasAEFltagHFgMQ2RHRqWYUk18kOx
QEhK0F9JbcJVlQXdhqopfC0vLn4n1e4EamrmGUGMbIh/xn7qSdMsN4Myq5L3Yv28QdNnRlVclhEu
9XbdZWton0BCj5eujtv+z3uPz8OVRt/kMktVrJeK+kJBeOEy4E9sCl2Re3O40Ht4pLXFyENTxYPk
x8oHMMn/stXev2SCyQHvhFY7m2IEa5sbuSB3aap4U548079/Zhx3oQ21gyY7Wn5QeNfXnq3WZMTU
hzRvmD/KDfw4BGvurm5P9Lnh3qN4dXUMIieYKCVdyPMNJJDwjniFsRjhyC41G4vKovqD5f1maD7h
ycJyssyaA/m9TeF1OZkzek53+B+aQ7vuISJXRq3lLKxXJ0SFaJFUd8VabFapZfTWukWmSDTNAyuF
6Qfs30+jN6RMzaMdkApew9j6hPi/ZRTpnTGZqEJdoXvZBI6WluXaNOaUMJiriCZs3UNxMRWLf0u3
Rly7bYKix2ko/G7bqEe1Bo3yzGweb9yikFpkgWYqzPbKDM6IufnT95q0Ydzf03p9Bg+W1Ja47Q3w
xVgggfZ4Ry5P8INEVXIjkL8akb1G9UcnuxO1C3tabuDr6j7O6ql9t438+6Uxho/pc5Ehy0ZgIJiY
dDWbEy8eS8qTukFvhlnjYq165mqbg/eNggod+jUWKnCQ2Q3zVsJOoaRTt1+/+Lia+kDsUjzMYoGT
YUZDrfD1hAWz38mpTGLRvSXI/gf89KYfi2sYEHy5RdxMj4aSy/6MDas/2pDKACOhV+9oxiL+ai5A
yDduDUrX0gR9lIA249Sdh1kkmcNFIYLHd9kHjHpgebVd4D+YgL9Jk69qJAh7gIxE7uGD/7oY7Bz0
c9XRGJsanufyzAxAtRdleHtd0Qwv/Yz0wrXiWgI4sgnTHKJKlxMZ9qJnuDwH07BDCGJ0/ZTeNVAc
71IAk2eo9mXdIkmBFLTpJk+SMyv3s657NvvrEdRHHC7vwxx0CjPvu1/GvZltRcpLMXpR45/Wbo24
YHG6WQjF+vviqQFK2FnxcfaYpRlppsbubyMhdCsODSPvuSlYt9ShvXN9xi7NANopolapLgxIh67H
dVuO/9h1MwmNf5BwTolqeu1VCi0UJ7l18wTiuGKMNx3XCLqyen0s7jt/qOk3eHuaXdEEse21gsEI
4D0HTKSPp2xpUaSnLgXyr8QmMop10CDcAOfMM8sRcQeJ/MJdNsO4uCiN5Gv2iOGZKKGnp0cvgLsq
p9XT6bqsQ852wY6kKazlx5p0ED8rUigBmMmuw7/qgTWLfm8xt9K0WmH13Bqs/d4Cca+iKlhpgdf1
UdZkcWDzTtu1FKjZJKYzOv0B9A4aL/nibcFOuVSoLg4DrGOu9Symll7Leb1ITtpZXBn7/UVDiRd0
NwqzlSQnZN3+uNFJy/gYjHcVz46K7WRucQT22MuPzgX3vqyiaEmWEIslm/ihGNFIiyPPn39x7JVJ
kApEElpSRKwUCMZ3Pku5y+i9bW3SU3VQsdicuH4+d9mp2/pi0gR1jrXWh3w1640yUDzRuE52wckz
Yei03OtzISda2VKuNiSW15G34xLb55X5YFBhckr5FTZ68h6ZQW36ME4VnVi/KUigUDuXBFNrH1Ks
npXoIVXP/ft4ELg35KhUORJgJiyVzg2QF99Kxezrf82nyVmhwBmm4u2oADBMdN8X2cSPDwA38h8M
44P6qrE7O5BYofC89uIl52vQYtTaP6KBTmFQXjv96F4c67jDeFLrI4FWnMu+uAB5lKZcjQOStdgn
dbKC7OH98jZq8sZ9PezPOysHzcg7l5AZ/nF5iTh9bvYmZVGxtEpcmLBak7uLtdjNwN/fjta6KmB4
317dATJOnAlJJKVkaU94HoSCLxpypqnIFzFoojZAjU+Z6P0kMoiP3qJKf1U3Xf3PMLBfUPjPj6vh
lDZ5wBCe2oZHywxZJU70L/K2ZlH9U+Iq9w/Xoblqe0qwStFOVTYVD48d234rtg5zD/xAbpCtljzL
MZDIq0EJltnbNQJROFMuYyoae4fHjuqQvArVTr1n6GoOCxWQSSO2eYw3GEig7mt9A+6jcDy3Hgty
p9aP0qwUAdQEoWk9JYChczmsTapgWLe9fPmZv9Bq1owecHLGRB4627dAyn2iS9tZ/UONo5Abv88o
0gKfS7mhZuOkrJzIhOsOdeywPFxS8eDw4seZbaHgo7G2Herpkkr5gNafz07pbzfXSCsgZ4MBKv1s
2paQ1m3cIEvj1tjLNOHvVlYHFdsRzaAh5urKBShRR2VJlqYUlF8GgNiU9qlZck0Yt/uZ26U+kjbz
LKb+jYx1fwfr9ZCu4OSfTt6NwCEKswRo/mIE3ZHADsf6fTvvyTY+gTcPH6y6yE/RMR02gv4UQD/E
q6Qwskr9ZgLvWN0x/tMXPV/WYK/yLJpx/7yUHLiQu1Xazk4/nb68mdaAo828YzQJXDlZLgRpmmVn
vgRd2MklvMnbGafF2HjNo2ybtamHLU18HuFSRTF3gunkIGoqu3CYL6Jit0p1eRn+rq+yEJkLcRTC
gpZhYKz33KtqrbrX9hUvaF/CvwyvhhJBqQu6XtB7xuDVX9te/VJ9IANHa0jzPSygBT0ZNeNF5U7y
yBRLgOXj0CE7W3CQ/PJVXkwtdy31MeMgggoI8vIBus7/AeoJAYQr5sr7EBYjbdnIzCI8NzZNCHCe
pkCWU+gjPZmghWzg8jhnS8qiZOII2zGfn7xbwGXV7rdOehup7i+BxnCnubOBu+gKJGXw+yQo5tnS
8gEI7TuLiZm1rUmwuHW4UYNB0J7VLXF2KgR7hAi64jMp4vks/fCozLYJEUV4fRHVTpSz/44gO4nB
c6dvRfePmHokKKyouu2zinHX332B7SXRteq4YSXvxITARDbiHib0R76E3+QpinGWqTq1ZX2q5yn3
UegxFZP71NxEc1Xb9uAN2tC/kyAyGwhEts0PTd8vZHnP0OSA6NtnH/qvVnp32Iy/TaC6yeGwhtQs
cIQfN6uRj7y3lE8BzhPRoaVdX4tT0D7aXaFZ34rRocdLPY9LhwkF2YFmJYeqN/vonyL6edQ8EWOy
d9Heg8VtC6NLrht/2+1g4G3heWFUI12GxI+glIF5V2EUTjkiu2DcQDnMLVqEY1LqVHPoVz3PhGVZ
KQTkI60+OhkTrdeab3wMShDi8SYCv0U64wnbGbfTaPm+2r6TEORITc0Rs2ZkZGS5SoKl5EDIxiDX
V5sg2w510xKIgWdHjkBzq5bMcr4+UxI5m8o/9QL39l2N2pKrjRsyg12/k8ppaHPGh7kYQ+1VhzVI
81SnVA6xD/H7h86UN7RNzs0iCC1RbuHslKQXWc8x/+n0x4bg5PaIAXQX/CO744guaepyNQ2xRMQ1
ETDaPZgUl+N6/IDcCMtuYvO1MiuvscvOop8BYLLNFYVsGnMxBtceJr6tFPzqSwCezAdNQdqdM718
Q+/uwqg5I0VHJITo7AlO9r+WtvgkphJECRjr49vZQ72XjhkFULsKeq0K3dKlGaiZd8GvbEBtdKXf
1hWS2M/pDuodSdweN7blVQVUpXci6W6DSz6AeQN6Ooy3RMsdvm3cSu3GdJHbFqtkWc0jdVfDY4na
fKhM/YVwbId3yMycdly3Cu4w63enmdUNFm9zdoYA25yCxOJn23GK8Mi6XFf6h2NSVqrPYyYtI318
JpjSHuEoVRlS7Y6fcZe8SOzFeo66QOs1BHUAeoCGmBs8ihb6oPxXrezS8hgKW3CHIn1uCSswUvCV
0QVVPbWXCYLvF7HKpM5v7Cups8SygneO4nhla9DW9iSPEvyrai0seXl7Kyyg7QBLBx5Puu7p7Hez
sVBeZVIXTcBk2teVrzSmshnRRXTT/lVNORq1dngRbLAoE5yYXEZW6l03MxbiD+KEz847kLNz1ji3
vLliWhFv+zaCsdlJn0zBu6NDDqwDlKfRq9Lm7l9bj9+a911qu04IaMgsCGd4ywGu/a5ONe0Cys4I
8BrstNutqzc8QYvWNvFaGLANMj9w1095g2AF68nN0RMdcylWawV1oYfHwkWE2wu4D2VdRZiFnvLe
2usYtYLHGVglulZImABn4zFZr7/viVXvgF8F81Cx/eejLj7FwBYjLFKj0QWnjtcDZKCDJlbQwnTH
ANFcD7Dbu7n+8xIHBSgwYS0hhwDTSQhO/7PBXKOmFRTxzSKWYi+p+Yy8UEFzT1R7mOGw75Fpydoj
kacGjcUAYoWrzHhVxhTVS/fOBnuXMdMGedp3zleaof5e0/RsiYIQafInTt1n166EC8/srbwXGV8T
OOE6MVrhXhPUfEBgn1+JAGVztRaeZ6pbebXePyQlNAaJFBICjF9qGoBfLPX9JrGRbBiBmzBD9JsD
9mU5r0TgtzgVzyLgVELoYQ/dB4jywZ1heEDzkjjl0Rjbrs3ryMPh505B6mdQZgrddfynwUPQsNZu
ACetBaH3R2cwhk7x5Sfq6slj2dCsWZ0Nnc8BogECxzlJP4YOj22J9LMXDO5Os5YWmx4aNbVQYoKA
q+i4EWSUuj3UGnl2qsQuC+tDRfU7zFgSJxtdr16M4kXXh1FsxVBPoUkdT7pzpxqSsXcahOHkV2EC
/ZJHdPG4SIDEPwoE1P1t5gRiA9AQLJsC992hYLMAqU8Wrd43z0OEj2gpgt/UcOROKpOmPkJcyv5r
OO9+6e+vQ5Nvk5MrD6JhXDLktwMgbxRbGLjAO+Ru3AR5S5E7wkpht+EAREx5dynLuId6nos5g8YP
eDQV5xBn7gg4+pSLzlIoGlf08v/EWB8ikoVVKDHbvta7HR6Nx33Ep+8vJmH9UedMB3LcsqzeIBx+
Z0fM3638cTZjXKLyCqwtbhUT5bq91CwWw/rgduVzORHNtwEFHHEH0r8vf5g5zIXxt1I7zYP5c3+b
9yaJZtHXuxV8sRl9I5vx1VlotqYM/v+IjLtGZQpBHf57aShdtPU1M11h6L+oycPKTG/+bruu0kCF
ovC/EPte2CaM4x3rVFds2oOXSp311n5TDL2pp/2Nv5XPUEpqEdEJUU3vHMKruK9GB9FwtNGQspoq
9641QwcWlv3ntqYVAEQ1WImUii8swq8VW1WjBV+po9ns9NdFMPmb7EwHZT3Ip0fvNaz/KHP4hFb2
UrpDoYrYqijk11GBItd5CMF4h//mpRctHuJAM8hkoBbJUoWRCk4oMAU7dKWEqCLGMbHPMWVlSIZI
djRLDu4XPTyrED3Vwgxc6ekTW7C6v47/aCcBsSPUgXJb30hmUHU+eogHM/eBbkUZG/urOAH86FsT
DRd1wQAb/Q5Nx5Z2svkyi8ufjXsJceF3knjmBwsrlHzFKV5hdFDBx9H+JK9C6hoY2pnBAv38x+MM
I/BnkalqWejhUvgucrfxjpfLKxj8UH5Qe41pWVMOUVivw4gRMS9SnZ155NqppadrwYdaaA/9Xcxn
MhvSCLdgBv5fkuJ7FiMVghnkbn1AWzdd5+95i2zQiHwDQkKXpE1xz8/AsWzeaHLAdt6wvTyyAmKv
VtmVHYqQgU3dL2LCtXss3HjizsKgNTE9ia9cHUsyzBdExdsTPuthWjO6DAKfQ6Zmr6yrhR2VMuPB
Sn9rlFvNcsCU3itYBnCxYFDDcuQ464Pohsd2FoVs4z6PssxqJHEwk2IIYwq3U7OgJ2/WHzI2FGnK
hm4fV25zZrvGmiheEgcWt0KMNfN/WcLWo3rzWCV4b+/WNzDa0FCc5d7md/GDaEfX9+7Sz+dhccfI
FTje3ch7Wdr8TiOEhsH7wLLo1/9Qe7JgYqrVqKHi1OxT9F8WplgYnmROTcRn/QLUozjaNBOE0XfY
koEDN8GIVkcn4+wn23X4gKNaLfhmto4hrcXv6eAz3A2e5eaSNv1AII2pbl5fKd0TZnH/6LSNYCkR
O53z43mhkZseUNSEz136mIZG22mPReeUCRPcbgopeHxa2NQPLDFVJdQ+qe3kXhS+vU/z1TWQ5g/P
1FzUtGCSFzr7PTFEXXel3iekE70UlSyxnqGlQD8Naq1tLxVZ0q4O7tazrynipG9pIqiKdOiZ0lRf
sMZyJJGkBBeMuDs9p2rrNnNZRMHvpqRV2CO+NONo9j4KN6JR1KcXFF4WaDYo67X6Hqz060sY392B
tPHzg4BVdBmtVLaPx/2U7LLzJxh+pnLBpCLWieGzIjh+ztHDa2MsOclf52Lzx5DOwGRbKcpGkxRA
8NhRWO6Q1V910/ZZ6GHu0RCOa5qXQ7foakwk4zAYfXW9UwZ9L5wtJfgrQp9gInvj2LeXQPlD0ZWr
2mrs7cNCtPQIjLMFQMUipuq3vudFPWDI9kvA8p/ocajG/qL+D6Ikvk3rTHC2aEX+Y9HD58uNUAyb
EoHGzX5wupaeI88vLzyb9fC6tz+RSKKpwWQj568j4/SAmzNqut/6LdiPZkhjj16+p/uyFz+G85EI
X/V6qWVCaWUTFskNTy59Q52BxcUxHWNXuZZAvJ+h8Ro+1e3XBQUUCro95HpZhA4VnMChmfuG89Pw
6o3VWp0ybQhLOOrjWmZEurPU1Uf1kXXbeQ9ixyW3KCVt6pfSKwqE97TpoIOb1S2cG+GG96bweh/8
qMZQq0JcTBTSgBNVgDdSag+/mpwwJp9nqCkGDNktMm/Iil0zZPAYPUzZ23racZcwTXQGNf5JgCOy
INZudfRLtnIK2/yPcfBb+vzVcNGrYrKCiH6LVj819T9Zkx5wT2ULLfmub9ctVJjxUkMCk6LzZ9PL
C1/DOdnDgsEcld67aJg6fpc3I5j5aM5WxUegiQBXO1FVDJZ1KcP+ubCvZrc7dWF3sAH1S1EvGabV
zjbPLkGjMdxtktk6wduJBrZRYOsMVQRdNj6Jp126Oa1zqhpoh6JxL/jpNVvsr7M6mWroxcw9Tk5U
lAaT2CCb3SHaxm1VwfboEPjfVavOxp8zweJ91X7A77JmO3bciaksYqqIvKJtfzuQUh+0qh5Ihqxn
tol36t0naFRMKYZbGiaHsz+PrMXcRgKaxljHKeAHMedARFRKF9kkSyWDt6mycieqVATObFk0t8sZ
Fwr0DHchAnVgvKJRrNu6IlahrPZ/0YZXExIBoQ2wJi9/AzJ8a6jo1IBoEWPMGIE649w/SeXcC0eY
LL8nv4M2qZ5iCMR09oPIEHNTyKx5tkfD0y+0jOHLW7QamZQ7gSbkxuyxr6Pw5IRZKV99yu6bABXj
+HQkxOoFkWji8ya1wNwl6Dixp5ymYf7l4xMG2Dv1MgKyz5bXbntUZGTtyRxsfo6vR4nejYJSl6RP
o98zde5+5f65bd/fZFmlZ9l8Rqlp1OPWyHvPfz+4vzg+klPee7l5FzbV4rEP8GmyqhWCMfJ28+s9
c15XnZDO+xNO7/GW4gCbrOI0LmzoNYpe2RSF7XfrZksnC1Rkhy8foHSLJz36LOUeG5EV38LLt9Pz
YL05MR++utL43/2A47VStyf2WNO+WJ/Go+g2LiGI8vCJOOhgkTW5oNYIJglZH2DcsuS6Yg7P3IkP
ly9GPuCWaB/4nB7j3S2DyK1xzHdIInvOv2ALgJQ/9iO1RHbZyyS2WPLb9FytD04wJQuhr9XT7OvN
0TgREiN9fLZJYiWmqksUrTW7RRu6uhZlqT0E8sMYotSq+CoSTRaew3dlaiu1g8TuyZ3XR0Tw8WSR
sg4krgRarZNU1NCbO694pjMgR+2A/jERy2hDbbc/9isPiSlFH/9QvZOrXg5lWY8qJShxsBKAXxjW
du3erY25NrDoFUUn7XH7po18j/yH213fPGzdeCBXeOA1kHLrkZN+KJj5lHJDqordho1/PeTqrPsB
5QfER71zK0iNzyC60HtObQoqqYu8h+LKuHO/pCFxtBnF35wH1ZuTBX3sbxstZ6TBcZkDZ3vMRxNI
lAjA6j7aqss1I5STMmuwR0RtPzAQpk1oz3z23QoV1CfUwR1mgdUukZCjfAkp9xJSGwLMzR5H837O
UKR/Q5LLXA4XCpEywlVW7zYRtFk0oB5nzBwU3iG1YfFMpyGkHcYj2aYroE9RVJQNF9YLTs4x5eEy
LLRnxnmU4ph6FIcB/ylMn5RU7glKe5m0ZUgllthAy9S+gfB+PhHkxUoG219zp4yN0ZU8zLlfGmPg
xf6sDWVAJIi2JehYIeI0G8LmRoiEU5HFEuggoPPmP/OaoP2lDQSAMYGY2rB2cjsYLxnYAQElTR3A
pxi9pR+jSpBP0FyYGX/CtVs1G+0Qzcjt0lNikkhLyhjfubI4g8MW//ZJE4aruLTGurnpc84s7zti
nWf8EPe2dKbAJ4q40Iqjk+B348OPduZFtBKzE/nPSmsS6uNJuUjsHnV3RqUOp4uMmhUNnK2CgCBl
ArbAIZrUQXt8i56eh24gR88qD27NpEM9FiwPV9cY6jeiCuca+fGPxYDlJavC/7CTL+1IQNpmJ4pM
YzoqSTyNt3cU/535fRi2RFerGNWh0UFbL/XpH49M3skvd31bSTsUeoykNdF4YyjdnB8XXhGTt1n1
Upm/a5u54dhTvy3Ds3yYgzb5PS/9wUrM4g3HwbwSF6aHETiD5QvtOq4oDQCN6AZ37Y271qeH9IUj
CnGshyqriS7AYUiZRRZm1IAt4TpoeAShQmbFiQRcxRUlMUuQROzLi06VmgLkwcaAk4oRegsk2sNJ
QIlN4iWcAZaTyaobUfCG8p8Q5G85UYtvQMIMHIp860VxVm3jyukEq22tNjWDdvv35n862qgA/cTD
WgztqARF92Xy9abmOkbZ/1G0Vh8Aqfh1jL0vIWT1U1DLDx1r/2c5Ep1cxwkgQ7ZQ7I6HyecTCO/B
zbLMkE9oMF/z/rt78wkrq3cu/2weVIh/WhJ4KN3DvArr8wEMmKILvRABIZOTAgzk5z8LaQj0gCBA
LGa7sD9/AdJuAPvbG30sD8HE3vDMYbrVe5JGmyReCbazmH3MRBkj5LTXygRixlWm3sB63I0AV/D1
doJG/dGqEK4AcB5JveZ+/2Fz55WoHT0AA6KfLCfbfd3N5obtbdUpu2j9EUj+965DXiFaAbuoeJ9T
M+Yxjz/0fVmqGFgHpCTfubt7ka9fTqgMF83YLPM1pbGD8AjLCSz25JuqKFKveVGUIxvCCmaSH3yy
aESPrLRqatqVHLaBxBUr1Wv5lHdSQ44rLFlw08Vm+p4mahymQvCZQyn0d2DoJ3i7tN0XaBYlxBII
i+5zGLASIutiMf503oaOqvx2vzKiTVLiHfDBn9uKdNwrjolwv+XawPFdmOa8qtC8y9ihxVZkfony
o64NCYhGPIj/jH7WGvFTBka4WajzTYEIT2HWN9yc998saIqJR2sYQDYMv8Y8/WvJSMcczWkcUjBv
zUxB0+EPGjZFv5FUfkxgcX6vfTQe28KTOy0+JsPX9KE6uaHvW3cTR2SbAhxMCsU5wUpbWyGBwijD
dDwm0MXNmkEkfwYesUfbId1xA1aRs9LRMK6O6y6ToU8CG3CEl2gEek44e0jH552Lw6nkK5TiMZ9W
glctWr5qgx8l8UTH1T4u6dhnPsOt1Eh43r9nKZIlKhifUSggnbWDSkuZfjmF7WXNmOEy0k54vpr5
fEBnyOIYXSJnzogHdUblnILyZWx0SoKYS+AWCcwcaoOzN7bOsz4m7inYz0gX+VFNMYg+gSepaZ/A
ICgJeFBuvs2htNMs8r1ZPgR7RhUqEOIoVW8wUmL1Y1TzbyCGQ2mgMTN+QtqElB8S05FcHF5Gtvsb
/T6VW2rtxP43drVb0vorFZ4yeO2B7G6AtL51Q50fnNtwk8BlXsxrf5n9i7Cd7sBO5uwtzTQAcHr3
OuGVaFd/vjXbBSJrvqBPKg3iQ2IRuVrqoLhMcyzwJE/53NfodB18/H2TY6f9MmO73VaWRQXqMyho
N3Kw5oiUtLHR714WDYQYLVtZhbE6eNkg6OqrX6ZevedEfd6U5z8pYr+Wgnhh2gcEZjWZHSOFdEwp
IttnP+stRPmqutwgHSYsVeKCUCAW/JrfCtnyqUQm37vRLU1kvIJBfSKAxv6nY2s/C9Tjdlnmrz0w
6ff89dVnQL63+PfysfLBvjxLVmeLX+J3oYicsRO0kp5ajdMDPvbViCtJ6yxcTnjfwTG1M1GYFs90
M0b6TGTkPIZ69HC3j1xBDeoDv4jE018qIohHF3Pix7VYEx6WvDjo57dP1LXMd+EEKUQa7p1SS8dQ
iU0y6W2dODFF1ITDozsM6BXzSvkqd3ZO/J3xNcaVAKrbmFYisvQTvmgNlru94o5/g9Tcm8Zo8JNS
Zs6zn4jFD66Sx92K7j+E2S4Cwmljw7TcfGkD/BuomoRhEoochuxqbn070UpAx/MWYAX+qg4BjJ9a
wP4QCLdeutcujLPHSpD5wx0Rcq1/eqz9AczMqKsIPtznx8nkjbcslqjJodf3nrJhxebNJ3f2osQ0
YcnxnHkkzrS7vUpNVwbCXofun5rxpRrNQgffOvoBjFNaWNiipcnCGYAmsRhhsw1+NAJNEqMtkxTj
FKVjdbuqJJthE4YSDg57BQIeUPm/ECttvpraVEj+EVbemZxpK3GVdcswqsGUQlu3XwfQiGvqQHfG
knIM5NbDjNNE5j7V02XZHDhLBBdX8qAoCGyTmgYOLbBKL/Ji3HOMmF4XSe5tig6zqGvMAvQxbi33
1w1Kvm57HQQLuT9MK5xRlCF6QteZWnamHOUkx2Zu7u5Uy6SNUfWU912WlZ0HD70MwEQA0KWWubWb
F+fl4aMSPyM9+hL9gz09rBpU+uqmgsD5MxD77ToMbnZzv7qK7/MQMOFI8aYFcobLz3/9CfLvc87T
vS0cIQLR+7I6WOD/RONQebUdz8V6ksrIYUu4yGwNp1XI5+GIsyay3P7MqeB0Ai/iQCmoZQlJvhKH
PpBBkZAzLSTEaI7iKtKbSJcuHt+h7o+Yu1uNUSg3mmxulI4rIaNaQlmDrG6dm+MPmyTRvGJwzsks
nb9mqyMbmPsbX+8S8fJALj/vgq4kMkD8DE9tR+XC8TErpv0P0YlVBgIqJsLzVGPqXb6nmvFjHCnI
gpV1HeZCAyVPi7yvTc1roAFNINOgzWaPfcK7Cr+bxg7mcg1FmLVOqsv5rsVP/Bq2+RiBRawHz4x4
RjVQ5rk2Eb7SI1OzMZ0hPqJoClUzMr/UzpRNR4hbtEktN9bRYedIT46y6UXvGWX6d4lSKaJkxixw
7IwlAcYgXOOIWnAE/eCG9kwX2iiDfvdnxnmVt8y8XRayV17bGTGxSzIzzxXWGfAUsr9MoF3GfeI7
TC0jZAFr9dRkgKJj659ShbTSMOUzdg6arBtwFIUAgJNYLz7SY1ZluwvDSXGbxLQRVkIecC5VpKHB
ktDlTywucvMs7WmopXBi7IDAD1n1a4zhPJr4N+ELQQxwaFDVAlvjGNDF1oXdZgXGALmfLpsRoynp
Nnqd5xYxOfijiFOHIBPhIKAxYw1O2zfLXSqpg7yx+Agiv6KpZ/zWF/e7x3F5/Ps5EXhhmUsdILNF
N8qlxOVwKhcVQfPYBQTHeVh2WGeSpB3ctmeq8hi71vh6RgwLyE8X7Y9WgcRfkUX+fo4lNaFQLSs9
wnT9wNKJJpkl3LgYFz5K7OpnhChEebBE6aMSsDhJe7/sUNNdfUKQs4oi9+T6pyqETFkmaoPRr+6N
TSvF52eZqoIhWFip3A2repr95hi8BOPeaQimUMNowPf4xAqSOuL1V8boyoevxmTUL1y4pFAlW88t
9a2BE4uOVBycx3aX+LaPT/eSeYZctPd5hLKmHpEPW07GNkQ8cMjZgCGBlrwSY1rMIisVh90m8D98
8pGbDamFirIgzT8GwwSOcZz08ks6O9AvGXEh7UEn2V37x1dgXUgf7sZAFp0cWfZ/Pw6D4Jm/selC
urN+piIcuW6laRjM+LzYqMMmEtoD4vcRBwi8z/sqHR4IfIkBfffGDQt/rL0S2YgpkDO9af2gvQxZ
ENyPqov1iYH4CObMdnOJs7ls+JjBIfb4GpakTKhCX3VWvtvNRfP47d7JNq/sd3vSQOoo4dXLKYY9
5ZCJvb7efOcYgDkHpaA67HrQTciQgHHg7B9g9BiYRAH2en1ChQtCeuHHadM1wHJzro7QO1up8IS8
De15plNU/KltJLS3+Wof23ocunTZr0CtrkU8xJgUIZmxufF2xZF6xBl8u2DgH/McICYOaLl5fYix
/xZ0pYiJ8MyfoD3ThkJVXDdpgpJ2DBshcfv1Fjx3iXWbk5yDzGccfNPjH6HDwoYbCmae9XGFh3EW
MxlbvyTTNGvSHav3Z4n0v9iHecB058Fx8iEeLy1VNGHOHfNT7If0zR4UoHFeca0IOqJ0anrrQ71R
5nKB/hZebSKFWpowbjkRZtjFI8p5G+SH9vkfqBSztyITg4RaLCC5eKnLVElTkitVRTbK4wmZAe7K
zcjtEKs3Z2+ywzrBm5vdgLlaPqhCQssmcYTEdFo3b2kLo9nHQclF3J7GB0IGbz2NmA4PoOYtxZxA
2g27uMh9rHipfGxwB8FpQWKVUSVg1nfapPyK3wMv1COluKMFudHI+n9QI7kCqruKuRKqzTGSAOQ5
hXoYL3M6bT7UwS4KfMlDwKxTK6dFlM1L3cOiXQ6pxL7OaXS7CDlGuj7CMUw9ydTBs+Q2KrPkzmpc
4zDvXvG9Nmptc7DVUvurufLcOgVtQdhJklT7RDI8gyaNcv+dDAKWH4DtCwfgaaJjDNCBvrCxWtKx
LyeR/Upfb0TqA+JyLGGkJ/vc1Yutg+MQDJREcnnRIkNpNK+EdZk3Qzzm8ndrKcZvmLqqMRbQAgFS
0VPdcrdjddU+bPS0UUiHV8s6Qvrd663EXuItdNEsmLbXXtedFoDqCZHvvmv8+POTcSBfnaqAcvTz
0LGtwySUDLfOhFGAj4F72liZ0cISE5c4Jmw8uyii39CjAeCcencwRrC+NcddjO08sfb/BF1jr5oj
uK4joXWIlF8k/e5JhuT0uSWZDqE/dsP1Iz/U2NfpTskd6D2DNluvs6tmKQtn2/BH3p41mxXn/Dvx
FvYzxAYk/LtPJxoR+CZbfyiDn+hvrkfEWAsmztdjpVl2Z0upG81BdUnv71/5kFLOvD3Oh6cPtKxX
FV7Kk2hlUatTOKXjdOgSA26g0g1Q/MrHJEfkDaIumGXdPuGTgC06wMxgYD4Py5Fk3kPT4p7OhjFx
y0GVC0QmyibKFAazEbCBuuUYN/n2KWAjTIEDpu9gWcxGfJpl4ZS7kISE3zF5RyWRqSYE1gEPy5Qz
Sa+dwaXU/zs0uca1boVUx3cHSKJK2q4Y70HV/nvhMSfxb35sFFZ5nmkD5XPAatXw5Gg5/Vyti9uE
JwkwsrZ1nFMJwGPHClF2Lq5BO6kGboI1HRPH83La4NF+v39WxRVKO4vEd3GitPjq/wVZ1LN/t2qi
sTp6lrE+9ad3YslV3bi+Hgk0PvrULlUdfmQ5QazwLKY2tgIA8CpfXzEQYxuMyHNHu49qStvSFE7n
B3tZtL+JUf4lseBRmnXaNIBRueOgS7q/uEb4uAdW6x9o0JLhFctM14E8f36geCjXJVKGyVwWFAUa
ur7/Z0JF0qk2NLB2Bi2/dTmN/RQh6Y6HwmYray4spXSIf0z2BApWzsqWXFd33PZ56h3TAzcfvn0r
EPMd+MppMY7Ppgn7jCTeP7RNna6MgzkwdbWe7iXRh8TxYjYJOTWSiX5RDrYCk/VOaRgHBU9jQSDX
Hv/1mr4yhNIN7k7pPoJszhLW/PVnVjWwrXC25wcfeJgsmVTTQe/zdEBtTK+lYCaPLLNcJPBhCwXn
QUBFkmHRw4nS4cdQLrYQ+oYJVctuAb+e4B43NrJAmYWySCOrU8T3G37WuS+zZk9ZI3dIzWoXfYoZ
Y1laLp8RCVCKICZ9HZR5AqaN7xRuXScixz56nQmMG6Oh5Rh+oK6hImFyF0802BizlFdDSpWOYfbI
ZctA6cNOp81xiZKmi7BKl1knq2pDyah0DGXVILqeGE2S286CX8zcux5En6hNHkI5PplJDbdwDAst
ri+jn68+piUyCAHFvPLqUCzUQOFL2G5Y0kofDCcULpLMCl3lQTd/eWCx/2SORcB5TUrbTWsu6H9U
Xgo50zgoIe5+bbU7caSUM7hBUffWasRoQinAwfz0jfcRa2ZyPjRFD9FPQXJPZDgmQIFvytrzixy2
XnQGdx05qCaCE2/Up23ezbtQ1SnkcatdxoXZRPuFTfUzksPMNgx9ssFXFIFAHy47HMt61H6Ia0G9
7can3Z/izW7gVp+NEdo0TPKOwB4f4ucs6Y5nyW/wuDCDLbJJNPqj+QC+IwRGNQ7xPlj8y+fPiwur
wzKI0rW0RmCTC89plrZXQt1+RbXiXAOprq/Bo6ietTXzTqcHQQJCNoKM2kAEAKVGXy7L1A2mrCQo
TE4CF6X3SVUunL6/6tFayXzu/BBdGxafZ4wUH5i73TMcQKnHqtRphKVob1nB1O2+HP1NU69c+W6t
aVYxQYVAAapWpzuZ4QyzJ0sKDCOojGM653BT8621Fl4n+Kvrd5b+ZjDiWk9T6HRDryAbUFQCmWNL
YXJOQT/kx690OJWu7KWm5jVtUoyz/t53fDpt1TLBJU0NniVVtb06rtfSNzHcZsKT+Loyv9XBpWxf
lpuGFtTbvDX4Sgu5wrLYnzQR99o1nIzPpaUelLbwef1MUB6ysDjAqvS8iYm7LpVspBvSaNSH+wfD
YuKJLk3n+zePkJYtsNV6nwm/Jvyf5eLtTYtw2J9qL1WORp+oVAkbClEskxCO4btspjhT6chpl4Ug
jTrVd3zgzLEjjJ/Zb5LcCGAstnPlBY1jJfUXsAARzFxgTIcmM0su4Mu0ZFozRnLaK4GvYuKwl54f
MHTb7JwuwC1X3L+j/cMpw1uD000bmAvgozi7+le5xJu67viK3fCr9IuCgYJKrQp4lbywJk8usXj3
wMK1hgZ72+Qx6fOsRHluaZsBWpJbF+ztGmXGpK9fTVdumpoPfsX6FMz1Nglrz7IKb7PTIw/qphyG
7RLFrd5t+XidFj7QTi+JPDVM8ssKoj1eD3X3dymSNJXsjNoc+37Hwr8sEpOx8qh4zg0wE45FBHQi
/rn2xkX1YHWCzHuejHeN+OGoJSdyOgT+0WQR5XSBuQUSRo+/o0yAG3IFOtokVmDCRZz0sfZESbqi
DEZqyj5Hz81jzCtNqvlEyMeBp1AQs6/nGPa5YBgXE2VXyHy3uLllqLz15yi5E3rDizIYqbXp/Nvu
h9AnsudVviBktP1XgvUV8+0OVmYFkAVrIOj1kuWvInlbejAtvHVRCFiLUAIZ2UedIoZEb+jvtbrt
Y2J2Pl65ChBsMFaE0zL/Roxmpfzw49sijdGAQrB11dnYzWJd8YeZJH/S+ik8ai6UkZiM1+yNmX27
T5i7KqnCbZSAvVPU/5j/TwPtsLF7Yv0HWTL3JXQrin6xx4/xVhs2Pt2T/SU4OStpYEHuawffwOAm
64ap/btk5DSz1CO/bUZKaFFNt0ddls58q6seRIeHYBzZl0Xb7Wx+/OsvJ1i5rosr1AdhYwUuG3OU
56Np5I9ZlBG6pgypVptWzrVQdgQRJVQtQbFBnSw4c9IkrAt3d7rwr0TnFRYjPvqHKQYXcad+2+AW
Pz/LvkEH2toHLkP7bMa//HS2EQELyd2yTE96R4uRl2G4S0osahdijvr3fiiw7xdP+Gr6qr2m85V8
mYY2XVTjH1990rGiM2nxYg0T0z8/+IwpIbwH3cXtpeF0jaU9K8+mnrBk3wOlSywCaShc+DE/1sbn
F79gWm9yBJsSdMUP6wx6qcclLmEEJpKXvdL+EsmlH/Mtgzwz+6gPftd0nGh+uoTVbJBLs52Agd4P
Q4FBJcpanabrIWFMvWEygkmWrfwOKT/uUXMw39pGWe4pL/H4FF4EofcM/au08rC0aJ1w05gYMVxA
L/Gp6nFplIMryx/ADdfnEPeXtAsBr5nDbGDX/clLNaSiKwJ6CPsX1XlMexd0QbIddIGEUKM0dAKT
xD2x+HwwKMISM9dvrJOlL1meF7H5LrxsIch8MLOB5ig0KHE13djVL1H9O5rZdfTb4rl9l4T4MXWu
Jw5A54pwVA3NLABioB9irLzUq41ZLDkfW+qVPo7wQ4m5/BMXuC0dPEtCGcgivq6KDeSApfllVau3
YEAyDLP0uKBMwopcZpzoTzKozw1qP1+VqNLDZd8JlrwWZf3zpgbsTvQbRftTJxKJYZYUhMLP26ko
jykNr49RS+LbYPDrD4TLOmv8bVKqkpzBTxalqWaxcbVrVardUj6DU0JPVU4lCbVaqqEj8MONM/Po
ERK75hyoJkPKxo31cuk2GBDKceCPlzhStHuY3zqz35EXcKU15Bm2VvhAdfGZ12qZTDCiGu8ooMhl
UV+k68sXhaIAABsRJ/nJ3WQWyi8YpOs3RgD4O+26ItBT+BIEGt8DwOJi7IMTLo1u+S7mWVkfJYgu
3x6wR7urE6bQYkG8+MUC6wE/0+pNz6blvt5W6b4zi8XX2CMvvwapiAxpmcbErBU6ZzmzKi5KwE/Q
OL1AY8fiLoPLVK6+8EI5q/6++SA/qAYXJ1cpQ3jXe1++hSRcFV+y7nuhdzJmktjt3h6iIcsvokTw
c1HDjhAM4IzHgJxynN9VxJiV85C/6TaZeqVFPIAxWbey39JSA4g76doacuQ2LHeOxzItjaRgB4aK
bQGdAGG6Du1SrCPNRrYflQJmE20xNTFlymJ/CvwIg9DyZS6uxjl4U2lIp+uVSasHV6RVd/Lzvpyb
5RNzVlZSoDF8hb7M+cLExPU/s3BrOUQVZL801UhhbBtB7apDxcGGcUkBz2rKBsXEp/bnQpTkJ8Gj
92dbVCu8vDDJ8vT4E3zX0jHV5JBPQdK7RYzTh1sL0vX/fVKpoY7SxKkJwsNLkpe7kBYLr4Z+I0oP
/2brMDtXj/FBOmuHaBgUxN3JFdhbQHM1aE+mSK3KsI4W32hY9VRxymARpKgYM6fV2ruhK88dJfZE
NJYoZUqXkFMp/Lv6he4IsElJCrT0R2lEsGa/1jt3eKao//RCDf9lz0nf4L+VLHlrW1zU72i7EKjv
2Z4XRVAOnrvKKvlp1J8fB47mjnCZIII8E/aHr4iqt5LGdJWhvzNaF3PFr4vLXIrQQVZDDZOReo/h
CYvXW24ZkC+62YIGyGa9vhq5UUaoqYaS+FwjMHzxvaeUyoT4MjubWbqDW3WaMmVOlMH5NQTgmDfG
e2wLrdZhiTfGNFKR2cZWIF/vtkHIuxJt4oJFkEkhkF0hwGuGQGXk2mWu7pQTEdoUzW3o/D+vwWnw
yK6pWSfPS5itRYFnlVpjr4vGsgEv+bf07Rx0VsF3X/QnQshHvFuSnC8ctdgtrprssUCwjJ7hjaZ0
nHJT0jygnEkrywCQXDXXHSAHV0TwijrGoPbqkI0VePSeWp1EAm0/XWcotMVKDopzrYNHVV6SJUHn
OEjQ18tFNk7WzTViPo3lzi41Kf3vHoVdkeNvxAHO0DR9fsucZzdhh/86OZjQ33aaW+gaD2YMDvcp
LFOEWPl5vpjM/s0iN8Q+QJesmT+zIkwJBu7sJ9+sQq3LNq6qc7bDT70Kvo3+1Tu+feSNCiiBB5Nf
YHhUNnrsSbKJS/1frnhu9uqbyrv9CXL2+SKf0Xvtm+1b8S4KoIiJ2egQbxt+B3DmOkO0qyY6B+k1
b5irGmZZotpVVqMvyAswbp/1OSoYlRa0/WCOcepBHcAyKJOmxv2C810q1miqIclOXjRry2v8VHYP
821f8WGXgO7K8Wpk9iLsSafxrs0lVlhgM1PQG4DM6zk/k4cI1uZhKKQpSyrcG4IYEvu9bc9p0BGS
wNFHSUoSejJKfGVLDBQ1E1ARLibn2VY+zzizGW9OrjKBqP9bHwFLbnlYm7RCiCgp7O6f1nHURB0D
NiZCCfWyGS8BGIzhS88fFLbKPsJ9eNt39MkvJ4IJUXV9stI0iYRejjTjEgVMi1KW0kTjA+FI6wG+
cCJwMSxRq7d5xoyOmmrw8Rt5yRaIb/Wqu/1sxDeTHPzfdtV8pdTrynPX1QSBuP7NnD6cyT7pTa9K
h6jsaPLePkxnMWP0OqAjuqtF86mJX/gpAOj68fXuPhCS6H+Ldwh8kBNt1AtOCXZVg+kt+yUT2CkD
9+p4Y10YsFSoQPQNBxnkHhJPwCLcS53emM1U+ko+wVTzK2P3da2X7t4LObm5v4D+M5ZZcyHOjHq+
AnXZlqxdIKAN9aAKzFEH20c+X7oMq5Gry1jBmaBG9deBu9eWJ/Gl9fECiUq5olE6hJebguw0Oa/Q
bG1M5TYIYQdBMgQuaKih34PyhCzJ/Pgd1mpCkP3qEitRJS6Sx7YZ8/Rxa+ItwKZu006kNPZ6dplJ
HeGhpBZGNJ1Afc8LMMWLCoQ+KHK711QQWtpQzgRAT6bbGl+bua9yzBqM2rJ4GDxCAjYXg6aEtlcL
YmqPguq5CEzMqu5fTJkh2rYJgJJtaMM2epe3nxawCpsmJ+PJHM4T60kkNBYtxfvYxDk4rIWr3Xbe
aYfNqbJiKDkwgkyQAHKu8y5/UZCO4FP0X8wsJp2qohH/drlyxeJ01po9TDMe3A6DMnSlH1ua854b
BdymLPhewgxOnRKbD9TeETNg6z2tpcG50LL8Oa7YBgX6Vgd2XWen1PGnbk/Wqa+ASi1G7QqLKt2B
YQijJ8/F027ugvP3RJWcbx2FaLtbdlxUtzzDXWwj9y0XL0Bo403Y8smnxmkUutGIH0MbrxqfUNMQ
O5qYgwRAAkf2SJMhx3q8hZwfJ18oy/o9+pFSPeFYP4AARFGUbB02/rW1vkoJp956yjc55ta4dwDI
e7bU4gX73XtXENiUz0f1z2iW1CC+jVZZom9BIf8ccvSFgO7RlwSiohHvNzcvWzttuIKD6PFKatpg
tOoHFWU3ppyexZMTiULril7Gd1dpb/4McEW2w/hv2ahMJj6YPgwsiLy3HQ0iRZsjGhalnWu19znm
9Pg7slQcBGuVz5vzGIBqmPCrYL6GVgolb0yiAxp01S7OGSmq4XanVfVArKfaOU5akS+k7+Z/GTZ2
N2dr4rA+se6tngHeugmsyGxMMMrO+5SJYUHXcpPS6PPqmGLtarY0fr6BP3A0syQUc2D2g8OW6S5H
+gAB0Rcx5iT9+803sf64Q5BKLk7DEHdQIXrqc+Tlvomn3Fpp9G2tYPypscEHSPKx0ZGtmOg/mtON
Qkk2Pu96MimRp93Hjmkz1wikjUlFsLvZIdXPS39H6o1+kmyxM9DFcP6qMh97JdgWsN00cQhkX9Sc
FNZ/eV94IqMW3xZEmYnlOhJyYmqGTSlk9uFU+JYCaWD7BCWIfL9jprpRdhJzCVlUAqsoLODRHKz1
JA89X1utLuSEVslCkkrjLE5zlE/OJTjkF/4zwk8o8iwYC7ZLsn51W1nkmZVDI/kWPp99bB5HkGrB
/rIsoiAr/MTtcicVAG0X7nbz+KzE1150MiTto2rsk7pbhQEBIqRBl2Q0PkqZ3EV3JNfewP8YugA/
n65H58oYHRcwyJXsOXfVwyBzrBsIZPQNPGPCpINRhND+DAgTQEuL6NoaQOOFryuwujOwhzXdKGva
spN0LEhVF+fm6rpskl3aByC0clRGN/WA4+Y5jJyhZzOzrL98ZYxf0XrlLeu52eNsqnLrp2c58O8E
iH/uGyv3g4IYwLdavE/60rY+wYc9FHIosrac8U0iwxBXHhFBbPqaLdq8bjcVZ5mZaTnaNNr2r8DF
YdJMdrkdfVCqeGjVdRmZdPPZVjaEddpxdPAEUowEQG3GXzcBH2Y3DHwK4pWr6ccCPz6u7vo8Twx1
pM57rLTWofjpUQol6474ZwxkuGZEOZXnWjwoYYV1PBmfEcPOp2XT08ULx9eJAWTW7thTCIfH4Nkj
xkxoEfHq+rKKI+CE4KrBcw+UWkEtPcZZ7l5qAdq4msyQHY5ouZ/7A2YiAR8mig/nHrduSNsgCUS1
gQ6Y5BISPsUmOBCHgdh0BA6oweWBm2DDdOH+QPijo+5Hx4wsTgB1rG4/Q0OZH+Viv0SVmrQjISgR
JKs4c5XAMZkZMvifE96V8mPX1J688yKT4cWHBmGn0BNvI7V+whoFDhQtFBCGAkqN86NpupjC6xkJ
ZEAKoRiPQdGjp1obtJCjm8w5/nmxQEcO5zfpqgTlVvwv11vvxdDAHyM43YhZb3qX/WJI4SFHA8DE
A+jCryHihF3Odiw41yqNDjCj5ogZZM9hDyiIJ/8OXPMVHo/QWPDR0S0dUZKK2QFEgt3neyjiQT4n
IrEsrFIliTXSuA0kZuODQBQvttxsIJOZ+2Ia5P8UQK0RP61O7hr+sYYKycTqKamxGKWk185+VK04
SC6rm7utya6LelzII4mfedpsTBOtcaYL2jydsNg4t7SYQrk5EtoIMDeCqmgYhyppyNiqwVI3Y+dY
KxufAbbkzTCz8dsbkQas7bN8Q8cJtWq/nd4+uKQ8T4+e2fIie6Xcqqk4QCKuNrovIATr0SeA+2c1
xZa0C+Vv9ydLHF/gUuE8chtOIQYb+0VkVjhmN1ypRI630cJQqsWcNdcCl66ps66KZnKkMpag6jow
8jlCWQ+XrwjaD1bD0V0HFVDMGZDLAo3yaYCklZqetOvJqWNmD5ZkJQHFUITtT4CxMVvZMDPVIWTh
9TpWMrKU3YP0R2IMRbymoGsbPcz4/1egy1Yb4YjWancxw3CvYu38L9GBSL4Lgp0vStgZ6sWUSnR/
Bih4zJM6S3vB6lPXL0s1ehGLqHgXMN7+RzIiv0ETQlAb9dP0EM/vKLUf7zGcEbcrcRUoWVl7hQwv
lOWC0swAEQlYdFCpxwIFtvCJZx+wTfh1zuv/9bLPc9PVMu33jo4xEZ2Q5VakvG65B6FTjEhzxncZ
k3DE05VW5zyvH1OBD1Lfhjoc7eQUW5ACbRQubOYGobBO7OAgGiD7u4P5dalIFM2/w9eTSBKmJEYE
c7gUtN2M7AsATrQZaq5sRDpPCjofmDTsgyEf5kUysesBQBnwuol59aA64UpAnkM647vf+bBNZ+dz
4bfhYNeLGmeGCvfvQ3duicAuimCucZCu+DTiU5tVBEu14BtTSElzzyLGUM/DhL0casG5OOHnRRGM
oFgXRAn3r/QvofDJC/EYaDMiPik8TJDVdYLMl/NWbCToHJFa+MfBqX48clJx9DzO08B2Mk/uXCXw
+lSwI1iMu7xR8gtWYv0WG80VuhM58SbtrezOTsYL5Sc1c1eODenkrGgjzDMvwOr0A7JpgoZT3RIc
esDykazseQ4nNtlnDKEcfCVSxcRXq01lkZ0OI2Qd+yNKQt4U7qlp8Lv3zlGg72WgJapj1BZM0w3p
oN0vFUDrD+ULey22e4nJ4Ftk4/HTvXcYeA9kwtcWH/y72A4vf3E+JR0WfnrCnuJbHIhzJWAoRdOq
8hfietAfo4qT/3r4AbvCtadnsAOJwR6JGpTbqlBgxFCVblbdpgoLvRlvOeCaVEEWTW05UFH8T3Td
KYw2OdmaS/gl9D+sW7oMwkw6sJaS1edY8FegtNU5xeu+iD8i3NhvQeRH397a70HEVAYGhKHRV9yw
gcYO26wAz9kmSX3NBZYv8vRr9IEvmHkoxxBc9EHcuGd/CMHH0OPHyLtjKNl0+qqBni6Gx67JZOpG
1Mm0QoV9dErij2OQ1e2V8v5v8+emaYb1lXbNjsAAKcMgeq0Iv+mplvgn0YvgmhtLvIjZMtWhJuky
EAVtHNw2fNmr2ZdBtY8YHzAeqYk1WqPNkY3HQEHCiIm44PaofWLJhaGo3FCfiwFCr2ftsC4aSJ80
gv0Nl++1t/Os0yJfue5I6i4Bua0Xkzj+K0udsgsfjVcIp8uY80qS6itk9POs8Hk5F4JIeaYKoc3q
TdyyjZSDmmS6uF1bWbwYo5hie+vUWWuO75+w432eCLne5W8eAGsw8fnZG00fmDM0yfDgqyCrYTju
g0JJpjrtlfDkzdowR0KKyFOqPWDVjhBYa3v+TF+YwVqLTs+2dGTYOycMxR6gY2/o5ayVuW9sMesM
omnDm/uMn/pzgoGKBcuBzvzWiGdKzSeYH69dZ6Q04NIYrc11skINyl0zaXq7QJvwvV/zr/pWbKp5
+dWqCOF6a1PyAM4taMrLHtWZaUYg5pylSjt6Kg6O91RBkiMnrTtSpcRkG/ZaYSsuqb3ySzcTsa9E
Uwx4sX5n+jjC27kSJ98hiwCoED58rzSSkZTh96m7KNummkmi6C1+r1jASIHZlOly1LLiF7fV7BqJ
d1OFH6vLs+DR2PTzNTKFIYcShI5k4TadPgeDMJTj9WUIzcuBFnAB17EC+nn56a1Ct5S++maQ90Ex
WxrNZAxQRMD49ztHK+MNlqq9Z+VHmS/Z9XIfl5c6ZH6ZIjKSYORVXXsQHF55PMb/J37mRoZQeXS4
Ursc2RR/BmzDJrUJ2XwiYfQ5eEeuTMyGHodGo9sQWxCB1hm6cDCD4XzkY2oco5SLSHwlqEjkNLuI
9YihywfMBkxLzmlC2cv22iWwTMFw7g/b3ru7Ohx8eOKnqiNy7EtQI/hUo5g/3AulitnGAwRb3dXF
N1nPxwhEsIW/LN3uS53A00q/tZIyxRObcxpGegbVABzQUwGHsfgY7SAN/C8GDskqBnc1zTl96/p8
JMAunVdWLQDhphuEAsreyjJZELLJ1A9+71OGskSW4sD8JdDxYqao1qf3YrCAP4W/jOkvZeKds2m4
hELXH+EbXE/dFU2fyMS4JSM0nu1s7PhIN1Db/nheHI9Y872hC9lnKxNepxX3owZFghosUaW2Ar74
WWK4C6dU1EUQ2/I6g70MR1q95Ysy9NiOZg6IvGik4hvzIScv8b7SKxMT5y73yyVl/MPaLwcTjY50
6yfLLD06S/v0oSrjMXzTFg8Z5ph18qTug8AgoKxL5EAhC4a7TbjMWvrELMsNFZjrB0u+Ka7Cn9aT
cK0YIY1Pr/8RZl0+S1pjZ9zrD7saDwJxz+YJmQDtYBg4NAYP6hZHrL0ZtGFQnAD1tDTvpdk1K6Ds
8SOsM09euUpXq3C2DZ84fIAJmQ3L+cszw/p/cWPba0swV29rUb7nhoe5ZDDmMmPTNyxCtLHTfyCU
uh0O4+bPerLe833LzO22kj4eWyrULpKeU0na0lR9MrmPChTYJ3BD9B5iSmIWwpXgbKPewt//GXiQ
igivv3hok65mDHivoSxVg4AhZDQ/a/IqsaCGby5XI7h1pt1Bm7QKhs8vcB+fWlRxBJ2gGvLQNnnC
PkhDgYsdelv8XXi4HoC+5va47EA/mXlBxghIvox49VR/tJuYvAwICymxcBF3DcLuqB5xiwdAdYPf
Gh30kSgKNyswS3MFjLQFnOSh+v1qbBU9V0NkYRxQzjwg+NiHN4k2tw0kq5F7PtTj9v1kEZzawI/Z
iOm9XOZeNGUpdO2CeDu7nauk4toXMlSMvEgaquX00E3kEhnQutbhocCV4ihPJFdze+UPmxmKcK6B
4y9TuKwRgPFElzgAaucmOz9/+qcwqePpwu9qPmfZlCrmEhpVd7KmJykagxRf8OoF0SHh62Vuo9LX
J4auDlI1rbJjGqd82mxwc1bWch3U+XiPdQaGKt4Qt8nN84fVhVfXaXdeLvef1v7q6AG2x2Ikm/cm
2m8s00tCba1Vr0GYI73oTtrQ9iV7e/9dwWIE5edWqJtfn3BnIPpfWOkGTJTolPysqc9SAfeHnolc
x92kUW8sD11qO4idSyXSmjxnfJNBApS7lvuXVOzED9GFamln2VhB1XjpYzlZpiX1FhYv/86tK4E/
Pce0YFE4gRSA480IEGbE/WmHrHkg09oiTKPce5+V0KYSMBA1+jrwmlOArpVVI4gm9CTdraA5AFSP
BQnotLd5HRiIuEjgqfnjDPmp19y1Obz0ZZZVzl8sAc/qVWGdBxLarG/p6vfZ9S8Dr6VJWUUU8AUx
3zwW4kpKrW8UHeZd99AYfJIYILMDJj8zmN8xSwGyjKLvUclDF6lD1Flzr3kbATvLok002ZhlsLWb
yFTL+DwzrgivXR/E+uiWzceXA8JUb0QCL79B8Tj6+W1tAlgeRPZhpytDjdyLd0jllWy5N+wojheN
vaKJV1NssKiUek/fsp0rjDOKBNd5Zt4OnZ2CsdhsOUsE9bIf0hQ+pxju6+vf4zN/LqKtJ76XuKTB
VmTwF1chP2WMQadBie2M5Fa++NybHbTJbPtRFTHKiV0tARyHObutSlAGwLw4BwAthrYnmmHjt57s
LkM5I+8bgdtUtdwRkLTxXtst7Gwhgi85ub0WLdQzPVffWrZc6xNL3f+khrcd3Nde1F2gy1pYiqw2
Mr5AXS0+M8+5fydNGHSH+jiJzfpHRS33O6vDpVUDm2QYIDnDoTf13HOGvJrGUwBsmqqEZuyJoKzO
RDfzB0Nj4l08Najby1Fehn3IrxB5p+3d4tBMiK4AVk7L/QD2slaN7kzhoK/zgFO3ASDdj98QMpLS
7Fq4hMI5Sbgdx16tof4vrIuHPsY36/7bfzJL7UPu47Llnv4htqsS/yoNMaV0PezcS/ZCJffV9OZW
X+cUCfJA6NjXtPYriWhKUiGhAoyyZHvWwYYhsPH/5MYdlgc3TenVQVCZwQIx895UIlrG+XWb/L4M
YTaG+7AZL+s7vlPtwZduoPQREhAcKc9LwdgSQJhICcD0uDHGeURXGbf3Dx1c75GW2ukCiqEgm3cz
+rWXjHhGl2hd5ycxksD1jk89cyzLdqvlupwBepJLlZNoYaw2Uu4zhJ9qwbaIo9JZV1qX/rXcs+kt
/xGRG3nyM78cNgvvAv2aUt6zQXTakrExjBis0eJiyZkR7hfro/B+bn5SJpXh9iF+bgCpSdyyE5G1
l48t1iwQjm0MWhC1HXmsQolKMz9OdkBpIuJzIxOm9hdhatJFx3p9fuk020oQuwYDFIT0qVzL4UvE
osK9PacX+WIQlQ4J9C2c4ajI4BDENPAaqEr/2XuoqjAi9RvS07HtXDYhDuPQApVgTLXIPPe2i12h
PgEYG8jKsDM00NGpVd77zl6j4gIyQ/fS4ceu9cCjuSoRaylVdqFG30nIlwSG7EL7N7FTdObh/w+R
aTD8/zumYnvMEaU0PSqPjSY0AWT45jNmVCU7+NBMyze9Mq5k1j5JthkyaxIYyjwC5djxGglxGla9
u79zAWlsQUnQY+yc4E/Q+1EVuTZCJ4Ab9DXVnpgbgFDYs4/5/qmNo3t4gYa7jFBou67jn1uW4G8W
HpEXGq3zb3pCD+gtxIQj6IR1BWH/ISjRan6rOeg42MexVxPDV3QPY++O3ZHrMnESWOiomB5c5maP
YRfQ/szEolZvS4zPmHIrZA50BebSRrJFatxCqGis/FxNnJaWidZArxylQ9Nfna3f/cW7UkynPOJe
0UlXHadz0eHVnWIlz5JqMGSguCmWLUxtCoC0+y4bAnqEVq91Mneo9ECZcE+T+dLzHOWASyoIB5kJ
fSzU9DTXAoO9g6H6adwxB2zKDEmUuDBZPV8CsiWIh8jBx/30AIMNvZbJmjGsXww/zmOjm6EA1wUg
V2lWMLdTNJ692/rbATuXQUMMCtRvS7xmOmoeT9ys86v4C+nMpxUVN2vt3DMwHc6f6xWdGFaXl+4c
5pwrzMrMSc6Y1eqnH5gBPDLf5zdIXt+VCAkHLeiuPbb2CpUsR25iOayuMHodejvznZSkIfZGt+AF
oCXpYsnaZkASejoWjXLvYMzcjpOaDzbeN6UrxE1LI3aiHvXavvSM/GOLvEnyyeMzzmn1yGFfzHZN
mA6Gq32SlTGFcusR7cgURx1RXQKcOJGskPUiHVfeRqnFI1h5adFCF3f4eO3Ai78jXgqRvymhHdyu
2+99QVS4vkY3Do/xjlYkikyk4PLMnQarN5570UF3Y3LNVoK2XDG9wGzOK26H7ezRcGPeReB0ScvA
5ZMMZ4LvC8P0KXm8HeMecmJ1VvKa2Zg+vASumX+3iy4yKFRnDIuxngiY5+Q0zgNbvSZa4pwLwRou
e0L3q3bXdxZ6U6eBmvfD/PhMn4x2mN1vx0aN4nOFFU7HXIWC5s95YPEMsfKhaHBjhbhQw7SWNMQ8
YODEFZiUjWI6bVZ+hsbJl4shVADvy4Ztv5nH4Rrb5y11GfE6KOa//fWGuy+vGVRyMQGk/nFYCY/8
JyQXfsgUJGrVruY6OGXTZf8sQdPHqdOhtwaax9AZ89odu7gBeEZGqfJXcBEEOM+F3VT6YHOGatPd
KUiA2amYPW+7iA5lfH5Vqz3a7OS8g0DjjdOSI/eX8UXIck4NgGpjIxWP3w4vombxZ2PXddFarr3D
fBff7Xd40yqyygioo4te8BKDWV0lOBtqBEHXHPU3eSO5Cuq928i8s/c0ZWDQci8hdtXr8Td9Gpl3
9orfoaLpC/iQf/kG04epf+ffLzbqSoa9aeTqrv6Qo60ufUXSPNkdTku1TLJebZhtrdzFa3IzviLP
3SoJbFnmN845nZNJbpiKAgISskmGFxF1WRDoFwMy1rS7Ih8mR88WingcplsFGuqEnkPT5BxOXApV
cmCCpT6EJoS8Owx7+SkepBWGJEpwN5CG77ZOTTsH4PkhK6nIHTNOxWTOisNhKQRMGyIH33CxEdE7
4FYuRrhimI215SoqVTq0hmLzVzGjmJocxXpU+a4eBHDw8yv9nzsnYB0rXEQyvC4qDY1dsTwaNl7V
oF9ALdqmLkF/dLuJ9P5PjXGwEkYsHrHIbyPA6ICFxI6pBrIadFTmwc8kWkkJY8HYTsjUrs2ort2q
2jPF7srJF66NpLlQgTgICMdMp4zSdf82YHtMvGVS23f+SO+KvddvbADYIPQC9I1MvyaC1kN1ciWM
D0AqoShBi8SjoKZKE7SQ8RJ4ADUAQzTFEh23f0trO/V7ccP3eAw12kU6wwo14PGBgFN5fZ3o+rGe
Bm4WxDHeVSR185Xp9QFc/B5meC1OyZmkWawS6aQA41PTu764RGJoB/uzGRM17zepahqblxaioYJf
fryHZqJZvaf5HXBr/xySZYjkd8A64GSqMcvWfAXY3tvNaTpLNTjXYi9ncNWSl2spNvKkC8J1MZjV
oAmPamCvIUqIlOUhtw1F9yyYFLrV4oKt3oQ20ddKhg93FIUkEuwLm1t/fpnYCTITrIZZxrpBZU3G
f0t4szjTAsjYgTMkBIqO44Ds/+B7JrKLL6a7Qch85g+F2spAAfLgR76cqO3Hpts99dgShq1NiVsU
zVSui//3DrqdO7N+1cSzlZFj3rldVJDXbGBVhPGNLNXSLIjJ/3YvL9hEo7iYm+Im/YQs6wv3q1Gv
rzB8xBBO23gFCsKWZaEPFFSL6ba/bRefv30KpSMAVFjA//HO4gvCOcSAYsqY9KB3WPB7bn02EvfX
jBBuv4Eb0SgC8sM+YlfAIlzPOYXqkdOZOlpHS857h2taLSgev0YV3nkSBQp1ZAh7Mj8xpxqLTnP2
F9pTVpH2Cv/3811E3cb/b3XQhDW/Xs4kzjp708jad/cpt+bhZx9gSLiStlLKlmopOkQyoo36eZ17
Jk9jGm6PL2CJkqZbCAuZWelW/+E5z8HxC6A5WSvjaFgk1nA03qLvV7v4Co5vGfaGzcMdI+9wu3lD
+PLiBwe8i7o1m+tCiASX3Wu8/dZVu8BPnW0hgWm9+JAKAZUVGcfSHAN1wzjTrQRzBZAydbwAxOOE
NqJ7uWZVGnHqqAuR6Jo2zfl8ZYT9AqAHnhJNiweO+3pW2t3kXIIwuIB5RVmi0pwimPD3WXvcdyNw
m+oNmKVm1Ni5iOs5vrDoZ6Fzv12EI+h0TZfyln7cH4AcAECRYUqrBixFRPN4fCoM0FHglo010AjO
7vrM383QBQbwCi41o6+JevviizGq3vr7u/TYE7n91rkPO9dSLK34IMylnz5vjEiiVKBHiKqcXsn1
7zYameL63Cf3xx2ALyrWqBscwpaVucYLvLeEdI5+aVw1FI8rwf4iiBciVgZgV6FrnTymK1P/qugY
Cu2yhyoHqXHpzyzEP9L+7v6JPqy6j+0jOBHCZoDPlNI7z0GD+cga7TruIIg+HexjtiwWwBVbFtaO
U1Q8sc7Z7Stgvifo4JBqnEpMwuvWP76VGyiUDzaP5y/wRnbFag9DHX+14xVaYgCeSoD1Rdg61u9Z
BYTQ7SXwNhgPmZ/4ulD5AYX3sDHCF4OAbSMlBVQYOKYscbvvZrq/C3NbWV3iy712hUqz7O8ESwhy
n0q8g24ntOzhpmRI4va2F2Hjqa0l0wPkizlBts3vlWAECHUoiKes03OasDX7lPUCBevMJAFOKxkR
W91t23vTmCHZoSdysmT4VCzv+bSfYscYNjpMWNCArtSm1WLuSjbpP6wHNcKaJxQXmbc4K2li9JeV
hbZYnKjF33j0EOD2DgIUVa7M7xTHTjAbKTbWjXdFiTjqxMWGhilH/uXADPPgef8FmRNPebTek4Mf
wJChrFac2cVth/6EIn9ky30WPCFqo1Ia0v1nc2fSlb5O2sDAz00EtsHVDgIkSi/Z9kffYwgUshaN
IGiJ6yiUQibp9A3rg/6K1nbS8vq3bFZVhRi+Jl3+SJbIh01tARlibCYbEahb3C/ghtuzwEaLkAl7
pCpy5BP2Da/NF5zmIS7TSKPG7UpZWKBsHDhwO7ESZNB5uqY3HGoPZCzaK9VHM2PUQUCTwYyg9uM5
OsJwSmI2DpT5WPvr/cXQb3WRsL0S808FanzSCm1tk1cBSTh/J9bw9WJZTD+Z6PFNZRybNbjLPzOp
PmPJAVP3arCDhEZCR81hNuAvX7K0IoKvUJ4Ws2NABXq4em1TE16bo9oMqWqGvYdLEQXpO0RQuGLj
asOcgRQzkoxXJ3k5HNIuKEMZ6f6ol/rZO9iJX9gilOPsoJ4dMIktzLom3St+WwUPDdUWT1R2vlBC
HC6+Jg9hH6HI8g2oJp4N8EpsuMwruv5MUVANigSrZHCh+ORcYqyWgUsdRfxaMdiveZZF6kYn9ERf
CjwADdmUDjeAjGxLeMPmL6Ren/m7pj0kXuxfQ5YHrLZX5j/q0xW985jPcCVkE8rye2BYmrW8SAJy
WaLQNGWZTPdfdNDXvFwF4f+lCNjsjgz9SbiDoedgZiyuGhZYsjX0dhGEpJc9J5hKbR86wRDwJxd1
BmJgO+tQZm1hg2VSnuLkv1KEbogYq8/BKLHiQAvIo1zBOtJec9W7nBYsfaCYRJqU25F6lwPMCpZ4
8611Eko/+uVZM+xbyGJ1lfhcTz2Yyqe3PgiArZWQ37FezUdIDG3vvMUdDcz2Mj+LoE95L1kkY6Hj
0JX7LPC+5dQue08kLsSyIvNVj/nisGbH8lqktxkIaiFfMuy8W2jXYdglzRka9D9jHBxEcxiGdJRp
MUod5rbGxvA+8BvcGg/CrTkclyPt7LhzzF9P30L2pywhXtgTDDpTcO+0Xjc4NeSFd6SNCO4sLJuv
CAGnlXxTC/sSiSoCTKNSmQWQM2JMGoXcH9srPd44YK4q76reWaXdn2hgzE+CAqji5HHP8/pD2Q6k
y/hv9oOUCCX79RUPvkam3A7a9HarumTPG5SlAiCYGZo5dIRczN6++ATIbG3gh92FgByYYyaWNfsL
AMK9yh29lj/kW+jp/2YwWQq5+94epNaUFGZmpNSsMsQxAg/8jvYfd7U3VNyuC/O4aKxon3CMKf+c
76YLVYwTLjN25jnjWkIBBeVa0CqP1T4RxMjNKjDg/sKt6w4vI2UoVIo+osHJOUGgqigQWL2jw3S4
dfRuZvt7uegYvFq4UFYDno9tKJT6OgaI66tsv1bdKIUAaEMDT0CHVJqpVIH/ggXtLeXhKZd2d1+M
O0jNnN9pKA1qn6T9qOQN/OtBxUi0c18Mq/62ZMzgZ48LD+CDHhh9/OlRVqFoapRY3cyUZd6TvkY0
BPdtU9GOe8NqBFrlUGmUY4rBi7kyqoz9dnzwp1GayZezI9PnMppkT/3MY2qK6gexEsTg9AZIJa9n
/LPRhC5YYJ88VMwOr9Q5MGirgYmEQ+PoiQxDlOKZnVV0zZOsBIZycth+BU6g/GYQ2xtjsrN+QhO+
kWY4Xn1v4fX2eQROS8NShN2ndSoYB6SmoM8NYMZQR89Nxtlk7yTxQT3mO6xTEKWXn0c6MOkuxgfj
3go4yqyCyVXzpwy6eSrGJW96OUTgrDso/475yKUjjKOzbs3cCRdOoOws3sJvqs+MflpT7sNuXNT9
7h6DUiLl/iCcDHjdNvQPZk1iRPu+3ImKfc7GbVYYMl2kJPnrqP5MFxLYqp6x3hC8c1gIm50/RYdO
PtMV8Z8XDjKV2euCta2SQFQixHnbgBFaYlvwIWOf9vBeORdpWCxhBx6MiHRvQo5A350zmrOW3UfS
HOupEunhMXYEApgFGwiFBzq5LRFO9UbJUxiZIbnahYiyyiAH7d2cLYT0NT75cJq3FgPePqt4lePM
gKDXeTwar+GZgV9akg5b5DilfLEK22lA3dYW0zlzS0GqS4WabGklgHeJ4I2g+KsB6Gdf2dJt+MZF
Y+xcZIcgwj67ZMFJEgoC/Y1TZutB59dtekI8bBtYdXA8cCxpFzI9cmtxMcM1qkxDm0rR+riMvW3Z
6Ps9VXcRhHogv/Mkkgi/9CP6a3jI4mQIapqGqhG/PEru34k4kujqi6CUh7vQ2koeTqqmO1q6+xGv
K6VodqFUOVtJN65tuj/sQ4zrSnBYloMODxfsDpWJgM7E+TkMn9c7j13/FycW/o/JVunBd0jIeOlf
F10qfc1SUtBFUinKs3CCBt/hFMpCj/ZYh9KzJTTFJuk6GWa34mNKfc/tO0gNalA+QI1NR7nSkOvp
SfgMjhBFfNuviJEA2x137f+DLvabPelV/5yqe6L/xTCjPaFvXtQP6I9L2IjK0dp7DPBfd0HCxM6f
ytxPNX7O5jj8kYtVFDqYgpnpEzOPu9BqhiFuFyfkKU3/ohvbfarBJ7wTAQUtixA0a0qAP/gBw8qE
I7OMuMndxc+xK4qSlC9oYYrOBZutl3J8gpPmlc06cWusijKHcJK6Zf41e7bTEtqLyO/zj2JTd/1f
Dik30BZV+/Z758Ann1CtJDa2j8LaMj8J6EpbLR2vJqIsW/rzTwXY3cdCpUz19iHNsGmUDuIJ3fez
+UenxtQg1CgwHdDNq4QbsMBEQVjkR8QQHZ3pgRbefQa9PlOJYIulUgPKDiazxMOOB89268+rb4J6
+WuhW5HCc01wqE8FBOuuEU8I2W1SIoOTAf1EQdycbTeYN3sjWlV3LII/PMQbY1/7zAFVb6eSR5gG
/b64AU/kvX6hKIS0driD/129xORtNsDKeqx0fMwSmFhCAb/JKyS0rGzl/91ElElWPkstxc0fxcYW
HhH9OZpcHr3yIywVsu3M3Y0Tc95vkpakHpEua0V1/ABlh36SIvdL5xK8HT27d65kBFN5cl1m+Jg3
H6aOk6soYZzUKrQTvYX2dcsxE2NAV7JUYWxNQHcK8yTTAMdMZfxFc2c7vakcDqDRdSL+cXEYSeVH
+itrJVqFBk+17RAwRf3/y7IKxOcRc89JL41+gd0C1Q7IsFr93RSGO2t980NBtnTY3g6iSMkoH16e
yyR1yt6XN0C08g3+EwssNKNbkUUcGrwmaymYJqT6giEfBnw3SvuWKtGlJBBIaoPAsvEHY0uDSiUC
GFhKpjPbfqVqWIzjuhtCApAEIe6HA1/Qww6eSpex1/qQNEMKkVJxi/+AtCgpl2i77OT5x+8rWHiy
mtHQb7oFajbudfb13FmdlUqeton0U9YeS9336RAEMGkh+61EMLpH+ka1vqujvVgOILGcj8A6k9CU
UbdAQoPtyHscJwt3U+Aj0AG1lRP1yxkav5m+cmZhyB000c2Nn5JtOqKNVS0ASD8ySbjawWC2Ei50
VkwGwnBhZs6UKH7njTbfuSaJIFQEbl06HO2hVAeTw2mZqT8kxnLidRmheO8aYcm2DawbX7+ptRB8
XJ7zReMyxrmUrUaReRflunW5qBTJh9Y3boBejwthDXzH1nIWxmyWiF4F6mPDgzsG3cUwSxJ3yg+P
xbrpwhw75TT2IFOLrO+eoN1QR5jQvEymv14jpLJGkck5CRclWPpxK0jwvENH0tS0dJn1g4i4ZkVH
Hj4w23BQy9XHb3BlBcw+XwsnvNfoCHIGWUiTAvx7EBfN3t4iS3A0YBj8blTpHgMQi3Z2V3CAFlFR
zTgC49kGphIc1NOZ73C/48bdTcdWedlZ8AYvcFT52T9dMTKrBXaM5EdYKvsx9FPUNbSU9gHtO+4L
FA29L0j+H0q+uOyFbqa0zCOKUDame9iIpRsHBVI8m43ZhB5MBgVYoErH7L1jAQGZrw76CVPpymKr
WHic69WBhKOB2Uq6TsnjwisX2zOuV8XPCFdCKMOAUqu/AuA8bqHl7bIY5je6xJp88ulQgbs6dym/
bv9wQ6ODJ1JdCBjLLPUzc3f6R7f7IRSKN62MEi4vaUekltl+u7AKCEUvLu6GVkPSxpZf+ecKc1ZV
MzZ7usVma14SbjJw+SnvennImz5gPTklkiZByIxNU8FDbk6RKm4GtoO6tVzARsfThTwOQ6CaXAmr
togYLWGbT6DWm+3FEJ72jEvuxBkkP6/LjhavzF42cISA2L3TjcJr5qVO/RjKl4XQT07paJhb6FaB
NKfBidRsvTLINIKfm2A6E1dQGhUAbx+8iyVrOtjFUQE1vdqwWHL/4HCj1HJ5yD9+Y9PQHn8IoVSh
FrTuMLW8ULFF0yM/9Bhm6+pwoIM5wrZ5Cvsrsk+QvhZ8S64ZdADV2OLtU1Wn3ZeQV83bpBmO3RPh
yd7rmprKz8d0ftxxv+VvPJLGwguoGjHrpWcNF6NYpg2r8Ub479SmyxKXyQ83QkGErY+k2xjL4uxt
ehGyeGCWlZB4FHKLnuPDatVvL9u+R8GKeoTbKqWm64k3TX0yHibb7CK8wXIYpIiXAtACJBbk2dtq
LiJtG1vm996RCNmaHu4yJr7DjOzoouTYAq82RELtg8BhcpIZUX3y2iVgQtAqdx8Co1R6uQW1BRXz
5rN7olI4hc9A9g+Lr4b5MS/tOnwicjYSsa57vM7Wm5tCJXiGPGSenb0OlX8iKBLknyU2DgZ/quSC
meMJ87PnplJsSQ4gM22I1q8moyPMcd62w5ShfF3VMGNI13s2kHHxye/Dgnq2zREajgWLEs4Jv1u7
1Z0FLzxmGe4PL+TGs1PHBF8p+kNr6IMeiEZ+xPdoHPkYqpLz7Hn9ncufEpZRYbKvWnrR7zds818H
p8xWkcttYYyjq3mKR4stUnbf2pKrQ01FiGa0NorK95vCq0BOxssUCKRvJXQHIkFb9SuXPnA2L/py
d8wsHn547yRfpF7oCQcGSi84Zj6YfpTDMoRIVFsSUMhaAn8QZRtZuNGk3rz9zVHSnAkMq/q6nG+u
mX961Vz7Im9vZ8EZM6Txf2vuadMyawjZUNlYLaSo1ObOVoA0HiJ/t5fYgNz4ZtesYU6COhky302/
LZnkELm2nHH+b1VJg0qHyIER6Bo5Ukc4QG+9BH+Zeuxi0NM4yTeHQ6BV8/ZySpA11j4Bey2v/OL8
UHj6AjSI5/HQ0ObW19zaRWmneDyZNnhIldJwcAR8cgcp+lCEHFHESDSaeEFhT7yGTHzsl4CbODBK
O4Gei2n1iWeU5fyAbcEHdanlxrsQvS807su0qYNHNcZVxY7Qm8vYgO4oeeBcUJqeqi/hdVGsCDks
zbZVN0UJn335Hk1yIIOyPpyD9ic+eITZOXi2s3NMQ0kZEtXsAaYvvu7mG5SHeA5FKk4PJz6jB4mG
8DO6IA6iIOCF/5zR46HsHptAvF5SeplRTW2jgVug+7JAKtVoKGEf5Dw7e+hUVASDlnT/jUiDO3bT
nYV2Cv8j9ccgKAJStKyPrOiUs//mRK5W+PtMSeVgkYCiAbAMP1miO1uHjuRil8TFCWjNoChnLEul
2nJJASXT9qpE0D1o/DE0wl3YNN+3uN1XfbSnUCh0M7P7qxQHgxylLmuKp5gMFsqJJJUO4GU8L6jm
PBKCP+KnRXqaiHyYlmk/bzX104z/g+PJcYScJsqMJWTNqhemyv9JhoJsgSwKRW2SMQ2nQW3CS3Kr
5Lz/VbswViSuS+2ETJpzE+uPYjkwVA38cSMR/c8l1RtRTHT579kClLC5GckUuKVoWUC8oBWsgsLG
I7EhISeHDwIiT6XCGTL6jndEQyF4hpzBgZeNHv10BcsHDg6hJupqKiKUBzi1548lPT7z2yqVyNSz
brPNfeKq9ogrxAR4NDVMz9SHRtoj+nvjh5ez+99qbXVHhaqnLeuDek8z67qwXOq+2AXCt2SGHfxU
t9z0gXAzKzvZDRPgvciG3CEefpAEj+c79WRDVvwpsxUWHbD/MB83J5cR+tW02LUZDHW47bkrYtRO
veBdEIs6prXtJbCDlBmxUAJUcDhwiL7i98LkROg8qb5k1VmtnN0hmCEsmVaAeRmxGYcUs49zFxYg
FsduXklsA8nprOJIPL7UsJe/6Oobvd9e6xiy1slMKVShPBbFIxTF/aLYtun5PUTN+W4wTAnKVHUR
/gY+z6sc3njifFRmHHI7KRkQ4tGiy1kZsgYANmY/HBo2BAkPN4fjEp3Usv/hk0TnZPH0b5zl6rZ8
FJSAmLd8k5K4JnP3w+MdNAh9nJ/7w5Gzdhm38Ik56WIiKjdcikmvWAiqZLglBgG7sp/9zlKJnoo3
HeUIbUbHT9uw871q20GJhx8p+44vTHzp40c3L689oyMLSUMFDepLfUTevG6sPCu1yYj1UZWNbhYJ
0/BdtnhizpA7Zde715zTDegyFnBSBaouiCPW4h7VKaJ1xMncm2dE6TkelZAR/Hu7zZCEBMVPcwse
Nt2osZzHW6br0z5QwgnICu0Yk7sYMOMKMzFpNbtyNu5JJ2S+0g2eBdA3y/hDz/Tgf5npYFCuSlP3
p5uVhF/WtrSSD+5WLaIAWn/upf7SZ1Yv6G7pxFw8szEbV2FzYq0rLAz07w2h0zIZIq9OoZLQOndw
+Usy3rgXrwpHzNta/zn6H7YoiBIa1RTB4SY3/PD9TjrBZs79v50mnzvkE0FfysqzwJxWAwhWpGdT
gyZagtlKeZf8IAQTvT6Wj7s3dyXU3vzdgehJTGArWf7BrocV8AzAqZV1Hwm+OJWYTRk3rk6Onvg1
VRk39nnwVPF8UL8UTFTEtvFD5pcEb6sEkjmr64gamLzoLys7FfWsAOlhaCM9ehO/Za994twQFNqI
eU7wKyYBqEVVwQYqfcElCEkV3Fqb5gc4rFL9HvIRWNUY8OJe2199otEyBu/f3B2b5nKw3hz7TbgB
oigON3tDgcROFSthhh1Zpa/sX+oDFbX6OF+K8OzM6UD/bgykL7rXc4Cr74Y36YRllQe0956m/Bkl
87XAIPGlmkehcAvEJxHZ0GHi1BMAIj212Wp9aj3EpfPKh0jidAI2uiG6yS/mHnpDx5OWrSlXUVQU
/+sRLpAoiDhp1UWZiWoRI2x2iJU4SQP1e02R+RB+H2Pl2iYJMUgFGB/2dTjjh+Mi2d4E+yio2A2j
e39hzqL2qDZxSRrPLryMOFX7r6VbBsuo8fkgeZ0RMucT7WtTipTrGG9yw98S8WTs8G9Qpqof9Pfi
BUWKBRHwwSy8jxEB3DWJWtbQgTSbZ3zfcKEOvK+7jaTQRlDJIpR3CPrzq8SOzeEOb/vzhJFyREgK
RMKVyRMPqE0xCTfVi03Aq9p5rMmYYxGo0rQarLihgmhwMJEy6fTj/ZgWjJhUT9pEQpa2lwfMGge9
Fcy9K+q0pHm/gptRDYhXra992et1aTQ317A/viq+Q5AHEaAt8kACscH9XP2lamkLsoceeJHOXH+8
Ui6Nv+nCkNtl2xMmcks4xztrLTBaMLRYU39EIn7dfoukLoqti2F7wTYgCBbUdZnJBiMPttwRHju5
ijJdR09Wh8N5FJ61GjL+QQUL8jPhqpAiie+E+XGe1WPhqBuebCBKTEEcXg62cWBxw/96bJb/A1mz
rqOf6cEU33oXghT/tIzu6LQ/QSHT9epKIxSV5jtrll4yr26kxJHbdPnrn+x3eZ6+Az5hZbaFOMNU
aSifCByxZiXTezAlpG6+I/qmywVKExXi3qNUoU6YMM0da64FFQ9TXSoHpEyV4WwE7qUhRxbJjQbL
WBTSTnFfjSvLbziaUUEyuitINc+wPiW2XN/MYe16IBnP0YjbYOIvhHCOzuaujkgQLbPEOItdYxMh
dTcnUu7xCWVkdHN8J0ctvikkAJ8tCPn7ijflLxZJ2zaZ7ynUVqwdUw7yPWpk+P1NFYi0S/0e4tVP
1wvD4sSl7zksLIgTfDqT4j2ETqLayJ1sKpKuh66YqnXt5Be/e1OFGD4zqRaUJyrdUdADROVYJmo1
oqXC+cNVxKiutrIOpYrspGmnrs4j+eR6J3Oac+XFfKj9b4OJwrDzkSVXXFwr9TZ1BtnigwzYZAWu
I/umZZTJjVeeCK52rPv96sB7puzzg13RsEslNR3iLsYrc2GjTkr+0CGenHsAztn0nLKkbztQQU5I
/MfF47XgsRWmsHLZmjfpW2L7gKPPh5B0eQpEudxL6xEFR5aYpWi6sYnRx09O7ZExoLrUz8d/pGrG
lz6bkNiFQi33t6byL/WeEGhCtSuG0wRw5vfyet0NOfjaECRCZLKXn/fu28/CPiBItsm/MkH7oPIO
dZyjyTSMYRBB0a3YVnQ6/DKWxMMKnlzyBYGwCNcBd6iz9HtRGT80k9GOanF7ad4csA5mJ81UG3tO
zDGHAZL450y/X/h3TmgxPlK2fZDfH8a9hHeEg//JON22fkH2PdEyOek4yKisTtflzyWhS1X1bNat
VxOvOJBYfnRghDik26JhxoZXg2bnhBfSshdCUVVEq7EvtTL9bFaMhh1DNyVk61/WN7FgTjnWqXZL
xZpf9/2EiYJRJJRbBeuB+eyLRmimMuOKokx6VOcp3Gi72YXJHkSKqBYGlN3SZReC6J4X9Q+wW9v9
oyjWyxBrJLZAOF9Kc4gPi9ehmECiYb+SWgFpBdFK53KcoYFuIPbBkk14A4k2PcRnKygnffXMHEQH
QW/QzwP2cuT5pWRZVMsMLl6wN5hkPy49V2+oEdOy+QOTQBi/LR0CzGQlLyNadLPnlWP+6aqvjtC0
lqtSw5mo5FnMV9brcznSO/IXVNy+XvjSDULUpdlNOAz/FJpR2Hpdi9/m1t0zoSr49cp4ErANLrcJ
momR2FB1ZxVMUWG+ZLr/t2Sub3iBLJE4S2196SQ/HpjUsKDMbt32f+a2mOeb7s0DV7HpK9/7V0Qs
jg2TIkz4ZEfw8wZPR9EuG3QUWG4g9UxRAMhdOGItzPrOHMwii16Y2dMWUgdCEexlH8wKp6MGKXgf
Vv+4PH5pE+vRz+nvNWZfR2dTF72DsF26e8rcxSgUm2rAsCH1FQZpnhzUofGxsxr1KmIrToOOYasD
D3HxMtcHjfImrEp7u6Wy1taw4UHff39CpmagUACmCX2b1wX67mRSPnL6HTGFL04sxpgEhtTcG6ap
Dq24dkWojbZBPGpzmG82jgl8FvXIDpEzVC1QWpSuoqVDB2WBQv9UgGrJIXUG5QTzz8CmQ8gBxAL6
fGRf+HtFaSswEpIstjVycQJrFBsnu6AkVg9wGMT2uzKnNZaH07OWS46JFf2bUKMJLKTD+TnTeDcR
Amzrs3XHcxW3ClJctqIABoFl6OUbI9hqoBJFg1ZyGY8DiEUEmqtkXMle7niM3VlT5p0n86qGhxec
5BOw51oPPhnKrYt00kywUIAip1iZREaLuLr+pRIvMtr8soxKtcLYDUL3ll7vlFvM9wpRv4v6XCMJ
+sJ0cK/XLcg4O+Ph6ErGRjaPRjaRO9LMY/2aCGLTt0jzSMPEU3xYs+du3c2vnbmMYaWdHaCMKeSu
UAdi1bNKfla60eRsA4FDfRVaqPNP2X/++pwuBYH39BBqWXjCWV9AHXdLsob9TGy/h5MswC1YJ6V2
w/aMU6+83IbD03xOwuaj54Jln045rdgfB4sfVLFQyR+JU1hQEmgRyGy/F4KBryUgEzdr/Vqx31tT
Ix28lMmNLOratpycv2xfvQC0VR+C/1T9t7eQPb4Q48qIQ0j1rmsLc2UO1It8i8tsUNwQW8iHIPZS
wBeI9X1RazpSoUHYU0wYY49mj5IfGvZm2jtGpEHWIuD2T+MCrTBunZfenxuqOt8BtT1zfwEWtnyN
DbDR9zQPEXKwYlRlsafgi0ah+cKDN+ShV6a0vReEfSBdoOEfIp9IbZfqFeSp16ik/jWQm/QwWdnd
h8tXJ1g6Jm6ll0OdYuQ8SmJ+pjTKNpjK1UkkZJicGmR18ZraQsc3u15Kex4hR170v/0W/D8xa3YM
Mjiklkwdok2UGaqJhRw8yQkVXR/icbAX2DRY3Gvsm6t4gbxg9K6G79waPFhcDu0kZdIq/2x8LzyX
V6vHT2B/gjoRMFtMYNAPV5xJPG++AHms7cm6lUU4yKxhyy1S0nd9IvVVAFePhQW6bHDC1mK4y9VR
lBJB5mgYGzforAiHj4D20rOLsKuA3gLONZ+6GnHZ9F62xdE3/FND7Bq50NapwgXSVfQH9G202KLB
UsVOkyBnqu8k2FSKakWZLAvfcaqrLtapBV8F8Mvv7ffTKGiE0WidqTtsYaCPJxdDxjYoUHUzlDlH
2st/PGdrXd3M7JhexslsbTrb4i8Rsaqgk371zmTS41EjRV1gnrFo0k/WG+thniCzfek4sY2lLKBM
cy47cY+4m8i9qf3r6pylQm/xC6jEYTU5zlvikczJzMF6oHo8TNd46Yznt3FBDeroQShn0F/az3fw
x5utxm590TfdTOLjiYhdTPaXY4AOntr5+kaOUg3URrxX6c4h1ErhcpcAZrw2Cs/gEVR6qgLwIgD1
+7YHxB6y1q3N8vUdmbIGlWG/287E8w9eJrze1Yu3Domrmrzk/HEqbCWWmgrfoEohW0qMNAbFJBKB
kPOBsArUgb//zyp6NChGpjqaaiGQhj0XzzZYWy1Lao8Jh03WNuGKBLxnYuwlX4gbnmutDcxHG8ql
K8TPx8l7lpxgdiuP2mJf5DEpGk79eJXyz6s3w2PcF3D9+bk37TjUb/KvOYlkMDaP37txDg1rM/Iu
y81bKf91UkmV7ANgc/QbDvOY1toFr8HFinBn7bG/8rvXWE8sxG2kI3aURhO7g1EFotel1cMs4Mlt
5ovFpItgAQSNOidH/69JcYU4OuYI1V1mS6BU26ka+C/Fu78Z+z7MdD80qxMIj6ACDP4fOes8/T+F
yXjP8RHRekSDYkfTy+ngu5vigRVaZaGSo74Mwzj/GL0S4iUFvbB2fD7SLXQk/lTe0l3Xfy43eHoy
+7aCrsfjDbIwIsWmS+Nn57R/SQtWSY9H/nW02VRKrHDMhMFYkAfqtdGZMWAOPHXQ0ozzzbXXNqnC
pXroTfP7egkTpbzY2BAUKMarKcNYbMfn1UGHqzhqCPweTu+tmS/7mdJ3Gw2WiLe5oSxSXxZZw2x0
6Al074AFIa1VtKFaE5+ua01+YHMg9KPxN5Yw0KTTt+jDWTzVi1oHlHoUGTUIZ0XvsAsLOnIbxMfw
GsIdYb3S/Jg5/bDmCjhAsBGNCoQ4mp9zpRf2Ks2ntvzq/H0uetpk20cbJzp/yiVo4Mi8HOLWD1eh
FxZIwUM83nwQ2yaAVcuikJ6qEdTIhMy3pdO3TdmdDGgEKcsQOUO9IWwsdH9YFtBATrCYUQfbcPsc
8jOPieI1yFjL4Mp6Fbc19NP9Fe6fck0jFB5iA2j6ExocSy15e/sVZL3yaAJKnDQZOFIoXm/QDgoA
/fNa6MnY0XHzMXx+LP5tdOyJjedygXKJyhmrOHRN/JsAo0X6/g/igaruEw3UkSzex8nNj3uUE34/
0QQ1tkqoJyopYqBCSkWpoBsBKkOQCUUD/fIKN0Wv9K+C1sp0/qdC5Bf4JoYZoDYAQSdEQSKyqu9p
RLeEtX5qW3SpUIOI7dxZV8gbvVfRoD7Z6IQdS8tKnPG4nyPyRqsC8hRMCC6YVK3er0cu43G6rui7
4nz+9rLayMNyX9qad5KxkAFdcoV/rhC6NkbZp0GtwCCqD/9gkycnPSsUzNLtbH1jjEA8WjE775eR
ZiPqrdflByGPGzjIoaEs+AZCHldT3T3KH5xgKHvWkz/t8e1HIl49Uuiv6Olrw8oWljFiIZH/IM8o
xkaHpxK74q7fAsN/YoG2JkfMNCuZIuUPkyMruFga2UxaBs/setgAKz8Pv1zwbps48+TZ6vZDVT4U
yuZG8vM1ZG9wgFuwu7aIV3MZrhYK2MyD+rBhdlYHUkM1i+wMOZ9owNcwZTO3M4MGE9kujLVlLZXt
g4Q9audir/T9uHtM/zOqigP8UNi6Us/TR8mi6SVP1f2O7umksv4q5EkFoiYSo3ZJJc9qhWZIIvnB
nhl7IDqR79+7KhBkBjVd9YjjDHtPNVsQ9Ev+qLeTrgFua1hmJEZSkcUdGiojBkbZKJ6raZYHU+qA
efbgvistuyU66bBab3sx3xcsUoFs05Adm4Wp5RahSJlw/WFWvNn03obM9iPTjLjGTSPwptx9nvoa
yBen0xkBRCD9e5ip8Vex7/R7h4UhYbehIk0sMCouMSwF5UMwwLZw1nICR6LXFjR9PlKvrVN5MHfb
qX0gAbMa3H5CYTNpnOc/eBGUdjB90wOl3MSEAfHyQGuw0ptmWCFYwN0RaITXBAuDBxQRy1eoZWv9
skkpbnHLX2Q53RzQ15KTXdmnagV8GRbLx0/YI5+rZr+Uoqsqk/60clJCE2Qsslx9iQSRSQeM0Krz
nIdSgIaeMlg4ghMxnWyIsB64fE8cMDB1FupVyRwQD6FsuIL9YQeVmXJ+u7fA8IT7daNX2FwSF7xD
8YsjevWUOIw4vicNII7Qn3gfc/RMDrpu7r9zvARDBiibleBwSiHcA55pRBuhEq3WpmRMpSZlEefw
ym06j6ixwGmqXEdN0dS4Hd2Kjm7E3QBjXPycFhkUcwWEWMVMi+gbYvzuIqH589g3X1RryXoGwEMb
2yr+R6Vi3aZE9s2GvENIHBmjE05Sqp7kgUKzNquxlWQQ6Bog4fouS66sqtKY5oTxnh+9IEWQwEUg
sguFArDwFaQ9sq6L2EHFZrY/MypKsUzEH62GusRrC4NNZbT2JHwkZAFGP5C6kwSqMlXImXJ15Ie9
/91z1e/HcCk7SsbdqgwkCAM7wqfPswxTJqhgpdOLokOCgE+QdULfSU6D/magx6CxcvGfIlpnfzT0
ES+VY1QDp9Ag8X4ZnsBlGPZaBtxqQj3q0x0Bz4UwunlS7TMmL6wavhgxBoGetnQsl0DbdAdYceZr
2VnQ74DMxIs1lTZs//nUDbyxQWlJlCsVJrdGE5rH6g7cMXusGbEFQx3QmR+7V64qsWg+0Xo7i/nt
aknjSgafftEY5ebHBDopJ5BHNAfJolxkxxIDgMu2LusFq33X3A8alB7hykFcXtGskXe97y5xqYDi
xZaD3cK637mMOyII11ecmx9C9mBA5jlNWLx6ey1nD1mehjyFl8e3uaP6K4B02E5/X8zWReNv+8nd
Jrt2eCKeB7rDa3XelE9PaqL9yaywNiixRcVpoRkG9ODGqKF3WNKxOSKFUEoA6AMR6/+D0ajQlgZS
QTVR0+p2yiSrMfQbze7XDWOees+60oolXMe08sckWoJtltuxoj9lv3BCCSNmLUBRGnMFBegkaeJC
iJ5uzTL7D3X5hr4ObLTKkb9b+AHRSnyeMFIedNRqO85lILgt/t6qUvo6U02fjfqy1p06zJ7aF+5U
jlfJHE21Y9HJ+CvsYv57qyUZtrOFvjLmeYvGnzMrn0aX735JRIms2suFiacc6Zhs5SOkzdW6d7/L
BOROmgHLNLT2D2zXSF0M2Cg2TrdNUnzhB0ZapgAQXOTh++qE+H4syOfjIOW/2q+sV0gM8MjQhPdb
aSyJHnd3yfLq3mhXZsJepyArU0agEpR7BFX8EsqDRfaK/lBoO2bwi2o8CGeR8tq48Im4cFw/hJF8
2hUc3u8BZTAbIwusAjPm9fKd15riDA1wyBeKEY6LvEZ7TNHlDNV0bZCwiCBPvSbRugM6z/yrZy3F
T8KLY62D+Z2xTzTymxWJ/xMiL3s+fU7StzAe3ZsvjSXexajOdTLIN1YHA8HLN8APYhMWva9AdEP9
jAxADR0N5Rpbv2OBedJjs3WsDzXfEMbDgsFUkhccfr0mb0f0anaPnQDR8JMbKTdwitZBzVKy4Q5f
W15erCiCFH8P4x+52efJEhPWsj11PQx6MDgptuywumchKi27l6TNhN9UPjjBDOrcn+E/w0T/hFI7
cJQQdiJQxnvzqUCzsd0JIbvcwKrnp0oKfGi+WxCl6FNFifPhCPDmVe67i9ITfReVZwXR+98OLb56
G+NI0WZPW9AM6eZgKIcFFplsRf4RVPWBmimr7nZJ8cpN7IhpnpndvqaK4CnxDyIeJFcxkCooZHEK
JDkrJ67CPcdGwkyko4yZfyYpqqmjqGG7MlayuMifyypCDqJ6GbGcJZl/bs7qzRjG9IUaOa5NuG76
LObfodx5Z8kQqk+sYITQvUaBY2slZorQbSr+oLADCZBfOwnUGQzcuMoAj4NlzopzTpi0w6b8Hrzi
0OdUOQsMbzjOcSg26mXcOWebnzxXTPP9KuwAOd7XZ9mNI0y5NutFE20oWEhTQ6LJn74hQFYR3mP+
Fuf2gMaER7UViEK7agiGJKD2g4kTuiykkwgmMciVdfUtB2Ki2PCeZ1j3JA5vJBRT3BV5ALgE8AT+
3tWRv27O78nn5RVoHIB34fqX5XJosmIDOTlBGt5Uilnskhm76+MWvyYIPiU072kzDdO7bIes3ibw
buz1ISLjT6K/myGTcLKEzHUZ80TBnepHMHJJCtrRZQSDqs/IBUdodZcaJozjznqr9ySyS2Q5ZwfK
xiLk5HwqaOEu3SMyNgIqNJDl5HEaAVoOuKXmY4mUV+ja+TqgnBXWT0+9MmOIjj+v3GrDVw5p7gVU
GylteymYdhyJBLXTj9wutcAWYSZkz6FaBBFEzVI4dhQZPEIK5Ez2Rp64HyXGRwx8vZLBF24cVXH8
9EkFVHYEGilthKFbWnNKMu2EsZu2HsKmoWOffDhQNVYmvqj0qFR0874rrUUCkjnP4yMU5JMqPtXI
61rOrmN/tahy/mds0y2/VHaIlI+yM6PKVX4OUzjBJDvI1UA8UOTjsFO1nNS70t5lkdW9LdBahkgb
Xl6BxZVgpfPjQae+tC3vwlEbs6twwRg9fHsEj6dsgtpGlaaIl4f4LWgjVC/a4rDiEzbQsafM3qF1
tFIYKfe4cqfcUhk4Flhv29N5hA/hRYREwFs4uyTwnScF3ydK9Doa6JQcZnC1x1GwIwIqe/XLud+e
1j4yBSwOYLl2L75AIRcN4qvqzlsyD5xuvqiUKBenwbRzxkgG6LK5IQ2QHcuXhEevywsPIw5XlLyX
slkbo+97ZdbnhbGRZufgyuAlGHc2fcK9e32bcv0+SvFU2TamPRB+XfVoQdNtgVUd2biiKpuKs7T4
D5qSvGZbhRFj03QuhS5SWlze9DgCeCxJ2biRrfLbOd5PAIxh+Bz9YeZTiRdzuD7oldcW2I/M3m76
C8AHjSF/CMHnvl9T+SmkswMvmXKckaY78th7Pt19SFftsTpReM0I6n0aoUgBfrxKELOtg2SltWiD
qlJD4Po4p2jzEUR+udsVljjQqiy0d/8q6eW9NcIL5KdLwFxavHJYdz1YRJU/qdb636lBjEEyanes
shNhxfSS2FUmY3cBDE1gogZJAFYWMgIM4tLrU9i8gpKEeZiEEFv9Me/S+uCd8bytZ4+S93N4beAx
DMLFOioM9RNlHzHHvdXY2blHSFVeFK+N880KtsTNaT91MUtUNRSesDWakISUPgYtDOOZaU7N0+Sy
AAGQIJmwhvr4tWxuVdbx9uor8B5pqaOKXSRrIpXaoxF6Q4DpAJN4krAvZSNDcC682MZA+y4YHwRO
MmHC/bpiY/q+v7npKq+qXZVB2dO23ZsxtnQktxBgZEKsOzY/T3PkNYCvUP6Kh8FqmL4pQb8r71rR
/dAnfnLCq5Uy87raOMJcXU/+r9dlk3aMpW+Mkz57zVoBe63mMnr0d8HXQnqDb6suzPVth4PeI2ks
bGom4H7hT88bW5J5uES/OKI7aEFweO+RKhg5i+FvqrrQJU4X6w6k4cSFvk4gaSgKxVMgnIJgQOvD
OyF27R170XF4EBSb/X3X0LPg1+Z7bJ81WqxiZnxFymjn+rAIy3Ee8f9k8X/fcBqn7TGTt5WxKbZO
nPdYMF0le8btFBwDBPw3KqwAYubDey2u3RScpfWfiEtObav8OWLOHmuvOSECkcO8zRt2fBYCt6uQ
Dl4s8dfY7jyv+xbHWwFYjKjlbCN6nKYsygL05xIM948p7Tvnlz+NWb6M9mb7RPf0xDh8gz4f4Lc5
ke9BGje4ZD/b+R/mUaZ0XsX9Q+Qok2IjVBUTtH5uiIjlIT5KhPUoHdSpszKSgJtZlzmvUjNVj4c6
RmsMujMn0fSbskII/6e4f9xocmEobKCCiG1i+oUJcQtHeFk4h41p2p3a9gfVqYH9cIm4Pg3uCWu4
86POHGw6bRJnH+u2pvtS19iYtSJFXn9uXnvYsdPrNhWvaSuH6OuzdyG7Q+PMW8pRJC8/5cYp52NO
9RMZUOK7vt4FKLHOfdZIRMDb4l+NBPRpUtHPajvKAySaTB51sxAAWftHu4pmN128pLLpgXo5UHqw
4Sha3TdWM6qfTHvgaZ6yQNApsquPr57iVjp3shKGWnRZ0VZcQYs+aUlnT6gBrBuGZS8Fm0RnZLx2
YzQITDCDi6T0qyJmtkRqegJq/4RTTvns5Wa4C4soL3bhXmfWQHwk2u04cef6iFH0UUsuYOuwxEjT
fGzoH+N+IEoZqTxzqClFkIFY/BEWvyho4P6cSpPiqDp01wByteTKojd0yD7J87G784FOKlm+MXlI
ug5dwqe9uB0LbzaQhIzrYBfW9UsYaGM9jI21PJ8IFsOA7XCeBF2jivo1jPZs9DFlols5NGjX5J6R
64501ZuVvqat3AA1lw/qWpd4qSErfdM1+Xk5c/iRGPjZ7jk8jEvciK58nXmM03aVK3QnfGQ7T/vf
groqeIzkWHl+EIxHIHEhrVbykFpG8ry88mQ6327BsvQWY7rjZfcmc+yzNpG2kw+QVUi8Q4TgQKSP
GWhc8bhkatSs/l+tRz8nNE8iEPYJdS+5hhyfmAdzBXH3R7u/EAGb+e1vf9WUD1mq6DIdNxS8iz3J
P0PllS+JmizHLTtGJ2J74gwbkIW4cc+rzNIE558R5gZumM7ApB+MUgwLWXU63uCNJVAYy8pJs3s0
qiFoO8w2q69R+yOZlzCO6AiwbeTamA5J92mWLfRl4uxeRtLwvDmZW8YeqFDrCdc3xgztLfAESJa4
bf8Ls5NJiviENW3y3aQW+ttIc/AwPqF3ztz8+lV11bqLx8+qXmi53ub0ov5c4lZvwHeFrU0OMZGz
i3gOUJEw7QNlTBgSdFmqrFHRN2eRqMgh57T0MhQkm0gxBy7OzjO6XvIe1gSg4n0v8ankm7wL4wpY
fzY47OMSqkpjYNxStg8HkCKAParQ2CLfopID2JUuiOAwztlXBgwBaqFtS1QPW3BajRs0Qlt4XQLn
g78BAyy8kQFMf6e37AejDRZSa900icwycxPfuMl06DX4O0mCQg39m+MoL/ot4QUs2d1TEXDzDD45
mp0mNta2HQ6b4OQpFoBTL+LwbUdEEIXSTZj9ZZ+D+6KXkKgwyUcoUcpPQ2xyVwC0GrzTZ16JOax/
TZqaJ8I5f7XrNWUn8RB0rSZX4Jz58uAjmIXJt6AazcmaeW8SjX6nAqowiIfhx0rs1Q2QGcY1/GWu
XmMP864MkWqZgHBpzHGlnGrORBhDODNZuVp2TjnXlukbN8qq0VQqM/Wj8BilrubqEboeuE7j2hxp
WAkeAnxzEvTt18FJTk4UIubVHj8o3sisbMIPxtSG646SLQQ/Mv+dR2BoWQ5ceZm1tTQFklsCblsW
mihS/kea/4oTLk3ws9NWkXxvaoCrI8qYZdr0Et+JJmcqO3q5OH4H0T4j0/PQ+M/MidqZfsAUwUpg
BLDmpC7Uif0CPQ4J3fKaIacMc9nuqIq3sJkOd5twj97Gan+EwXSkBVvMXmD6R6vr/X35wmRxIvPo
EeP6WHFiX/HZyc0sICFSB/f0oTv9mwTtDBhjusdtI/ivwHddW2evVqx7Qzg9LkWjsBs3F8juRZz2
RdN6apf8VnC8g+S++rW/Jiq5RJX87bWH1vJ6G4r8NADo/tQ/svM0kz+P8vAfOcHjb2ngWrAuFdX6
nXVNbgbGXBTRAANuBWSLhk/AeqFYX47PFVreBovPAff/5ePNRgFoAbGb3khCIBnFYHgHbt+HQcmh
yAZCu9G50t7fQCflY9n85MK6iXWdbMD2kWFlGqKliJw9C6SpvkayzYM81ky4J2YkC/DmIEg43LjA
r2F69eO+KQ9HXUBgiy4OlJUpPSDNFSVXwR9Jn/wO1nk8h/3Ytey+J17fAu+Am3jOCfe2URcQvY+v
WVeVCC0lJOuzYofbujR3NjSoWcvIPFuhJzzw61BK2q4WdmfdRm4eFvBZT8iuh9ycTK/s4JZInNJb
jIg2lX0WmlKw9rK29S4ByzW50XBD/ttQpkJzamh0h0FxZsfWRrCXIhdVmJ/rXjd6PI08T7oXSb2F
f1ja3NySgV1shvi43W0Sfbbnu0G6l15CAmOR5i72soIG2sxjeOU+Paw8boRfYR2dikjrLoFD5j+P
OZBZk5B1r5Hnsr1bMlh5pBZFAlF3F9VMsG0yTrRPqaAEEN2wmO2suBWpW4I9bat2SVuR/KFwn4qa
+zhakCxo/JkFa/gMGq3xx5xS3OQmlnduPJzVE1JVo6Jndc9mywpUywwGCbBAyEol3Pck31ya4fWD
7uj3mUG/YaXaave5581/uC7tDgqsDxwvzerL0kqaW39oW9MOi9EsXliUoF8mDpta90N/yUUPbyq6
4t1Em0lTaYGLH8PO8upbkj74U0oH1v2kWmqYLcv0LFvY2yMlK2tI6bzT4tgvk3OjozGjW3Ljy6d7
8H2o5D7Dffqiaz1NhbEOsfkyYh2S3qptQi6tLx5ol2tRe49GQs1mr5fXVsV0MrodsYKrNLDFhpzn
9rTT9R3xounNYT0CZaosrArAOcV+9xSNBg3WJ0OXdpKEjL4+OcE/crGiYZJDiXmFTYXcZRZ3HcHB
nQPG38l6yO2KRlLPFbf6ZbIQFjdytdPk4nlv0eAF4hMBTxWM4U+tH6uQ97JRTpAcFKAqxQOGUwUo
mYljVkDv8BOXeRj46qV6TQwojXGIm+m9O+gpIJRd7CRF4wHoqAKhCrJwTWFBf3/I8TjvTAtR8Ld5
NeuElDDreVCRytH2ano2D1HtGpDeq8UiUjv+7D3SZMm/meoiGgD6UfO/Ow9nO0mugPTFUzxIiQbq
I6fD3zBuk/9sA2grFSbS5wEnjGYN2xAYfsSFpOZm3GyUIhWcEwbM/p4UKczuNguSYqd1ZHfCu9A8
Owj/zCFsIZzd9Zjs1bjQD81b0xsbXGv1eZtQlhxUL3F6Jv1wXa1pDtGNI2/M+17+LKUreATypQxz
vUpIe3nDH/9Pcuh6XiXjegoZEqjFpoH8Z3/ShjNrsqvsKz3rsj2ce5g9wS6awJ3MnRATF3H5OK1J
2aNCO5tSSeLKJlRSP89LFvkEuY2oSI/r14phoSte3obiDpHSWc80ZK7hSo/D/Jh0JUGKT7UjmXkC
ypSO1ye40yYVIdysxQioUrt3zdJT4AsCQoo2ZSy+qrIBYtQsJMyT7r73bX5oStSrj49mnxBZNICD
OGjrYPSl+wQBGUc9DWGlqZv8lBu2TCMYqtPySfkpm4sEi8bjSNcxqR2TVDc80UHhazmmk+8GNgKB
zY2toEgxULnAiJCufYyDRC6tjPxJ9sLv1J8EMdPC4fyBVNM8xcA8O9DDFbdxAsI38IBxYYkH2dGQ
h+5+LJN29GvJPotKd1YJZ67jgfJ1oJvZoYxVvJ9iYJs3x+BmjywZXNZq9dhOrb/nUqrdLoB79piG
0ylJ9P9cQXoWgSfCp0qeNpZ7yvxqlXlaEIkjUtBbdxFw7xD+srzryw3GQupXdZXE7y+u0IPfsOhy
S/Lpq3CnSDVbiIQXc6Oh0mlHf4bIZhMkuW2iRWsF3Xbd4/o47GH7MT2+lsK+k4RBkFSzV0awkkh+
l6qwsASNOiVEvWvE6SckpT6GwR3bKSczaQS+sslaQPo4T0LCyNoiuRVwDJPUCPlhQhHGyciuH7oq
hditk+9fjlz5fnjzoqRkUYC4ULvqd0t9P/+btxcmFLrwm1PqB3nhYBlae8C+4f3axA7YAqFFzC0G
tQ26Nkl02th52GcN5JCA4MsRiHXtDzLsu6ZYTLbdEcYeNMwPpuYClfFxgEx4rNsCtI+cgUHYYcfZ
DUQcDFN4wvkQFvJQF/JmLFKTrSulh3W7NoVTZS6TFxxCvAz25CqhUO55i96lMoH7GnF6wLzHcFfT
hfxz4908oeP3KnyY3vCg5AeDUBfD40AXEF/RLi9fq/hKWZm+xKyNHAe06TV2vtqhdg2ietXY3wj4
hRYT9CLSZtYWI2YRCCQ66diU8eg46CA3CRGrqKwZAgU2hCXRLSZbAWFbNaQ4rm2PtmPLg967QrsJ
H5Jsr8r8hQ+iKh1ua2Qy8KvuEL1gJGvSO6UoByo7CQDFnVLLa5WMmyznxDU1wMxRCOozVIpBW5LE
rWBGaMYp/mnms8s9YEJK03hOkRE9X+jMI6gsddNUuLlkqN4iOIqUxCN2wIjCtIF1bDaySBVHsAj3
p+8y41vcEBrRApZnUgTWP6Q8ej0A0iwYGfbGrt7LCgK5s0aJ9MW/q1FbARdceQ0Tb2TsH+O75g/g
UC5GSg1n/HbMcG1VDzgBycR/wt/x+CgXqY+++rjVn9i8ggrmzje7yeDFAgJ91FChb93ZiVFBEBp6
JkWbLXmHTgjCYIcYgBhkjEJ38FjTOLOGWwOxcTj+imBQYwiW9BocBK7N4NldBJ/MaKRjnbRCIpRh
mcCSwAmyUeUamebQXNyk/1oEIId7OOWWOxuVSql+wDv8UZkYdIXx8sxW/u17qihjSqWXRbXFVUJF
yWIzZSMfwBwEdFbzY7u2XNJ5Ta3sDoq6UOQFIoNziaqSkGCgfvN+X4GYQ+0l4sJelw3GpesUQ/4W
j5HXPQkIxg4gto0xlqHOyCjlpHUqKtkKXguqMT99hN0IYljuOz80uuCCzN9lJ+l+kNpxcNnqPIEY
r1Y740tKPQQbdEuXFibo1s+J9pykpZIH1Q7Wy8O5JU8mDlwTfkfg5mUIRnbQNzNWKtOyAutomXYr
l9/+xi3FFa8P+1jYWn46sVyhdklKhK+qNnPKVu9bEW7tjRfJMAdeTxQnTf4mwehY+bXO+Vu4smK5
wvJNX5mZ3maWhXfdaZnOJgQopVwUFzupCvx3MGeGwMdO4wV9atzT+t9QynuG1sxYuTKx8aKNrACo
Ojcy6rKScmZ94rRV8z2bvccyiAbngzuc1Ax6GqglhKFFjFQq7JuJ3pWeqQWebxuExFQTeN/uVCCW
soNpP0uBELvgLNVbqpqRXSmaztrOdBy+Qjw1jF1oHaRNL/BfLXXt2drGDNcEoiLeGlPiUwPnGbQu
RDKxnj8t2PAS95YoRD1YkTJN2hsjq0jpxVWlQCKQchX23rTE871ZUSMPoRWwWQH0cHP2OQhzLUZM
jftgb/1+V5rxZeeuHiqkN+BwSHj9YdrgBSOAlXgaacdNtTHRPdP7uqkXuxVtTvPuybPkZ5EMPUyk
xruAVfJE+XQYl/9lfEKQ4dQ4st8TmuzvHRwKAx56coZPrUM0nLd0RTzp0dUzf8atT8hK3/MF3Jh8
+he+JcbNVNxDGdVzEzMdLikBgXybR0C8z1UNKXCg7gqk+j7x5710KQmiPgzdF9o6qBD55L2uLD/H
uYYIAIo4a0xCuAorgGDhgeU7vKSSmcbdnU85U7oIQxbG0q1LYA3Em3JVUvaFP68AWXxaxsedEatG
oJ2jsAf+vzxYEVKGj8rH09kZrVrfFu8xWckbyARNLpq5V4NjyIbXm3JyXgRB2j4LsSVAyFK4+ACx
67TPH8Y+CUjYVl2U4nl7vXanLh22G8Ki8qrH79OyHCbEVDVCID5bMXu3tjxOfS++PdbOSn4kZcIy
7UKQQsWHvYln1liWNiNRZWLV13XWF446nL10H7E7X5gtzNYV0vxr3034sV9hS7foKHnAfiiHBd5G
JL9rUNh9mr9CLFlgU9B4qJeHOKHccF8Rcb9CWuG10jT2ctxORpD99YwWWiSYyMZEZN2ZJKaPQzcV
CFRMcsT8ykyYqSv2ZyK1w68YeiZIaEt6btmUfqLDcknZX2mz9RS1zy8TMpDk7CMnbNnC/Vsa9R4A
CDlFEOMPEa9tRvaFk1VCq7GWWa5bzFio/mlbtT1kgac9B0N/DLQ9f0BkwOTAuEhyrNP3yqHOOHR3
Cq7yI3xWi2rS1+4vbAletq2NOw5WQzUhGDfjXGu4K/xTqJZceZwtI/npSCIy6sZhyiGRa/YKRpiL
bW/oeHIva34yeCRA1qcnqgzDxfgSQ9fXe+RslhX68nMnV+a4QyQlTfzLzWMQvu0wRdLAuJZv8Hxa
PoLtk37Hs3IOhf98WpmE3s8DNrRUlFc+jTxUZp83ySmSRybC3MAqsbgUxmNnCNB4/Rw94v8LLC7M
O7suLAX0ckhwx4R0H98uEkRV37xTldIC2mQ7e2hichvLB8xqM/Loght7vu+Gq2Q0QH3uT6/6HLJD
iMpYi8JhR9JWbnXU9IaDUk9BIZPooYNUUmPmW0+FROMP+71GmsY+VuuGzl0PZBOZY+5Vk6WpdBBA
QK92VT258fmuITFrVURJpA+PlX5jnSGKBCjJS2Ug25lOZyzfyCLJqUulvEYqX4Y8e3/T75aAIxXe
UdaTMqEBo6Ql5CR1VgdMu+zkQhLcxzZB6DKSQh19rIpq16qzaGsbDLdG1iL8iQgUg9KPprPiXbXN
Y4FCiIuHz4LkfZ18x074JQh6PTbXLNbbfvpzRZvlBMYcbp/fFOuPgHR8vssoXY4f/zmj8F+iaBXr
Bh54wsePiCJ3pIZPPUHLwbL1Fd7/4li36eRYM0GeMDyycs4Z7KMvlOnefOxf4SbXPVsenAftQu13
q+SK/GILWrseg3e80aj8Sjcb4+OjvntW2ObChC0Nn1ZIbm+4xedL+qtRtOL1k4VDsrcSrDIqORfS
lekLU/iuI9NYkCIuweSy5pyek+B0vY+0f2jNJO63vQtFSHhhOVoc/V22SI2qTKB1nwzaLTyr5hAj
Okxk47tgAeIOyHxVnYW6QVhMMARfglwwW5U5APFfHNTERCBVTBxI20Z76YOSB8LmQ1tVKO7C1y23
OuRbOf48i9VrJQQVd+UEz0eVgwVcnhggMYXW8fLWuCwI+92qf2sZT20/6CWFi+lgbbK7bFSUM1CP
xltLeo8kVGMS/iV3imWZpnUsxe5kQEoQWeJfZlRJPycBs5E27yBf2D7ubFR2udDDhwG328XUH/pZ
h2UpAHj/iKboGsBi00wFqOS0P568wCMCNhXrthXFmZqnGrG6zA5aaOs+3uGK7ee+PzXkeH4FE3vJ
aWbjK2tOiguQbBrFZE2zDs8T0/KfQSPQ0TSFDiDYf5twZbhWz48l0ZfzOzLY3q/P0lhqZcz9WJWm
kWZYRQhHURnF9ORXDq/fMiUK+JmTqsIVUZ35FclqE4znGlB0dTXtommlslMCCq5G1k4RA6wjJ/Lk
MRDdKPith6/2LkJvETiZzne3W3pfXgHm1Ku3z93otcBYnphYU4a6BVe6yztmP/f+ZeAT5E6TNmYv
koJI8l9LqbTCCZI1UyLm3NeSNe0pY5uKLZIknJW50U09O/ETgfEQAXMPQ1cV9XYDtFivcF4Z+CEv
GuJk3FphsrLUQPX9CIiK9a2jZvp4t3jSu0xA7aawYI5PxF1DaUIgxdFHX48f3zll2aBjGebJ3m3+
7mkmzkFtI+w71zYmHXiTw+EEBYlBXR1vEzyeW93dfS5Ye3YHRznsgg/5/6uqq2P18GtHl0A3gAYz
ivJjvPnywSO3aJfDDPiQneMvMaCwupHC0/Uedn+2+5Xs7RCNcwyTLPN/Tp+4B4U+TF/hItJY8slq
HbUepd4+k3Bl1/dSBi1BAH55vufbEE5gduM10voOepUi4TLivwJOTE35ekzOvP343Inyf5hxp9co
QWqivT5EbglYQ4iivK9i0s5Hnd+fVJ73LaSSfDjrOhLRBtZRB9mVhucFpFmc8fy7ib0nsO4HM4C4
OosrYO86JKzHYhurqcJ2oFEmH6ZKtU5m9xbUKK++CQSrOTIjc3ooxRj9v81YDkXORBlECcxTnG83
qupr3CIu6EqL1qPjEAUaZuQ1x0FbR8FjFpB9e9xIWg8URW3RY4DEQLfOYlUeo4nCp7hCRxvsjxq1
CZqi5GRi3BEKnEEF7LTwm0omHu2x+j+/SNuCnjwMuZz3djV3gA6qMW/pQ1fR0SqjH4ldKXFRtOXk
MYhgBItj5oS24wnDGosn7YKPVJ6R4iOiJOXkozi2u2TFxpesqTwDR/CTRljMLhZLToTMt1yEnNr4
tYDNpHipAZ1K+GS0pp36EgpOThK7zXzfSt24Ru+J2FMgTk2/cnaJT6MnVd38mKvqHrgBxCY2xnVd
EG4xbn1Ty/DAEOavHz5/P9h22lHoNRX22XWa6ql0/ju+sG7oyWqHbUkKSdODaV79+lYIsacuBEgy
Yr4+zgPE4RiMEzN0S56BFuVSJR1OkvwbmcwPh3rh9nOKlZ+kCV4i9reGvRgO7088ZvcdTl6sdxki
Wit/y/MJafLIqp7mK4hjAivMZKxzseVPH/bKr/VBV6GHH1RvpbTzW3+RBv21XlY9ITbK4gJklQCA
sqxjq+XW+RIVrtSWIO17gX3bd+E5XA7e57kSsSrfebmsJTpLjDjVb7Xn61YjhzdW77lEJQ93hMVJ
vwYt9hUOAMqcZf43RZ9lkARzc/jGqmzhKOkb2ginJhVX9tCzF8UWQGqTVEwupS2JhsETB3xP41JA
QXcRL41KXdn4Sc9QuCJsyal8cnXSIsUzykMJg/KJ6yUXWCt8SA/ULXfCqLedzscFJOv588UOqPdt
Jfhtw+W01QmTnqNVDdkldm2yftUJo2z+5/mjlSM31PgKLNqVY+n9nB8khBBh1AE7bk9IRJpSx0r3
ZKIPsQiX1D5FjHi7ZPEjb0TYSqfhlB0SNnN6aJvDAUbh3QSF2X1of/aJ2jplhLdcxawYUdtV26/H
4kDYu18N3k+hV4vIHPCpzntmrhPHK/0WFjWBVo2VrY+uODam7bQuR+XkfdWsmjhTJsPYRHZsneFi
mKrvyxQoAG4tUehmx/pbXdexyvbs8UGlqx330TtHlUaZpDycjhfqbhJ96ms0T6fckEcO0xd+beOH
GKWOiKoEo855SbTvgeslhLRZPATU42Lbxa6/NSR3sBA6+EE3T4jlkI8AYFvo+QtK910PkGrJLVzg
1YVHvTIQzpXaT+g+0XfaWzN9roCAhyKeerpAQgn6bYnyQ4LH3ucPe8p4py67zg8vZU052fwFjpa6
aSUPi4p0gxvf20+YRgYEjgo8rdifU+nDss6OARIMja99MPkP7Cd0JNg5cy/7e1F4p4Y9Rc3WLWZ8
shO4hudUUEHiWnGqRmTAWHiNBBv6K/QP77EGXLeEVp8ie4iVyusjzNE133CE0h/dDipRBJzltfv8
yZjW8bjsXEmovPhdxidlokEnCgVfoD/TM6+WhBsKo2OQhSe6E4vHRrpaVyYdSvoHKEOBeW/lHwe4
g4RD5bl45Htl8YREWNkYu/jJ+cgukMnXiSv0H2YnYz9AIrCFIXxCDmvaKBgm0ho92wv8xHZAWDLy
T+nEzJzPrgX79FZT6hBM16JXEzKlDeig9aAenjAJiWNUnT+r7TCjJZvVeOeTgYrEpgJKSomVDTt/
7HE04uddo2yOtyPFeEI/Ql3LKkAN9KTJ1WEqmrypcC0G6q57OV4IfEXmhHqEZSUKqlOo9nBS3zj+
ETXjnimgkPI3vLDGW3DqBgsW+4bx+7IoWQ6P0iRa6ehmyfON6ZzsxiM4C1E8iuKQt3DdUMapPnv8
SeWSyRqBzUt3cQ0CKduiSbKk600L50zbmo8ZinTBOlqcUIvs+91fTFfQSrS6jiCM/xu34qTimvL5
PkBIn4j+LDPTo9Ce9mTnmEdxYlUYK1QbzhGxRdssFFbn0NxBih6b6O+lu8MVYzlpMDTKxuHwn0p/
q6KzTidAjSD1qMHLY+iuslcxu4bWDAD4V2JktZ/rqedn9p86hD00ZzKqgekYYpy1S0ggqNxbvC0y
GNnoFqjLrO30K5piFDNX2lGHJSYSTAVZ/hrDsTtcWjlhgqRZ7Dzl5ZF7wngTy4hfV7RCzVN8zGVA
sSZrq7GoI3uEcCJC4Bz/6hPkYCqCeYSseKPHTrmT3J4RSeX+q3U3/ClYuQtLgrETv/HtZwt3lDMq
kqFFLaS5mhfz4mTNVuSiTGIDNztSr4J7KYideeGJ1v29OLw2SYlgcMkByg6b68h5I95UDaG2bxkF
ro0l5Lo2R/G86lIUZg0riE2IwwjpvVOd02IF/gcp3DhAxbHSSBt6OPyzKUXniVkqP5BkLQ2eYmui
k5LPBCThHkRtyf9xvcVQx0Dj5M8/6HihVxA2PdzcAsd0aVHUG0oluOQi7bagByymgoFhVio138lr
/ZN26Ic2OsMabfnyityiuxVU4Rtbg6RlYpYM74syRtkZ8fcctdJUyBAR7tn//4drkiplJkZ1VbbW
6DEccFus4HUdGU19RzdjhAuhEicUkkYyA/CKa/ZaFkYkrZGKb4CyeEmgAs3EX3wzUjgxDj4/0J+U
gigW/1ndTjAcOw94P4kKdLfoeaxJJSbPhmpxM1+PDXE1n8zpQZ9Foup7z2oUvlzYU9Ac/MM7vA5U
n8zt1scBCBS1S3/KBHenq9TJY6vntjYXXabH1ye8+BWN8a5Ycs4pODUKNd26M3IZ17Yshu789Wjf
uN/24AQUyHy+BgSe/NuFj0z7sT3yg/TR3SOvHvbrNpAr63b5wN2AbHb5pmi9ZEuojg5OZ+hlXmE4
/WdtfVlzLGMneRwFjHJPRKlEVA6bVsuDSO11512ju6ToaJ2JD5pkJnvwdHDBxAouc4fNFudzYc4q
5tsQRO6D9DamuVRIl/jlAJGoEJQKNFEHxvZSyJcZAHRQuPgKl8ukkJU+Eb8GvuJjTVq7TIwm9CEm
0FnUJYUKkLZ4gg4QDbpyf16kxOaIKSOxFaxSwgLzrNK6Qi/w28ozujamfZWQxxDOCltN1TFVkUQX
6cGXh2+3qCIjPPFAh8r9nCGsvNL1wrKdmtWocN2xPm0Fitcm2SfHYmDxCD8UNwwHh49pPr1IG7bx
+Z9lsAUEjOxhnURwOSjSVdfxZZaDXxG/MMegbIXjeUhFCiDCqaQOrnjSzAaQsq/XHUuYkoVlia5H
KWwfZStOrWuU+4gaZLWNpEXlpZRWCEysRnbJslcP2DipTRlkGCoVKz4hW4LlAhbk3o62RSoeiNZx
3foDDi5eOyMRvzm+2yjwhVW9ZlH+g8kW0G6P51ZEEeH3M64Q931bFjSqryL1jG+5ot307RNEG4ia
Mu74Bay4pyiLoEY1yDAB2FDI0ThZz/K1PkPUNSo1C0HLPFrLMlRoK8c48HXxCbnnLGalAnwtIAbf
NhQLMwqXkV6blQLJW5nyIYBW4RAsUH3vEXzdp/YH/NTETFFsKy+oKwRn9wlvb9s+fijePbZsXPvV
/Q9Rxj/+GiSwpOphyVlUZBHBZ3sGQMhyGHqKTUKqprPv7WIeR2AQXnkXG5gp79fiiHo6Un2KtE3P
ygD4esolSduFogGRzfur3OK8dFhhEsNjZf3FS2/gxvE6KrsAmR4UtCFkP3HUfG2SiEPF4GSjYDiW
ynhj9V4nqeCjEL7MZb4bDWq8pepCuKxY38qbvyRsSkE8LfAbs7NorqJ+etHEZKhnx+8HOstISA4Y
/onqdQvMmtwFcyd+ksiRAWUciV0NI1Fxol58eJ+9QBXicRmXnbnHCVtSP1MZAWMo2y9T3ErPC6RX
/DbtzY/yYikVBUJQ4EncgE/mJap2wOfYmJlUvkn8NkN1t88znn2w7kJZ95sR2ThFQH+GjATOT9Pm
iK6rLvWCUB173l6TNL7Ni5mdoFjubqHi1Ug0mOzolXvXM7YSmCW/Qqzxn4TGan3cB4MtgsZ0KRtv
8BLoDFa2PZuvU/B5Eo84Ur0hGqAoMHbeabjEobnxGIVk7Jx7fiumDE+xXl2lShz39rT0Mlb3x1Nv
mwi+unppJG0reRgAIUIxbxDbuQyQ1yWmBlEbVJlAyT9Fw5na7slSiv1MJFXcjJGiVQmo9sXjZ9Tm
pVOZ+1tKZJFN1hJoTd15HFuCEifexojbQhEYkEtpZaoLgmW9ceUuzISsQMWNmFnnbPOe87nwf1CI
AQxjStyWfoV79uqGEYkSMcHCyGaC56IxCB0plh+4WB7it15D15nqoR7KWSuod06MxXtFh7ayxYJi
6zww0Wfem30pbuy4/6tC8tPgq1Sk/X4hRyQr4akS9eQO6Oh0q29ZOPnGSkjJ1NvyY9JV4hyJZZXk
rzeURC5jfGjOi/03w/4Zx7GRGrU1nFmEiNF7mOtUcuuoMfvLJ/WnC+mqHohsexOGEx1bGl65rNpF
W+yZADV9n+VUtaBLdXLMVobTKZ+DKfcgqjx5wpMwqxl/U3jAcBxpIBMpUPfXrfn4V8vHMcbTCNpS
OCm/aOl6x3xOXR+kAjfYK4BL4pE+PMU9lDu7ATEFqnLrEz4bONssqbAWpQL1Q1Pl4Sq5ii74DS6C
7q1ZGwuHsHK3MDkf6S5kj5iQH9eVEyvEqXIa+rntSh+kP90C5HSGzfOIihJBdkTgn0V14cRC8YX/
nhIUtQvoT2eyNAUFmVtUANreVxsQIT3/UrIpkaGLLdX4206YYQv+Xz7ee1F0olQzFe4H6GmyLWxH
pfz0RhbIVGpJZiekhJ53pqRW0cee8qxJuj/+zcVCsTsWvK+toYnCRGAmFXajxqrIHKlKymaoAdIE
2ejWinpiOnfiIt/SRHFYuTqB6eup/NruY2FQ23ZwIBT60IO5y2p80IBZ6Rfz/k3IKnabbcZavR+E
ZeQqLPv9Im3rdBLQ4saHfyL+eYm0gWi+3RqThf+gpltKB5F7mbUy2mAtWkzXQEOqOcLYcHQ5QYM6
dC8RaNZzfxGandAbiwa00kqEScn2LU22xD9+vTL4h+fqCgx8pl41nuP5vUqzPNCFD37W/Jh+D+bq
Ou4XASO8fJYhKXSTUE/Tkk2ov/fmt2cSqyxp6serb1pAcCFD99YMZdg8EoudBP+g+mV9Pa4Ukum4
ssI4z6ygCumHqsgFWuXIRhF7R/2WBj0t94RZfB38p5jb6DRl4bjg6GA/wwVs6vhL2zpx4QHZdstG
YPHeK5Kv/H4CxKYJylLadz/k9IHVoFu/QFD5HrvA9NkDMWLyY3aMQwXW9J8BvVFIxdSJeOl+W6zX
St1LEyQ83cylSwwPWcteDRP3dEIFTeK010zC+oy0wi9YDKGqS8ICVPJGJtzSQAkVpavVFrN5nMXC
MgpFL94+x4TLzhvNorG7kwXFpUOmgnCXmwqoSjNoVFPkoY4N44jrVs22r2G/wfliPWkmcDyUQx16
PXxKZSxy+W7M3kVrOqZL0hkYt1M882xzCi03NHMI4C+q2aqpmF/b7F8JHG3PtK9c030TRIb39Dr/
Hsv2+A/I9PjGhrr/GZT2G3PAtkzgCcgHw0BrUy8QpFHqWnT/JIhKrfhV62pbjdYQ0BrpzbF+tr1t
7ITIPo6eFV/UDFtBAk5S4cWNsLjfYKSgy0bfexrBPaujEQimrEXpbDLQRFgm5BLG2tIPUPSwgC4R
AsVDgBzdEcL0oqtJUptHJU4K51fWddBCMJOjuRlDHnFs9px8Gi4iapbtI1OEaIWoWsni2ayfFea0
cKkK1WhqIla/THawfcpK1xWtqlqTj9XFn3TMx1rXZfhho8pBVApvGbWHofGCdM6k7iy4PdXPitis
rrLXhPFF7/TFVKRRTXASJGMk7kcXX/LZ2RWUYG0AliOobx6VTgWPvXUI9AwZz8YUtyXJxyALjT0b
5jjuKi1PJWGRMMyfAzcLTIYJMbLchidoT8s2XHLArGqHKIiJ8tkYKIlQlvdnDSYOwjDcbew9hvX/
x4xLx89bQfx5CHQbDAeqBnYy5f8eF+g10RfH3Ykwly00rC9AzCNU84Dwsa1w8FcbdZSYo2NFsFdO
7bGAGEiRKVu9jUNMT/uSOP5MvsWtErXpYyyQzc6hlc52q2s00GHBsVXKIossN4bkhPwBbY2TjodJ
S39r8a59wtltrhDk2wDR7vrs3/JjKlWvku7inXdm2WmAQgs5qLMR/PPasrEeG6BBCS7kZq890syA
HvDVgFdNKxhcNMwe1UZjRtTgQcWy+qWokudo/Bkvsu0CkwUM6xPWQohKAKBQD4P0gyu4PBQoPJ9L
0zgm1DRQoSid4Ph2dRgkMv7nmlRSOQgP/bVUKGp09ZSWmzUn7TFdq8QJV9xTbPmgD2PhptP1MLac
foOOET0NSpeqEd/yGa36P02pqeuWE/TeBI44wMwDt8arNZHW2a6CmHMhD3EcE3VNBul6WKMzt8XB
wj14QcgpEVgANzIlwyjxOZn8nOwtrcu3qDTFKFP1iay4D3XOwptD3ysdefkSlkBiEC4Ez/TzZVxA
3lb/vAEleQSmFazn7jjn1NSSA/TMpWb6u9bSBHFAZAxbrG5rBTqhBUdTPDNMXQ6LmkCexpEq7UL4
BCb8WuHo1coWo6eKM07SOdubGJ7+y3hHymVXUn4PUacB70p/bArrV3UNKd5260u+4Xk/xMdJGZM8
kv+ujcMlkCdKpQ6UN0/GTfb4OCSQznJGY4UUylZDG+L8U3XyXWB++nJQ1Z0v50ll5ryOwJVP77J/
MIfjaNtCCjLFV+uSVD1In1o4UVwCzs0aQ/Kiq+pT2+FX6c4cIK1cVCGWpCmXjhMPvABRN0tprlCZ
FmKkQ2CEyA95nNuMWeV+rfGdUyxx0ToO0MEqlFBLy/Y5AhPpPPxLqb9mtzL1M4d20OBY/ZjeDEHJ
SONfzoWvbsU4kefQRzquT4m3a0txZRCHcjKLL5quRCqgRPSAdIN9d/N87yAHiJREZdeC8+JQuDQu
uy6IPa+PPe5gDhK+xdJW2kJwGPQo4Df7O3DE7XETxM53qAXijVHfnwwOY03FrmNO/OYZ9+/7i2Nk
V0uZOlXhWIpBeF1+i4Js5H5hhfjoW32/WVwzpmGe9aqMW2fxdXPH6+9efDBHhTXEPt6ewNd/hn3h
IH9lRzC853/cbV+SU2kXhSewwB3udJ+mHgPtIeIvdwj8DlxEW+GgbHZSWERrJA7SsIJnNxp3bgjH
C7tp7n8PxpDd4hoQ6EvF4h0VKhmCUUQKyTaFg9tAAWpnbYE8GOdpEezlB2PE/Ie+u0VCouBkOfKB
qBoE9zZWYt9d270QiW2Un8M2LSJPLr7vgyWKoxGNFZ+jW4Myu76fUYwHSJ5m0Ps3pVT+rxSHccQk
t70kgbOLCzSKtr2m2o0Pt+5w6qTph1y/nMaePMAdelw8f/tHJNvsDdaCH7m6V1QTO8c+UJk5Sa3a
n9+8v6LZ4mCdxfvrlhqZxj1f3ORO+319iC4pJAKL5Dfs98aggLG+ihSnNqPfcZueflqdeacokpNs
JUiWUihwhRsJEsn4ekN+Zn6DpUil2Aw+V9j/zt/pB7GQMXmyrCf1QkK4a41REhZozPXVLwvtPRsy
tJs37Fek/rWNFsxkr3UTTO5wubNpNHONl9B/sqTRCq8rrMj3cwifvnBLvAD2nqSKE6EfkA5p0Rym
V2mBrruMNL2RqY6Ou3it9qsM1VhvXQZw4HP3xFx3AGrk6fffzUl6/eZMThRu9bW9QXxIOSWAqzQi
8YbBLxvG5cGCrLWsC5+98EpdFsPFoqe6aRjdRqPOuM6KeECUog4Kz0UilV2TnykoNt4f9yNCRCOg
XRg0JRJ71NjgR8cxWeF64MIg53lTcdUp/ZE8QbZYDot19k4KcWVNRXXZ07B159Y+TKIKLx/oNqti
6fbTmko0RluNIHE5RM9PncY90yVIvrhK3JsVuMrzzfOZ/a448LzUAaZbTf63Pox9KHOOKqK0y3Mk
lH4EUweppKIMFMe1WOr5xXlbnyMNMxRVg0HyuMG+krH3Pa7gbCsd/Tq/VSFc783AjCkIDWDoljNJ
LXElDwwcDE/Ok3bEXodfYUxQAGbkW5sJGMUhAdo9jG5ieMVTSq6aZtuZQ1woUFFAh5O/e82FFOek
6hqt3x3JDyM0pNMBeD/jtgrZjHP6t2S2ICc1Hh1p7hEt7fihCQuzCNmVbRBEWsy7qsHDtKt2NyNI
v7liBXHxaF5Y+gCSQrMrodPWMdOyWOM580eIWX3b0OiD4hrGmV/wpOp9Z2dFEZaJanEDEXMUsnxU
qjwdvA6ugJM35H9WaM7d4PXOAs1N5+9ncBp43APME9OEBiFPyu2mIjwtv3/2CTcMLi3S2mcEEWFM
qEQwYtCS7GBmyEU29kgfe3xi9exWgiBSVJ5KTFG3PeJ8TsXkg3DjoIzKj5b9OeE6ZP2MZeRj5XGd
gIMAYOvYtQgCRLoFRFRLyKuzdq8WmzRjE/nqcN4sI8Ac4k2DxrWmnujl47JfH7b5oK546YlVRnI/
FEqpnnI+XeNz++x70sAFSIxEbKu0pbz3/ZDr875ZBdMsh4mKSET+M4mdhHBbZPIFP/+sdr88IdA7
dLlIuaTQIW0JFUHP9vmFLQJqVswgIsz7JCeAuya4rdV8qI9R69tRq6m346yoTTjd2JQEmiYF5HBR
CKx+xwpiiYCyNR20HIMqxQjUv2bhvVzb1pH3U23ZXLk+6LBj95dBUAc7QW3kP/oUay5dL+32S2gs
LDaZMzPTBz6pJnR0c2UFd3iQ/HhiNgpRNMpAHz/O2htr9gWSYy6Tx1E3MVQCD/FjGEfcu3+uYUQ4
NVyEWSH0esvNu4ybPy4mNQjcCr792SAfQbireP487gBrdPLzEahe1mw8ShAkbf9wOQntvN4Vt/mL
9C4oj9Xo1cMbEq/PRMphe9KJbbBSxJWzY2y6YJ+hu7IvjaQPXLkfxhY+wIOcNE/Zkj+HlWjFgyUm
l2PAqUluC0+aC1ByrTp2RyNVo/r8cbjkL1H6fq97auUndOe9EuADBxwb6VdEhMNopadEgc0Qukym
OUJwYu8PO5Yj/cGkNSUbBJfZMa8hQx8oJCFlOBvi/OJZ9HVMvAyLa05cAMVe3q+YKFUkor8iekQL
rPh8mCdrjEedEADhdXyHO9jKNSTef7PeAEQ3cYuCJx0cOUuHwVLX7Zg48GVoxZQbRollHkZN2ZUD
ceHDKWHr7oStYC8e6VuI61cMnDohggBBaoqwz/JzJXGQpnm11Wj5T7c4GVtuMUiTmampKsUjgMSv
xcyknoT0WKwPJStvG8roFNffnBtMyX8H/gpyGoFhcfqgC4xsmQOAv5tVbLEbhmncAHg615gamt7M
hc2Y928t0DpCrBGuuusRFn4w7M9jJOwd/yroDBz+TSst+Dordsq+/SmAC/hjfxM2v8HrOXw153h7
trm1nq97QoxgakyVt8wi6u7ltGySP0lza3MQXvzsWmCFJKY6jygqz1omZOyo2UVPSIC3f8UE+nV8
aaYEL8l/LjqJdiUUVyCAeOrtvACwUAl42Llp1DTask3+aVaUK/U6VIJfcAiQR+jbQTKC2bTifPRP
KVP//MepjOHoeLPNPNiz8idHXOu0LYxEJe6QMMZ7RZjkawlJsCEETLRu2jB41icDFjisyf2ieH44
mKjac+ZEDf5pdU1Ox0uf2+QMDy9u6K8hnX7bixOCL62+GE+2i+bW/deZwMZfn6OoJ6O5dZnUYoFS
O8YuHeJ/L9ci7oYw11FrAJXiJ05G3MLRjXqlh4Hk9wbzZMkLqiq5KJBkFHzqB73amgtW+7DCQPtB
axK6TDFmiTvKPb/8+t+3npcRa2xqeVXN1pNq7nSs0hJFz3h3vlZGxmE5wtF53HNMS8IJfIx49uPO
J5tAYLTeuSbT0dcUWYQwAA2YgNIbAvpNlCIjqkzjLJXE8PnDSt6+ZucoV9XPX0UUIvujDiAt9gSS
YY37Yl0zncOzA6d0d5VyV7ldZAE/E5/sbqynlsH2Vv5tTcLTaJr0S64M2jGLST3ZrAbroGMeYbsA
6HB13tWiOgUMO3K72QcORRr1yDcdEm9jplHZ/TSUawwCQHnOWhSDLlcH9jA6wOsNNSaJCfQAHSue
bu3wXEEpoDKDoJurplC99vZ6SmzNZbBZmTxnR6uPB9dec5ng3HlU2mOJVYAmbaHRbbWM8qRrmgOp
+R0iEmAvSyUzAukzNv076nwNPQ4L33govwLmWdgsfe3xcvHmJyYxFSvg2GrZvMhOwubvuSppcbt9
wEIsiSHE04mo9O+eaSPY/thARPPKi4eY5NyvgOfTg3ontF4Jha7DzuC5nFxSYaKvR1QHBd1lfUUn
dh09el06aUESqwaSTwR9q6cNvrWFSM3YJkB0xpmJg2bq1hd8gKiRs3xHcg6uZlIj7NtWiEZKiwrC
+AQH/jQv06LSW0vx4AI9qf9Lo4f/kBujSjAfUVp2vR9qvwx/zkvtsYXbUY4PcdwEF+wfkZEsXMXZ
KtKQKEStRoGevkgzEHpwybh70ArUiaGrmaCr8bXy2KwS9xz8zkWHO7I/+np9Wl1K6losGVA/fEoY
324EgKSCpG77ebMOC1GAtAOISSg1VyZIPKrPbBjSY9fj/zlrnMiX1RpcFTu2A9vPnGwYcvDqsD35
jlFSM8knEUyXMXupfugP96fxPF3I68qe6yL2x2Cv8PEvH4mH0VHbRx48A8QLSB8261GCN7AQHlGA
ngUGeCg86tdjV9pAdlOjpUZeQv0PG70ClNeis5cTRavccXPj4mcUC1V5+MLmqwE3u6N+d7+547EW
6NTwevx1QVtuEEZhHbraDBQKR/x5TrrrP735D6jLppgpWdeafg5PBI2Z7HCpEkUzYolkAn2RPDX0
n5WOekLt5de66Jpl2cScF4w5C/XskcuGROdtNVRNWNoHbiL2cGr5Kvi/CtWv6f625GqRWdHGaHHi
MiOA8bzCth5Ma0eVysSq46lIuHw6DOz6bGwd4FDTGK4gRPvRkejRTHQTIum4ZtuexfpaBq4tHsxg
nIKe/xoqlI+a/kB34eu3NpRcsgR/I+RZMSAvAC3wdBlUUB8wvpEV2TaFYD2h80sMTO1a/G6zlI/h
96N6qR0e8tz6eGHcNN9VlGMIdrrw9VXpljZLHzW9y5JxGG0LXyrB/x9Of3gyWjHWBWudALga3fV9
EwyZEdZ4ds+1P1YT0D0VVNEp52GzVuMAlXClQGj9G55adPXDH0dcyJV916nx+k4EJkdvrPv1IX6f
Dh3d7xm/gexIiC4Ts+GSrpQOHYlKtzz45K5phH2vb5xLtCjQblA93edXlWH2FGY2dLRxKqVKeqpD
kb7/jYFj/vB+wcawy8Y+LFbInMJwD6D6BWv46c70WQSZDpCQcVsjdIIt4xwIyiXAWOy4e4ZROwSA
Fftlu7O5oiocY3afxl7jCblELTm16JYP3UtRSdHfW1TAuS6DaRUiU0j4gmg7jm3IeB00VWu8NoM3
IU+I89T5c9Ke2SY6ZUHNFWFwjVMsJUDIj4sPPRNta7aQl8qjZ+92rs8h0dpbx3oFiHjqIKtvNejG
0z+sUZa1A9gBy32f2OW4t9L5AcSQN4ThVRQeAURmqluV0sFMCKf68icVOybegK/h5uaYNClN4Eqf
itPJXT6GzAqj0LLDbbkUZJpXSj4f46A0r+E+CbHS0KwWruYssbQHKrGXvC484mzpPdgoCJHd0Tq0
q2dbHP2YP8rfdnrPElAzuN0qgSg1hEUZFIcxDm9K8tJi8+x50uQfY5H2hrPkA008chVr9BIxlUpi
JgvXly8KUUu4By3wKiyo5TwGGx3hyb5Gy4o+ycfHd1wXdyNeV5XvNc53xGOvL5PAgSu9gnBXsf4Q
7El2o7LBm/VzUZAOMh4wVPMBpgeam/qx9+ZNmi5y69JMONrJA8uOxNO1j7r7vbzLuvpAWiOXQQLX
r+4uUDOyOZ2wyvi5X2Q29fLJKk3DoPnW9kKk+eD2cPqDCB6GEijOJ/5cuA+pDcg0Q60ovhHTO3Vz
Go2aTWKHHibSBy5p9/+G+wF2yKJE0bJ+SWYEYKc6bYS5CvOQDoqXQwCDy9n+Qmn7LXIYynpMPr6v
Pgimkh/nhV5FnIr+TDep5PBA/KQ8Ih6/VwstnN1VmO/gpAONd6KzlRP4C7sUfZVPeA+kY4xLSIqe
KPpHsIAE+agFimjCMo4r3HVTShbU9pXn97BSz6w6mcUBXajKSpZMGdImlSO4KDeO6wfU2pf0gEM+
V0ZUTtJxOx0pGQTMO6Y/WiAZeEabyGa4V6SKRbY37lv7sjANICSR3Mi4HE7zJGPBx5C6uWyw+AKW
PWuwtTx5sTQwIopwA2zug6d9mHXMT7CZEig4Dc2mN07/wk/veWtcNCPcgvy29XqUApwP3mUEVcX+
GPoyXt3GsJAPGo61lmHi23sed4zWecPIoaqCOJ4hQkX+Vuw3CVOaQOdXtezejqwzBTnA6op7AfNY
0xdrB0ij9dYK2ZNZOxW041T6itcPGCPM6dY1YasU5lzJ7RMkXWkfIgWI6VnI+UArH/t1QF5JbHxI
egyz2btKY+abftgv42DYdAdhKMFzlAmh+bxxtW3BLGzyCTj6BiMAjq3jUCrqxpWpblCbOaQ39KXK
4jhG67hZYS3G6mghIAMzzATgdq2VFY2MvJyH/XuW25VSCG+wQn/rZMR6Deuy+rOQWwYeY1diGMIz
8d4iQaY4HVT5ie8Lm6vAT+Nf+kIWH5nU3+mUMEI2OOSrIlR934oRRfznD0+nHoMjfR15cQ4WzJKa
TjBfE9VANPktS5zf+3511pkMfXQWcsa3EbZ9/QSzXAnMI3rdA+e1bvLzHELav6pcL+borjh5kfPU
icw8TWT08Ac0Fd+VwW37W4Gb/YbLQkkxDI5XcuFAHIv0LwQNN2fVwalcedRG7fGWDfVt+LRCnwJT
W0pn+RqIJ4ttEOM8G4uZyGqzy0ewuXcEOznC3Iw4YbBqwe16RKEIKfSNs2u2yvvEhll8iCmc9Mwr
lqqcHsUpsNdOoZsnuOrTY6yNdOgw9euXPvIoIgF6v7CKR4+W7PmVxtv5yn0iIaRDMbx20KyDgpFo
htEBbjIGrRSK3fup+qC8qAQyHsjKEJuUg96yj61m6sJlDq5dKV1SM1vG+k4KG6LA4PMxD74oOOI4
d3oNnPmk/o+CcvNKWEBFOgT/zoL3XzuW4Wt2Sm6aK4qcBgXKs8pXf3afh1W79O6+YyWpEBmRKcvg
n8MCA8vSZoQ7SVt7iE03UuutINTVwuyU4MKkdUYYcMBwo5iIdI6jJv2JWR1L7ku7wrSxiCuTZXnD
nZr0oATJTJnNAAj3PvtCx5RzYz6hJy03+3zmph5IleW2/kLpsucSoZOWA0nX+YaC4CMS3MiyRdNX
fzO92Wb46/A26MBIU4Y/TmHDWKBuTpo05VPcOF5ZZ7Bcpdcl46lLG3E3g5VJyZiZ5o9Yg6lxsnd1
bFXYbAR9oWKziJ+3ToWfZykmQglq2Gmq+XtHWjm7Fh77trM5SGqeUggZY7F1qfOGWSxJ/LuXFNDr
g5Qjf1MC8nAF4g9qASN6EVDW1cdneN4ErqeqzORiSHYgFq3S/uWrTr32W8p80LaGgtbGhUostSMB
gVv8iHT2056QudUfKvS0/CZFOJaxkoEGgaYbciPydwZtORq/mxxLZ9O9EruhNn52vbQDTZC1SpaO
yciyBEfSFF+EKEmnMW5aUHY3jYsdDEJzmP1XkD09cVOJTzGmNl1CCpLPquMJbwgBCHZXg9KpR+z5
MtEr6B+tXhlS82rX0CdbLaW9vds8RkluNdSVZc7QdaOJ1lnsTceN5504jyCjWHDQqVdGr5u+6cig
bLspKXXeigS7sjGk078fcFL3vDh9kluLCVdclh7SAVf4nClE7TkXhFHNkXZIl6cK2Whr60ufwzXq
H7k3md44ytcec3WvShXYXAWd9yFskenL5i+1UE2I0cHxci6eIzUF0FQBlcwZ92nZ+m7PJf01OrH0
Q9mx5ECjnme/ADtNDrsD+pxsDni5acQy8vWrIBTBDEuNdET0n2qmvuJeAfuixjvA44w/xaKaFUvC
rNiUEACiYnavrhNFiLrpYvUBko8CwfBCrp/8fXpn1KX+EH6ZP7T3Az1kX5XIeN3NY0KZ/dTj9Lj1
m7JxffxzyaO6wVcAqEUx1soxiDtTX9Vl563Rb0hqlhhYMjuNAz2XsTQINGKjHwV/PMImlHv0q8nK
18XiPsLl+7ODeNuhyFDQ1qXLlM7mhFVguozthezjGdRxX9KSDJxxmvjQ7KjRCtC+p3v1ZJ7e8MzS
IXTbA7c3NJRUXbfZbQ93e7Bgv8yvZliHB+ZRi7oD/rLppqmD+zH9y7liSI1kJecyZK71I8Jf+gKZ
vvZTAnvy6hyAZISHgDzSzVsuHe5zGMP6Rp5op6ABoGcEnCMaLuKpHWE8AlRHyT7eS4/k78zC8+K7
l087nsh0tWPYUs7fVT38bvNHlD/PpRPn1+/28sM6TDQgajWtjPWOUM/9D0ZCapEzZ5Kzy7WbpPJY
pvjg8kucjkVivQQ2zYKvVcTSH4gCUI+xTygPhF4gAhKQE/GVYuJomIKYj7zkiZdNgubkBa2vYJTf
OFkRp+8FqkcEPx5jDWHBR6DW7mvzbG8EhxLiAynie3gL9xo2FirNroWIFtUus+usG2hmOHffW43B
mNGKKNFBYSDtrHb1X59BMSucjdywl6HgdKkVjN9pyfj9e94WgoKo3Sh6VjpR/kk/MQtDTbxcbO+2
PIEURk9dTgtzUAQEOnclm9aOAjadpaqKGHu2WFCfZXrr2fqL/SceJ5j3R5ghdv+ABssBiQFhWcYB
loUDLf4PbXwNikiKaXE9BN/jQ09WmlF/pGbDRYVj1V9tJG0llN/6RboH32RyQdTENyy5RgpL5bul
fHeUN79QpJ+x2xfeCnK6diOWqiT1zUXJROsn8Rq0pbx74CIYrPNpNQI7PFRHLZTm2O+g0/4WvWg9
ap/2q5P37A3G5TWIP24PD97w0664ZWsM0tM3YH5I+13kZ+X4tb9GhOPIekUWlWDlNIb6sH7dAFwC
lbXjJUFelNVB6RcZs3aXb4ORwnDwfvxPe4P8Qh02eMUPWeR63UfvXh/N5qvXj+SaoSNqJWWwUxKT
PYuRYWqeVySpBU2T/zugchR/bXqk8ZyDq2XasZnvIkqmuypbnqHEvUiAuYbt+QxSWgIJxqQgC/6F
H640NudxSpQDUGQWXklph6WxVENv+tiwRD0Y9zeKhJb4Xy3rz/k+RVzh5p409OrRzy5P/Qq/djOr
SmODZVd1sg/KrooZnG/c6F/N45sR2H0S3UEUDKpMX9+VKANECcbL+fgU9XTONTmkWvHgaeKe6euZ
XTrEM9N1oRvfiQusKebIoG60icxlEyVTfsIPeRhA7Vdm+rzyuMvt8Xsb8P7borS2R707rBkHFwiD
YC04bmWXNrTQF57HG4QXdjlI9sjs7yWh/oNrxYHRNH8LPEWpX8W4lXQZOvw22KmM/wqg63KXpPku
Be8mBxMdNJya0YPmuwtwxn+AJRH5IygtyrOvKzuWtDA/lnUM5IQaoFZ6wpfw283pWkIJGknWSy8j
+JwFCo1lK3LAADpFTM0dWm+UuFiWcM3K+5QfdsKTpKcOI1+AyWbo18wIOn+fQHo3u4Pygzw2pswk
4pRdbvI5J22K2b5onOx7jPzfzFNfCcOCWnrFr83HqJ+NJz1pkR33oJx/JZk+lq0x48Q/TTqFobZJ
h59N34wrSw8K9CdJQKK6+oacjOE5Qa5zTINmVBkck/MJt7+z714C0VcK9otZSyVcLMvEajQIrAgY
PtMHqdbQ1JL09X/DU1fZ0AI/fYGSmgQOWEuBCmOlIaErBntyrQnGXVncMV97eGDuYeZsfKTN4BJ/
zoFGtYbSd0rVtJMHbo7EQIE/9PtVIDogpU+RMpfSH0PFJPLmYEdNSVUpGqmwqVKIlcgOK3DCYjyW
wYyeOc0pZN+2mdpdr5MKrjUuj5yID5+3Al37OhOS+cslsAyTuAB2/njifpK8YMvtBCCHMuxuUp7u
v7G39G2/aBP5XOy6ncUrfHik9Mg8/aI4szPJK8wt7NRtijX9AWnWdXpVTzOQPGJpsyZFucJVaT8m
aD3iWS0NRNfkFQvk3n8gwHt6ZrntXBgFBR/66Iibq96j3ck7QVCHWlxAsfwnU6mqbiqLuOz9X/AU
muz4taA6SS88a2i8zSEA2PWPTh4LYcqe6JgIzX0knBho3L6N/SlySmRcINFxYlwvxlptTpMR/HSs
X60jm9P8APL1ZsrTHqtwCJnQXE4bzLo0KhEu0+bCEoaQwuZuh5xVq/bBMV/7KtPaYqUn6d8hmhYW
VAcbRU5mc4/Gg/AW0hmmWLUhB6+td1PqNUW/eoBd1B+umeb+EWtH1oZVHFHTdlj+s0fRVpWyZD5p
NEgr3D8o8JFTkZvGfyQNPd/ymE1qOgSRn3jWMQXUPaSYltatPnzor1qI94oz1OXeeftw0zxY8yBT
4BdGZcps2atdhm00rEY1sA773MLsTgoXMGxAyf0KnNr7G34fs0c5oPLxTJu9aq17gZtO9A1Z5wVC
+v20mmoF12hEmEw3ez4OJy362rHPJC8cOwvwf3Dsp+SHrhZo9w+vIPBlq1groBlBUMQxADGgR/Dh
VreH2+PPPWZP21qAnTN6B/v/2TPGpabEKB49KBN5wVPyHgJ6byvWJzjEipL4VjwigNVg9e+9jyl6
9nNbp/lskvW4FIlAMYYyCZEC9gTLawPQh4UsXYMUIehQK2XBIS3xHWXx/o8I3LH/wYdQnbaCGOz7
o3QZy5phY3QenH2KOrO/o8cyDmNTsUVmc/CbE551dzNE3HHo8v5dC7gh3jVqsD/DEEe5DdVnO5wy
7RhlKvJM6cFbFidVebpDi9eatduv36y1MzIzsVn/2+kSyGnj0qiW8WmmiE0Hb05Hbaai2/mXETCh
DXAvz4z3fPd6YA9eprEQH9IGVZGAVmhLWL2Sjyoje16WlMLabo0DPdwI3ZC4VQnj8c1UhqteKxpY
jBV+0wATHwSvbYsQ2fsegbOVEnrlUGZSpS6dupgSc8PmWVC3/rdxxNnQ3GiPM6i/Pjxzz7oKTfOS
sPqhD7Dps6jvdoYfEMZY9v00OqTQWXU92QCbtS4wutXeUdm4KZh6qXKY/G+SEYXv5QbF4ZKD8ZCs
UL9G7VdwY/EzZtQIPRsuUnuDPgCW3Fy6Ulai6mhUWp3NMIo+YVST2gaDqTninnflbCPIh/AQChp+
BEJQDh1mJ/A3ng/Ewh/1HaZyTmYhned3L/4Utww0jdnuiMiZJWJJm9xdXq1M3wQ9IGsSWRf2102o
n1lp/eX2IsZDFGVDtxtPqCdxpYWFK7KJx6jmhVLmlG6FdYbAH/kb5pHx19fEBtSVs3n8cW+HW1kU
0L+7ptC/gczb5yK29U1zzNESSZlYdotCVH+PLo8eYoquNFCydvsRUdS6m44wipEZsUEPVzAzFfby
HlH5rRMLFIxUgqaGv4R5Y15HJUrb65SZGUd7KJSILgZlsvR2OhZw7+9ABspUtGlZO0UVMecnxx7W
ZT5h2YrUz9jkeNN0eHpb0957qe4BicDJrS0tihj1gChL5nIPOl/GZk2n19goieUxgGhkglvIfOhi
XzEKPCQm8vTGz5u722cnQgQJL4HzSn+1hdtj3630PeRapEyMr/Mqn3MQCvwWuRu2s9Iz3PL3bRH1
WJEe03H/tryTnaLLlhzIKdy/3P0iEFVq2IWDsMz54jdC6k/rXfjuZoGQO0ThIIq50ANgxhWOoVCH
55P+Vw6+SkLOA+Kb8kZykWyQpgd18nFyUy6ds8PpRzzwVK1R87/3+h1hV4RcWO0UTL91zkaOQWdi
Iswdd/llbbKNIH9lx5hja0uM3wqS2gAXevnLv222VIc9h2FRFJOVM6rZ9dw9N+bmzgNnSUMyVG9R
NcRzKmmLzufFLVvib2tJCyt/0/uShUFEIO7Qj7uzDbbg4fzVMkzomfVy8Yi7NavYFjWe6f6AusGp
tvwNKNVEtJ/ZqqjhVku13tuPJxjEW+09fa8Vj64cxMoMgYRKe2NDmLDf3NweG0i/ADwPfqufR9D+
e1DwwoTvsiXWZC69Waok1SIkXVmoLkw1yyNqEDMo8vE8P64ldGy/mSrOGde4OQ2d9mxSnW8w0enc
SVPL/tki9NPIqQml4cIoGOnUyyouxgB5WOP64rTEX/j7WP/Q5KvYkvsG8GLcytohp4MsB5ptPxdS
qEyBrD2ZdAPd4Kp0XWkGL3amaMH62rtZsnbQjg77N5RPrOCsy/J8MMRXrSVxOS5i1KVIuJRqY7oa
UGaTKDs6nQAf17HqyR9vr4B2hsJW6whPlHtt/qxUkqziW1I6ctmWOHzYywMHe3bAHw1HER777NGn
rmuhN/v+zCAvcGodnym+7HY9M8qBUCzzvYuXtAsw+uC4UDWwGUDnUp05+0SlkfaCBV631z/py1TA
109Wgj6uFOii/nG3Uy6Rvk+Gsjt/9PlD0ZHMsbNvNbZAYBFTBKATzqjWdiJtPP/LMkS33ubW3e1r
dYMA9nHN1bH2PQm6+m3RnTN9HJXTfjNe8OJBIiWbTwO2bMMuKq1O//2bGXJlhI3a/Y2VxjcBFFUs
1MpnQUVn2WKazyLllcF6y03Z3NBPWw2oUfbXpqYR0COwJFyE3hLwDQr80Ws57UfUqIorksxZKT+x
gioocmvK6acaSj3NDGqkGI6UQVkk0uJbccrLcNRbMM+FdSIF0arp4Y0Zho08M18PuKT89vtA2d1O
RWvCxdn+zNHDW9gvmSgfEIG/a0OVlCpVq1SWy9VLSz7NYUKY/5NiqnfoNGtLhP3FIwNDgN9aNW5s
y06uJ/nXmdFWv79OxOCGQFQctby/dnsAqiNUPa41HkNdmPSxMBiFtH2CpUyZ1rtZ+DHH5oEPVPdi
xK34l2GOg5Z5esHF7VqXWFlzQ4/Egxa8bCqmIS8zXlfGyWYV+dYERAU87CSkVMRNPsnvc6lgDVcE
zSOaC++v3IkP587bU/38AGX0fXN4e+rf8wVJqmJVtuNtQk/rKPuD0ta9Hl+NqnKFGN+EvMTq3ijJ
rvKH2S9AFpoVSvdXjlexaVcfK4FqYc7KIoFodxKuCdcW0bLnVdT9EWO9qB+P+ybYLdhFhuDZV2AU
WFebmWQ2i290H0+GzWxPkp85Mn0lLTkfz1L3zP9VXkvW9T7ev2PgfbQ7FBVKVPElRtfIjKqlejFB
0fFm3mPG811jj0dC9nD5phGFobn5x8SElinst5cgCEWB2Yq5Sf9tJK9Qro7KxefHtROisqaG7Hj4
9dF/GwXQl1nNLN/+2koXR6cZf8iMxy+vpELd2sBp2NsnEH+VzDQRzPeHUr2GFVH4mgfV7JYPgyHO
ZE76ErSsSSh7DUEuvWEHal1PSpk8krbBxioJeh0KXOewuwKD75aAE7Cvbdee0qR59gpPlkf0wibT
F1g/qiKh6KDji3vSDkQR7d9BVFf5HaCrGNVgmdUJ08oDB947h+l4Pdnrm5zBWpY/ACkSzOzvE+bt
zBn16hO6gSCjRtRspJzbU7KVQ2kJYAfmbkfVzd7CzO4fVF/7CNFICDvrlbc5qVFLoy1uLZKuFiDS
a7mYDyG9wfNJMoE540YKdRy1fLkMGaDSFFlM1Zvz+6RGIjaOA0Dj8PlL8QxU8DQgPzJ4a+H4Jft0
TO523ykv6Fjd/PKEudh8ieXeo3htCxAld9foPGVrDjNuDdOyLb4mDVoEh9zmN6dfkJwebgc8Wcnj
FAo+EkUYujv3rHT1/5VayqfYdwBlpio211cXu6TKvojFWLQC4xwz28RGoprAb+QA3dCIkbiEB5Kx
MD2r7pGL18OE9Fqlzk8NqXt8Qa+g4MS4IADjfEFI535yMMJ3YfMDsdnj0SLUrChAybZzDunp+G75
0Y8HYDl8/rI5Q52dY4yVyXTdGb/RN3LLPC4/pCVoRYfbZRbYMeENkUzzK/xPcUhyFYPiguMcljJ0
B/5AJHknZ5esIfj/HQjMuJ1YPt6/iaYfwOT9jHWxoYUMcugYoL9liSXSXcMnHW/q3UgUNi9X9kIU
0mY6MKayMg+9mLSRLIeCAev2EaHuQJdWCAN3rPgqLIPLAYzTnN2n10lQfLTNQdOnjr3kOVNzVyQF
TPxF5LtbwmoN5hezd6y7lzlZUhf9H4e2UG6M/Qbv27McjsYkXWcKYX1YnWymLbdO5qz5231o6UpS
5Nm8Rgz92uTItBJ+ax84dgVNnh4gsKr2Q7nApZxhrmmTBgjVFeCIog2YL351M8a4k6iWEaowvSQ4
KU/HdY0JDV6FcdKPL2K+8gmHRiNTEOO8uY/j10QU/Pi8QoD+QOXs8vPno/NxKtWsnuF56Vg2LHzz
CLD3By4aYjRppFJ1hzpwYCdzbDg0HrLGiN6G7KY0Q/o9uaXLpGX3Ku8pPuY4onDVYppv2vdTQNgh
h656t1JLFoD8ggjf0Pe8XeIFLvgO2fXKwCiFnd6ikkTHUDN0SMCshxy0jo4tW96gsq1KkfAbYbUq
lWa8E8z5XJ96SL2/q+gI34sbDj+4w+WfKy3XO1KNjgYeUFLKbQH1H6KIUvM1iV/tWrG5A1qiHqFc
CEj9CEgb8jEPiYgov7XXNYCsM/VgWmVXLd/G3KO6Un1v3ml6LCIJ51L+/DSRq5YInJl8LujTZhUx
dgQPM8nsNBpukfbQ9UMU8qBA+u+xUhvMoTDctxUlyYe28+tf6jkD+WVTwuLhiwd7KK92jStI05EF
fPMS/+v28L6P66y6qdxYSpw6+pY1Ii6V2KGvGrC3qGoBQBe8wFjAReCNnCyw1vg8neHM34Vjm5+N
e47yDLE3TQHFuHyXhGRx+7TGtybSF+8Ltehat97ga8+Hh2wXfcTHOrz0imO7z9a4sQpmpRYCTyPG
aMbjLerj5Pu/Pmmwspr+AoCemnGq6z9hKe+3a2AGWiL9ThnIhSyzEkqEq6zljkoP24gxriXYf1LL
yBg6V2BxP4zU8flksrnOkk7lpp9g56A0sUj7stsGftPANUKP36LdigSUb9ia1Sm/AGl6Bp/BVDZY
t0/Y8AxvYMcHNyiJIfqJEkw0HCkgu9K6jWyyTEkcttw6LGJyL+X9cP43IKzNGoWhC33+5mx+aG+c
l6flGuZ90t2Sk9ogUjC7qb5E/iqe16V6K0sDuzTJaRpBxvRQGNUnbSntBzhJUzfLf41+7fvGhJh3
1y/oaXL/+pT/wEv5YhJRKcgVd/W27/08hamQGolxmdT5f+Z9D5jMlm6IexZUJXjb92zk3aFHjfoy
C32ywuJgGwjD5MtxO26Do4vPzHoMCbtHkqU7yWJr1B2uB3dFu7Au4vGc9tVSXQlOPf7sbI/zKyZe
iC05ncgVd2IlUQfS5IsTX1l5PO5d4IWTRiiNKe3EBng1QW6ccSEQEzX2+W8IuLLltW0jjbBpDzrW
rPqOry24/r4qdKOtjPYCasfcPvhCuArDDyBZvwBKdBVbu/ORfZ4Q003gcx6xkXAacaohgufutIQK
dsGqX+KsG/2SAr4CzLU0FurIyoxAOvN9CpHTLT6ZaSFUHTBgD4XLEMARrtt+ApmwF5pL3CFrHo5A
yL1h2FYcQWDcn5mu5XNP/BQ4LHxxX+w48TYfZpY3u6Eu7faYRsTmaEU9uwZhFBcP73ynLdIpTwyq
Mz3AdZ2JuVIaqaWNoPj43putdFTgOz2KXwK/B1T+GCx+N4wJxglBnb9m1uh3LCh0ceVkgbnCVCLW
x4OSlPumT+25ekVy2C+0GvMo532aADzrTEkdm5zGAnwUSS8FJPTwrjqQ60abds4R6JrKOWOiecTt
outpe7SlrtoihEMrGT+Bb43lyxULxr4wGqbi+/hB1taDd/ma4Gop/h2j2+irW95OU4ftf0whCKYE
sf/SyRn4++MXs591YQOo0vtUcswkRAF28pkxj2OQjE4gLzJ9EL0wvImjRjXpO+NTL/xA35BhsQeo
XnEJjIiFYR09wwuXRUlL8WwoXF7NBl87RowZMZs/26dNOhp8/fqdNjQ2aL0WQrT6HiFL21cEbNxf
CSCSOWeNIY+cJzVb7hRiuG9Pfzbp6OB/fv+gzEuuJuTO96piSlPt73jjmzYIziawwf3+wIa/toEh
Shty6Eb2g+eN8ptUns14DFZQO9BUjWJT/ks8YQxn+bOvmG2JgWlhw/4+lYFsG4Rea0yfth3qa80q
jdxMdKXvvid63IlUXMgiOlaP5CK6kIPccy15q+FRt6TugadTONSSF2AdtJsKHNfai8W29Z0uKEZD
pFoZFZG70qxdQ9vWjISIYPaEo3tW6EftEVmgANvz2klWAEQqRNdStY8zSZUp5bGT9/aVlJ1iBmYi
AcDx8h5RyGSA83DbVpAV5aGMtAVyUonazwndL1JFCDJUo6ZlM7Ng11QHBoF+7JyIhLhWaSxo9apm
59blcNWXcvCKXQHP/G0gH2lkrUwAT7XKekiSqATGhGUGFUXRWqQofhQurgQfzVxLCBhoZpqQ1Xk6
2Pm94izQRCshtWr8B6gckdE/3k+UGDsct3n2tZEurHAThFD7s6ulvBPoUgMP52VX0o1Fgw+GJ1dB
KqO9S/d9AnZHnf0N+HlR+CViMCXA8jafXX6WEDs1CwIm2EE8Hk/KeGRzZPaNVOZYCy7UnCEhBrvI
U3mtvpflAb5mHJ4zbgqQ+tg3mp5gKmZrGD7ZZPDVpBzkiJriVcLcYL24IY1INpHSN1JBNqbq69iB
hhj9cm19iP/Kr5Ey78bPpB9If2mdGk7FkAm/ul+MFmHLL6nkmgBFcLojvypb0ttTqv7VL4deLuWL
L6ocy1tKOQMaRWhhi1R/IDZwYZ/Br6oe069LwtQxJ9oEDGStCH8/L1WVfN1rD+3g/TabCG7aTZwl
H1/CHQ6yQ8l8TDB3xbSqaakFcdzHUtAiaQQ2mDcdVzSs4ZJLRCog+FC2K+CIT2z6zQ9kzUPa2OZ9
85ZuqWOD69uCi62n8Chgpy8fG5R4oIQQ/4EyiWlpZkErV18g1IVCQLHt16YRN9cXXb2EFl8tzjPe
ABriBuU5XpGa5ZUbuCBI4jAGxVBSwtv1TzoLlNbRPBYCfRxVWTWNIgjfN+29bpM7j06DD3emB9X2
qBeTUzlj3GrLf1K4uVSlUJHmx0/pU+SqfpUmJb5+ka6F6zuy9q4Z0FqIhP0irxEFM+zpKXLup//C
2tOXSOnoLRWIf6HCAalWSO1LepbvFOCW6Tt9vgyEuC0o6KtUDkk0n4/eyv6+MWCl8xoHgA3Whz81
F3cNqPFZZn4Xjob6T+PBdMq/vroU4oB4cd+z1tQyqn3xXVU01os5tei+EEbkl94u6F2cEgGxveEd
M9MdZV3a0g/UuBH5crn8Q777mU5xJBof0CIdVCh+MTgWO8ibDINM8gmm/3hBa8MNTF8+kTm5l4RH
fECjoz9jO+OlMs9bqeEEnrBUTuP0qdVfB7uQQxowb8W+1INwcjlRPEFcGRb8AqegyhZmqPfj7O3m
k/pTHzHP0V+FEJG3z9djjao0eVfxEBrS9oUhrySwi2I1gzQEsQEJBGMttQ7DIHdKlgBHugvq8UB0
eJ2hCuJE8krtXMujs71Eem1CjoEtrekFz8UWQMHVZqOY21Q6J4MpihsGgGwtuae+fZcW2dOIjeRz
Q2sI/etk5Y375vaabrXg3Q80aiqwfxhFPVYLkbfNy7sf2BKFSg8K2oXsIBv9qK6EGDRgBM2OrYF6
O1kv2z6+Jr0/S9c+Mh9X/4MPOEjE1w4XVWkbd8HPoYNIbkSR5Gby0okyYScrtv8X/VgwCX4iwVnu
/TPSvbcXNp7cbAvSDw+RR/HxdL3znFNvC04Af9UiZp7cmGEY/2Daelwe8VCyJwQvFSfXCogkAiOd
SXrokOB9dYZJC+E5r0mgh1dH/ENqlC8q2VAjcETPjxkaihszQoNdIU8oM/zh4JPuM1uy+DzW3WrK
n9XuUtvX+ZrstyNpdN6+jxcNTx5mmoirFpEtEbTERDxKh2Qi7fFxnXF8qss98IpUklzRb2n9TqHy
e4w8LQ61euvOG9hX5T3FYHqRonV1dDwq5yZ1TABnWslOS4MPhzCrgZ3MRGq9khFls3570Dx1NvWr
PNBQb9gzDgH4jZH7aO4QLzDBf2lz8f5XoVC4gLdsDCsJnmAN1js7PxoqHrVG0GYjoIjpCy7PAqgI
fNQ95QeblKrxuhKTZutvIDSMJS3HCdefq4Oc724RerkVJXPFCrnlFdBiQSnQ/YwYOamt+30xHJjk
xjxD9cd+l0T/cG490y/UW7EtxMZSqcK2XZzTUaWBgvIG3XGK7QJZOAtRzAeCD/EDRWyxj8NSeAL+
+9zF3XzExZ0J+mlvj6Emi/lIIN+xdjP5Hs2XLfBMAhLH5XvedMvZ34ng6XxahysbTScbn/6XCGxj
e5pzLU5T5J2K6F4gUfMOotL35WGauUNiZ/CcR6izfM23J4+WGlVCGgd7WcBQI6LLcll8tP7z2vXq
YnBoekIwHSLOLB7BzW69QR1AVjAJOj6wlvwB/SAJnJkBd6/LEyMbU/IhyMEfbTzMCnaf1wizkG8G
MlPViY0xqFhIyIuYUS/Xwno2IEkCKhJuajHo5Dn2/sX0HbMVUAmcD10wos9QRMPM/3/tTycKCocn
zPDDUurWojvvPkh3KgfFE/60rsPuQPUOaVhYz8IYtiHuoYnNEdm/x1a/11JiRHOqsWhdymARsme4
n08MHMCukJhvzBvnEeUs2OJW6EJzZiWFMbjZa7C8NUo+MpIL86wqaZRSFPLMyoOL1spagNeXWSu8
81OwLAcb7i1ccWhDjXJ0FpAqNHexmLxVBj68Ff+oHirZYCAVcqfgetcCZwuDt/UBCMwT8aCpjtW+
6yAaX7SdSN3LupcvUYGwUx75AJrubCUtZoFCMFhH2KW9dOfQL6q7XUIZDhoRC+BB+uecTHZntunR
bz7sazeUZsTJbE3aaD98UWAm4be8HhXMia5zhTHWzYP7GpPomGnVsBUawL4OupG17AIVZ7XJpeKt
snbd7q/csPF31irRYQBw2GROesaSxyRBLDcQLOFnSTX1L0veOMqZ1TG/BaojtiCHQBwg4Mod8mps
dN3PDFMtn06p/Ga5ln5CkwBsvgiPUC/5E7lz+/L61nqKw1YEMwi4hwgFK2a28Mn6CiDy6WlnhJAd
khTESQmE5NAFurApu7ZJCwrRNJMMDRKaeONNH84dFM0LDwMb2iKCd0p6jFiFPrBZ9d3gPCkTtS0G
K0FUQsrFJ08BLLTwsfhvai3QiIxYwP0PPfpsa51VB6fBaRZyqEnaF3/xfZIxcLoCLBfChKNVFx3C
UA4mLlCVfmP8qjQ+D50fDXU+/TadxlrlgXRBefP1TadBy8fdj9f2yA3D5t+/xJJfq2Tklg78tSFC
Sax/zL22lNXDz2HJvUEXp9QbwZpElAzYs/9yPkq+qUwuxJAZo8JKhWAnkZdAlL88EiON9YsBaUKV
GtQXy2VEo4ZGYL7+fDvruwtWtvCSwvvLOR6LnAFPraxyufoEwbyHQiRu5QDaPwwBYOWSl0BxBI7j
hAFRVTcCycshLwZOljZDs0AA2789kfRsNomiLtfjE532hj6Bc9dIbxLcKpKEmtJzQN18Cu3FRYVQ
mgGCy/C/OSrIw8NDhMm5jUVVUZVtgOM1xvqBaJ4ecQeR6TAspSiBgqBqswkXVPy1yLCil2KpXgkQ
A6POvdAzIBf3w1Sx54R5wLT99QirAbyY5OJIfuVIVqPOOZEmR7GBHAlF7eR4uFpnP17oO+aw/71+
At1W1IU1vxtJVJIZQXmsBJzxF6M0uK5/1dE/ZRr9AtcVh5O58bWTcskAWYGz8JDPKSw3qfjw6TH5
e731N/K0nrfpCxHii03mUyPSCMDher3j3j+8yqdWUqrqTzlZAiJof01tblSvRF3NbmWZwUijHMrD
avwEde4NnIGUmt7xeyjMC64soo80NL8gItng/woMYvVdStpH9LIaBGfrufLKfUjDwvYegEld0Ow6
2M2PIewSERiiQx5KOUUvpPvX91eUY7+fS5E6/RVlu2wXePujDSjRUvmyKQN1lnaRkLc4A5TW7JCg
p1NdvZRuAg2/AIIl74hg5m4vlvwVhxvKuO5J4p6qMDd9WgLieXbRwFFdKGM1jw92EkspqmIW6Ebv
28Jo/so1omdzkrbU5Mc2VbHxyG/gb5aVXMfQeE0NKviK33uB5R4q0mJhRCalCW3vO863bUty3wNC
0b2jjAPctbaDDRyq9IlsbZ+gC7WpUwep3Ik/4UR2frTulasDTMLqVHa5oj1VPk4nqw8KClCzQ4t7
hUFSn9XYIOn2cR1YUvyhDdW+tPPSO7DXgKQ2N5N3EVieI10yjdCGxD4BCZSxeP06ghROhFhxULKJ
m5iNFW/ukgG8udTggaloSPYpxSIOCmbSxaDuG2pAZBvDgwxdi23S441qAeEn/bRzQml8oJVy0gRH
wRSLT/FlXqSrVhBuR+z7GTP+GQs1rYFb0gbICX5n6u+ztZzRcf/gFAlY74VSdoq7JRn9Z+4SftvK
8S4RsulWxEocQKEFQQrE/ZbZOQJ1V5ximuGsfYbmAuAqRfjbsR20YoMFWzUmOnPUOUp+X12whk27
XVo/dscnUohr8/lBzmg7yYlpNHw5nZl4zxCLWNPM6GPyI9rYSbsIJYkeA3AVmGaQbSYEKkNqe3Ml
wVR/zvjMeaPM8LUo7yD6Vm5o2EkfuWdT8nlvUukP9+94/83vdb7GSjkrVZeOPI9+RpVB6E6qGBCq
YIVIHDfMXkJ+cR1+q7xVKhToajcpzWkujyxRqBz0Aj46VkApOGkNdu8w51p8dbxf3dHHVLv8c3ZH
lFlrUaXRKyu0TrXj/5PtuQDGFFzaZfwc40Wq4DvH6rOgoo38jq2hPPViC06bw7wTnt0kTxPW3V3P
R7xKxu3tdu5AxWyqJP0H/GbvG4hCMHOSv12y2RULFaupDpSwBOClFa5kXa/zk1JMrJqk9mR0LS/4
mk3pEVjLUiyDw3euoVKyDVL56+XFYlHiZCfHDbp3/ea4Ad4qH93ub54/GTB67RbgcGon7mNQVU9O
9HSZ3PFCeZ7jOqcVl48Q0OOAWIkyJIhuwoSKHsbtS+DJOMUusLzPsR+8Tht6pB2/K2f1bbNJruqF
O8tYoM5Q1vOOphZ42fW2/wUTsnBdcsoeAaHCicmD9pDoNM+jqCsl2YGUYuhdtpz06Hvhe2JM8lGG
42kcJzauyy9JQ7EKeUxnNOU7vEB1g9LAfuNF+hBtU5spGEQRbAhsVqgVLkNjTIkZNHa71q0CipCG
u0hth1zQm21yA1IWl/SmVr4+DYgovQFJIJzSboMnr+bh2KemHBv9Ab1bES8YkVUi/ivoElYoeNPI
KYXS6Yy5CIwArlt9XCLh2YH6WxhLtXencCucQobJtSbVNZkXbPASeaUWOdR7wYOHIzuDCTRWIDhq
jXWuIbZDuTiMGOSyEZwNy+U4RWwU+4H/LXeiIm2OT1f9mBiaMsdR7RiqylY9taawK8HLg4ZJQJsP
v9Lq5+DF1HBztsA0RaHoV/mvWciG9WGBXs/cBGHOm47ksYJuSdo2SJ4hCt41B9Cpm1Lctu43B8D1
FoO/psR4fLmnDsV8Rq7ruAXk4V3VSkLTrMA0MaOZ1yA3t//l+Ftl4d0ZuSUk6ycQSGqzKwmRyqUH
I6C86s5h79RRL28o1RB3uXX9v3OdDa+XalHV5KpQWPdmo1rxmGjOGckqYKUhcs7hCyG/NWYX6fXo
AgNSQN6cUB6jXiK3ERAkVln/O+hfMSfpoA1STpPqvc7xdEoiWy5uSmFXytmCD9ecPABfRhHZTJsf
YX2LqpBJ/q49iGGBugZjPkeCLPNFP0mSy49YkIhRSnCskbf/KEViSEO0u8qGJjAvsxDJWOfNh3jT
d4q0lXX1V3N5AvmWxXkMWB6NeqExusGeIQiMghs2vZreNfbxOtQTmBH1MZV6qoZ9HbdkZzBo/K6X
2uSZHgokO3LR2AVy4C44dhU94zC3pzeYlETc4C/Fs8bw9EQ2hhdqKuAZScnCDOxh8Eqouo99AF38
DXUg/D+Cq53EMweE/3eh+rufdwg+m68dfVLG0VaelYQFJIOKBsCUT+oto/2w+/l9oSwkxltFDQCq
oVwb8k20cMWgeQyVAqOG/YVw3pZm6ZkIuQKu3e1BzRa+4N76Z18+s+936kpku/WjgbmwKu+gGsy7
uBanen/5LuzX2gGro4POkCL+owtKk0X2y0gH6II1c1liWqal5IqRsu4qvdyDJifKYtdvb8SaP+YY
VFGEzJBJB/skTNQyDJ5gc35NcNsajoU6wk4QATY53fdGbmxYiNlkK4U44YVMfYuhprbHzwHXsOD6
si58XWfXEvaeffOxmQoNSF+kSSW99PCe6vAfBKmPlBGBVqCRO1CftyjljFym3dT05buE0xWP9ZDv
guzia3Q0/xYiixdVfBLP6jkMF9OjuuadT1m0vKI05E6iP+32V9R+B5zb9pWeOEzhHbemLYAt/199
4uSmkUVSqM0BgMmGVUr+hxXlxBVZ2QTz9QTYN1sPACjOgZylpXaAUf2WQCrDMMdd1NiVHmq8Nkis
2CT35ekr3IWvGQvcChQgaxKKgv6DLRMf6J80TKwI4ZvQs9dxD7mLw/kpFNAAGk/NBz9IxnrJprFa
BxUXYh62qJU2OBS4RFFdfF4USgFiDHLzkm8HMFYIuvuLP6xIaEfAmKr+VLy+8mqK6ExvXWk8w5OU
/7y9e7GKFgiEyI9GNm8nOyGt08RXRkrt55dxX8V8SWjL6EoSGr32XuK7Ar2BdWt8N/TJR9Lm1Z5k
wHSTx1rFMkYEruZTxtERPZddbpFFfiog1DfqC4uZvUSYwKhZNYOh8kETUUDPptmNXk08vDNAKn9s
s6Zq4qUAuPemg/UxtPcvSz8hT7Ss69szN25/OUrri5qTMbXblkVKtSvMRa17g/vjzRxhOyXykE/d
IltMMWmTfVSp6tKcBVU1gtcToZaWTyqO6g5RXJ9YexzW6hd2I8DfNuSPAAeZt0Rydrrx5iIfGPQS
KZEGAfwJ2gwoWosbTZXyjIruPxHMXIDoTDM1yDcBF2sqITpnp4S668tgk3eEVmjd5VgO36iZ6avQ
VZrr7ET04O5mhzUN4EzKlDG7IBqIATFsGMlteNxR5Yu28ruYRThgQsHV1WdIzBImyQDTlGZs7C+U
kOrbBdIuhgpMnvlPZA7qhk92YtUbhQGe3w4kOBXAEUPgxB4OCdXRnXoCMFUPWtcQO9fsoGTf4LZL
l3ZLp7WdEKYg9KK/4iVB4on9mMzwCtarTJMztTYzE5QRxYcr06fXAanQjamO4mcfDRa81IyTRQN+
Y7AZ1/eO39/tA9OCAqEtT5uhc8pOjk5H3YHPbzfD2lyaCu4oROykK+eKQwxDBZFqNyVeo8TFUKZo
rJEbamTEgjwMy8qV03VXUjSrufPUgEIJ/HJnWgCAHTKfE6BSsfncmqDJ9Sh8bKej+6dx45we8yTg
oP6LEfFaD+6qIh2KWFR7xtgbFtO8MJfncii6LJqUPov1VQY/xcNuecQPtoYXvHHrs1dIAFZGt5r9
l0yOu9kKiN5i0mbWtPZATNGgEBo6GyNffQe026E3Q8+uVQfRr/YweWJB899/GZqf7B1LbcDvkTp+
aXrhzDy6d2Nwt3f+zYOuKlkoAGj0D7WkUS3z8KsI0b3ZT+OjvPlwDsj//md04c+0y6v7DQtWtIsO
rgDll8hEhbBniD5QGyx9LMGJ3c3kPnd1CKmDQMVWawtkBU97GSqfMKDv3UBsZZVAO4ieQJb5R93b
2KmCRT4Dj3jolw0fVvHU34YxPJGWaNE4kxQtuZNrNSbhKtXAEwOh8HlAPm5CG0qEACU1JdRLvF+0
PC9+0LamL8UXYTba1n3c7li+Xo29xWhojaju7GgGES4Vk5pQzpOkvmXqqfkbVzkFKkjum0nlwCxi
sZbcLXKEDzZ4sVsFzQMpy6MCu/7jtmwwWgVQv1gSo6fQyveeG7HAuf5VaXH+ShYuQBcVlZHV66WY
QU0vtbMToc4YuXVSTFBG7hnWOX4OgrfnkZ5O/Zn4qYGKuM06HHgLPkY5bK8Sb75wc/VuONHb0uP4
DmWmRpG9MtSnjLPVTrDtTebeYwHpXyVDURZwVxiW9iNbG2hAanZWduGSJVodfo6B++lx1cPnT341
7C30wrME2oMf4RmF20s4NA6esdInsHM+gOXx63JrsRWidyhrgSnPKjV9XnWB+nJCOP03amlzCyVo
CtAmzrpdoeVAKUfI0dSKMusxaFRtE8u7PlJqKeorKK70QUvHj5By9ojTHHnEHtblFzFpcOEJpCU2
9BZERRTXnKO2eDFUbmrrBCCvacJrAQjJo07azsm77otokJBCzINdTDgJaYeTfLRuFC1C/20bD7ky
fJueyWDDXNLpjj54EWvJlJXjH1WNSOPDHanzNMjrUIaRgGRCLOf7FCccTmeqLujdmOvux2ZlHBXB
jPdEo9NXCLvQdggoYFOuUNRrhy2Cprn0f2kOmPOYYNTrjoDPVENZig4TTr6v/AKIsMQD1hcPfE1J
7Ww7shoESzRsPw9Wok/Wpz0erS4LY51NWtmMhO7JPWlpCxohxx2dhXp2Fc57hjxqZwUom4tc89qW
pW4Zq4gRpgYWNBZ2J6Sk+03SRH8G7OXScgtriJ0HwxqsWrOZ9za+D8/plAAFFqdxNk0A911ec3pC
4kntpBBWUiZcUOW85QC1KeT7DuuPC2u6ssJtR3wu0ou8NXMZQLGuGYOs1iXsCN3Pn5CDcsdQPWRX
vYWbNPo5xFuF44nMO4yUt4tgAzvm5zQ4YLlkJsmnjiw0msVOyZ4rZgVU3dAT+7pJEIWDbtQRDgYz
bS6+qbdRG9zigwPJxQVL3df/7xsDUyAQKdyEo0+MGLOcCb/AcY4PYSimR3HsgsFd46892AB+DA8m
e3ek9KukUXtZcATx7fTHTW0d+9597z4CPrTjr7oO7i3MnbfckWIYoDW5QG8t27saCyJVHh2vnIMe
ontlvYLThq2JcE1v+xDXRF6Y9wrAEkuHCFSDDWPbQ91ffT7PONrBmDD2fwixA1EFhj05iASg1yJt
ADOtRTRoMYOD6S8pqv7lN36KKBag2oUinFRW2h6ZQgu+tbT/goaz1OJdAGgPcxZP3P3mcaU6VAIv
jomO288QTf+qaUU6LNuORBv3GjFMB/LcvgJgdlaV/myLyaI4H6OkHFpwTSASk2pjB+m4iDw2MKMq
WiHjLcOBZHMaYFSta9MIrUBxWxap//7TDg/lk34mk/Ye4alCckXs7xfODVnW4XPwzzmowINTb93p
aHwNjkf6tEoBwYg3zK6dwYZi8B3m2SmMMHzH3A+vGh4BIQyQx0fsti5zHCPIgVRhrUexFQkUF67u
i5TND0VKsfx1OwGoK16KwyNWMznhTT+xIe33HSoNzy9tuWWZU30hhOPSndh74Dj1PkJmfqjknL/g
DVncGZ2rmqGQ/HIuZBguYWHsoJYFFs37r4O8SBdKoj8wKU57ciqKaGVtX9Sxa708qaikHTtWurFV
IxNKpQUwF89bjrJHtG6FP2/WkbFe3gbGfCe4Xo6gHXwqgx5eQNjgfky1qbKweFo0ppHf+EwC16aM
Vu0PRsMNhx8nyR9qGgn87w3TOxywJZexyh/hxcoE+M52l46FIVCM86dQ47BVX8ugA6Av6QzlzlX1
D9FimiWw3Ts8l5nr0OunrRvGlWrpcueoabHLasysZbVAblpHMNe/SxSWmSnzSLPrgHFNTkbg2Gb9
eKiwC960Yc0OTq3sIb+42YOqChpncX+OOaUV0ycQWjZ1buyhDO44Arh/M3bR0rFqyRm2Ixi1BrBY
w8ART7qJY5GF1ZGMzxURv56OKnagLc3hefM+3CDZB+u3kJl2mv6yzVy+40vOEgU8EJu0nVAQuuf4
KRwyueHDuFFqzbdVE7vNuk4sKNw9B2XCHV2aywtwet8Zre1LiCw8quovHlLw0i4CDNgij5IZ8NoW
PJVYSJRvgeF1pv178VXGDjbS4mhA4stjFK5SwVKqW8yK9gfhvZSUg/bSjV+1yJMH7PQM7WDhseR4
AWogDLS8k+GEqBmzHpYQd7BcErTDGBShAGV1x+17+94uMQ0eBQaEb9M88kHV4l+H0kcaED6ubaKi
7Vrw6f9iJM10QdpmP//pMfCXAggOKvrqIuSlc+L4G2IKO1puQ6HlIV5HSCk9+7um4qhRBoaLAX/S
UOBHoRiUEe71hXfy37ZJ8HtDQIJZ8nhX09VViAt3ngYErQP6njmMT09jmzs7t99g6KL3cxzXijnq
cNrwhc9jS3NWftZIXOogM3Qeslsv7h+tZLOEqn7PfqmVxuQnZUxMx6rv/6I3np+JNCX/kVwuhn5b
sZHFhbqbYaHEHeh0bW7EJCg/LHD1c8tA7JcKPZL9o/1aa4x9/IEnlRHzhejiX1HR4z6Z3toUy2zD
dZjrNOofyAYABupRdzj7Pmj7AnqQBgZEyq9x+rF5c5Q3UIXeyUkEn3rIphHtsuOSUZLlM4kDVsEy
lUFBmufSvo2VXyNATzMLpvANzDRVgC+INrJe045BpcSHGUKQwEg+kQJPVTZvasMxKXpQAyLe9rAB
Beo6++Xc0HuHr0T7Gok8eC9HvQRzCsQJjJAGDX6ULPfAc0IYgdzjx5dxpT98mWE+LoJWmPB2etoM
/TMrzfwBRBtRd6nYb/xSY0MiUwlfQf4HcYJr4NdqbBD2BYlCG2LlZ1p+LaTZrIWqtDvrfhrlBUbD
O1bZmQMAqPb+fDNSGSKbJpetd0HwZqKBs1il8bEXDGybD83gWRRFQ4jFVqQ0wQxQAM6GkIKfoCD4
O7D2nX+VDa1wzvG8IjnAGKcrANrkbTQosfR7TYdvZWKZ4JzvW/xllM9e/hmsX8yzVt7ziR9FnyA3
sqwjCCrA1Tk4caBe3hCjBxDoDfGf4EuCUxSq9hZBnL02+OZZM4wK+gz8I/38aStjd2cJAfyEzo2V
2irBoFmVuUWKuGZ0L81J2wwAj77it4dm4wQsswfEWDL1C+Ub33wVhAy78meCFvpyxNBL8yR+Ge2k
7qyJELbYEu67t2ipk4/F9f3VreaECws8Gy7p4v+pJp1v5tjKzKMiaOHUabpW2BZk/BwVEmuz7Csu
q9qGv7WFPM5fCLx3R9J1bYR67N+XkvDaCV7+y/bMQOrVmUTji5kgMr2IIVcQL40jtWRMCgLXyWGg
U8qXBezBBkXiKY1csoOLEPc7Zrj6iosytdxx9D2VI70tMNxvlY/OJDSEu+ivvRIReWXuKcI0Irf8
EMyVLqQZ2MaZLr+91DvhzYj9+KZEFFF1DExjxxu3K9mG/9kWAdK+h7XYl6Yj6WkiEZaTr9NbojJ+
7S2qIRsQ3/GwMK+O9ca0ylKjKSsZdgEskg52skESbqlEac3/eSD7SYaKnMK33pnpAIFAyObvVPDT
7gcMKqVITVXTHvOe5g2hQR/Maolg3fGwIXzpsMl+1/oW6G4tSLZLeOC0hma8mG8WjJEYnZfsB26o
VbuvGQqXZYY+QvkCIFFrqYPESL29dxGKbskv018/q2XxNmOj8AUoc9UTn5hVQ3VmG+8kR0rRAXg+
RR9pdr7CFtVmgtyxBNyiX/3YPftOrXopoTvN3vaO6y9BWSZHRyqXcWCzjlENUoLMq+mKBkFEm2GU
7V+xcJ3O2Og/N65xRkNiceD8BUBavufyyrOtKS9/4ioc8/PE/k7aRBulCvdmwjdFrN4pefu64VXE
XHk6AER8/R1npDQsEMAxPnIc2kPHqgiuATN23lSpeWjL2V/5xASRIuOyjcEiBYX3u4B8tm7elN0k
Cxv8Siefb8jIPMIEKMJZQg6bOejif3IWOUEtbgvBPeNy6C1nPlFxCRB/0lZVSyCSDHOMZSIywWeE
QQcRjmF8INaU3ubAL8w0QnlxLt5EEvKzTVy4NmtJKSBKB98i9qXBvyBKhdNjdW/ZEKxvyfe3GIc3
1eMPMY6cHxtkyradhBKoX84ZzfeUxZuHouRqMTiI2vcvwQ2OggTxYVgInoxko+JXRWL4FBMEtv+q
RxdEa+MxIvMIXJcNLy50qpnhX66gMoEuWE1QcwFntfEuB61OEE2OXF6MU+QAkj47/ivAQwZzS6Tg
j8QeGzpunGUSDPEGrAVO2P+qQJYJa2CfTF33xRPEdJsFfOVP//Wn+NcoOalmlr5/xIFs9wjRLsVN
Dw0NuZvkgENg0JO5TkRg5Aim8a4IcRqhj5AHphEPIH/IFIV07XXwo/aLYCVFX1g71E+YsjD8SJOO
C/zEttD39IqK8SzY6l45hMLS4FXczun4pVAaVQwvEQgr7lWFwuoD0svFMH7TYnAxG09S0mvDLIWz
DsSsa6BWAskEeGNM8p+1lvzfgHSXgXVfoQhpPEMhjV6QuS7Z3EFhKnuYEhk60C9kIGJ7a7c7a035
H5wYLm/tcKIyunEZg+SFK+Qm94fL27rqXB7uHtoYZJ9b3gnFgu/tQB91Sn8Oqkw3MmepUsVqR2zJ
G4h5zYfv/+B3///MQ3C0mRtqyBECV43YTFMWP3vufVahbU0mxCaDhS+lX+3he6XnhQGY1xhJZhNi
Ldwq7nxCxFmWOahrMQYqZrfwZgKYhLWj0JbYHLdqmxFqMfUl/1mkceJtUj58Iw5SUSLyCB2IhtOb
GG4JI5oBViTJcgib5K5tzKulD6rV4ZxRKVvWFjN9OR3lLkCrsH2Q+FOI7byDE/q+lsl0TzIk/axs
+cOba8XcoQz8CsUimqaZK1eND+h/Ps4cqQU3r5HW+srL5klNcsqM72QCeG4R1n24J+SI2kzssSNf
Gb6VAzAwiCp883ODGAoIJ6l/QamVq9oqJgJAvHge4TWU/fMyWucW8Q1Ih1dnRwmw9F7WcbrW7aDM
29sRTsItnjHkKldBfxJJKVbrbzum9Uh3DXRnuXAs9xZT2mfI66GIHsGWMECnSEzpzHgNgcN5ND8n
XOPmEg6NpU+dwxJG8SFkpOE2Vlp0p9bXCmvnYi2g4lkppPwtMsErMu1mVDgcVZqx8U/iylvXXFeQ
lmDUCDnGfJghTl5PZ63pTs2yMhFNyqQoqSoubPLkPMdpkLlmelQkMDgMTAhGRoPzJu030HGhY9Lk
3tEa+6d+a/TTUdU+dvKGNxe+diJPg3iW/LDHBPsm3x8todJ/HTPdZlXViNGkX9t/xw2s9kjMnlll
GlakG3NKJNNXQBnaRjukaPMpZ8ha90GUWLPaoz+eMIRa0s89s0phoDOQ0FBag0KPthJSY9yveLMf
T6uaKv2qtxdlVnlgUnIIMzsJquOJSnaZIDClGsKA70j6Z9xiAUw2Wb3r+mJEVUFEnc6dQhmYzeoa
c5P9zgu5oaeujPxb5WGXd4ZLYQHJPXK+bOfZPry9P3geIPlt+KUTCIeX8vXfgz26Hjtu1Y6vvqXa
hs4Ykp0/7rPeZTlyaxQ/bmA9ZAaQ5l840jAYawNhICfU429u9fyzRkLQpxH00UCyhOxF5wSAWVsA
uSFEkz4EXAyyeM2uPKPFFAi+xT1F2AV3btFTlnlRhtfp4T6Aqv8HNrht7WSS1rWeaDayBB6sdBsi
evzf48kFBkffuP/kaXDHjL5U8QaJDWN2Gd16csYRdv9takeFqs4a2NBAjbOKlv8FnnR9rPUXRZ6L
ygisc6oxnVnBkcihYxL6WAck2XQGKPO7fGwMgeazYjOLBxWXClMXQzZq+uUBm+6w6VcG1Q1lOiQQ
Mdje4mrVLORc/+jTbQTi32OixWN0KG+8WqI/Gkgl+4CjvHVTUyzp8z/aqCJzGTT2YAc0KUbik7QT
87dS4UIoV/ywIMeB5hKUZGP6HicVzxZ+iH0ivl7EpYL2Tn3ctya/C0kDSbKHzV/4hYE3Pmr8pFr0
CbziudT1kThDjHh2NxDu/t+Ufvj98bzwsD2t4OZxhDpqSYDSXNo5Zj2PgJjoxBBG7UwPZGYq6+FV
sng/bNBMj5yUCY2aJlKnSm4xlrXkGHW/C8Uj9cctTLZboWgcQNjcNLyU/1QRVM71gMCnLoPhXHYJ
AtOk9mt59f1kuc2XjGN+FP72q7PeizYKAcuUBOxHNbH0rTdGtaeyJjrN6mIuhL6bc2iiJGQANncd
8VTplq72ZvUOjzF/N+jbuDws5WaFJMVtUA6K7/uc38aO6OGfFvCEe9+LMthO9zfbAD64UN0toxh6
1QqWTt/DKyPx3ZrvowUeKQnj8hDL74yCvx0U+PTfk6L3gPkfBhtyhfsCeuZDIEP0f/yPgXgVhvo1
+ZRtbhUFzfuXWQNwGTe3EwZddIrnfUlgZrp0VtXeCTiA9bf2JSeO8L+tfSEDjIpzobaWO8dtzNCX
x+y81Vujqutd5fm2OMPsThlbvQnAzzMazkWsgQ3Kf0qfuIGnBMy79SI06gYg+hgg8Zzg3iM1fdXb
TAenW+EupX75cQMn+Xo0L8kmpBzuleoEY7c4edLbO/176bkqdhpA8zxxSb8fw/z3O2nnuPIFAuEy
xa0H5kez+8ZPk4T0lkqOhQWmIjdbFZUHJgL5e+hDTAPHgLlxd38zBzDedaeqSyb8Hus8IDUZbR7H
euFLspdG+D6qCxtMFmWoVnkStR/dyV5GpVaEd2BVRRjDIGMPfRtBl5I8iZpva2+pADhyuZF4xunj
x62Pe448uUqCpShrFhwOm7In5N+vh+agSFk9s7ME7ZN0YJnhqrcPxysOzNwzxKzJNih6o0sQEei/
IyBdn/tnAnvNrhDbAyS4HzRucdO2jlE7h9JFJKpZjpqhGMBnMK0f4Iwjxf4dYKnlF2VrFmhLbFAo
nnRTUnm5DeaBJbiPkdlFGoYCJ1Ia99lAJfKb4xVy4CcW5V2a+yt6igoEDrgL1mi0A/CNHMZp+MIM
FhQdxOJtO8iqSuXz4rs6a9XVIuBCDLozIgSBdOQBkkH9bJMZ8sWFYTcuMXIA2Tg0XRss9D4jgkNV
cAUbEmQj+A1E6138/2lme4FkbmLqLQnBGqX/4rsR8L8JQ3vINoCnE/VGl0T2usZwpeKHnHAGL95T
8/SZafu+MG8rCY096MjQwtUtAuv27Bcnl8C1C3u1gn/3L4VZ3YlpGXBNCuWOjCnHDSh4OVW/s/m6
oGwagpY8ogEVy3/0Tffzq2B/QZMWf5nkvuoi7660Ul19iheVR75+RwcT4ln/4gSmHdjc928RsJ0h
MnbwQ/7akNwHXLv2faxw0ZAzh80AarDNa+4naMKzrt0/39/XDQ3DfgnMxtt6UljVsmkMMIruAT/W
KQmDrrc43iZOEXwlP/CAu7kWm8M0en7JgrQft91L7iFzAQlfQISLWJVYXHia02Nh7+FmSfTSYt9D
X/riS7i4PG8m0md3ZS6u1QIFzebf4s/bpXoLN240hjrN/Q5ss+yALjtcKKyNmbqaOPTdMXUl7qPk
oamHXrAzt3QgiBM79ZxgX22oXCUw/2J+uDscIvuHJ4P634xSD3X4LSS4Vu+6CqvjNbGwQJL+mUCB
MNMANxq5/IL0W0PnBmpNVrl/j6NMbBpS7V98NZlfwkPugNDqUHtu0o/IlgWrw4rWSj2iM1LRLqNM
CeD9tadjle8HkrB4on+PtVuX9myoKngeIeLkkFH8uArjDzUW/8cfZHNJE1S9eWxKaTJb/gSuqz4e
s/1GUmW1kaWgJmI3yhdrC3CRrWKEHdyxlAfNQ5CqzJkGNWURX54FxjcoafHzBS3tj1Sk/7eXdzmM
nhkpjr3zdONl83noIuMKX0vZ1l66QbZGOvK9utv7/p06LTQ0G6ySF+s4KpVLY4mLLbvkQN/3KGKO
8CBoewjqDbVRVj8XQh4rpFuWGH1X1xTX8MXUiMrTKk+TAWCGXdzoi8emnORb+5CRVuLyPU/EcyZx
klVOK1l0WkZZIsIIK4QEE96zHeuzCqJh06s3W1Ln3KmHor5NG52XVs6qNmiwVjceBrRJMdc5xzRz
xlHa+cBcZi2CWyg3IvOmzBvrwXQ/jDZTN2Ek0Dvn5LTT5mxMmc9saSylgD9PkLoGcV7ifeheN1UO
rwSO+w3mcrBcWisLaQtGIAE4SNDCbFB9YWnEtTn+tArCbWKmqZDgUGudi1jeWDPKN2cyYRMuOozl
keTS8AmahCWUXUZ1RCrpoSLru2uwIQGXdmHCU56QETmk3o1SOi0DE6SCR25YS6EhbIw+2AyN3OZC
mKNsTv9K8DIrwtHuCgBQ550kLOdvz+rKGdI2ZeKaDHxL7dbjkfbZJt2cf0v4ka6WdR453Q0fKBsQ
9ZVsSK7oX3UlLOMUtytZ9pEjLF7WwfIGlCzGpD2Ya2xTEbATJReQpeQcK2X/Ko4bDo7+nAG7VsaV
ubkgDzrBYZ/AfME6xoK9O6QsFBRUNgDkfx2arcif7S8yB+CKS7pwfkMMRVHphr0vL5GF0m+5q9LB
R886clwggotKDfFNxU/aJlHsLPrG+YZZ1IpZHaQdIk0W+Jfp//s6VoAoW92qrUlrgfZoYG2tS4h5
0EDoQMTyDi/7YXoWwqlKHvMbXMytcWVVv/ncZkCX3h8yHgFttv/fVZQ/tQMRJ1IabSpw+X0Rq6RF
FilB9KbO4iiuuvsh920ON4n2VRmqzEBs8T/KGr/t9QmaQnRlM2ARNGhcxaluP9KjM7Bq0ip186ct
P1e4qJzp44Gp9FICq4mxJQFxCJ2XGafrKHVm2/qv2/ycFDIh7HHuCpQeGuvGKX49KYXf4ftw2bzo
Kr/NqPdVusmVZcHxaVktX8tyl1k1tLmjh5NDcakIeWPiiKgHzgPzcDzTHQ7EJDTmK0fyZZ1EicII
HsPADXi/vNPFoxti7UqxW73VheTzrff6trFUm8He7P3AR/8J/nz9ad8cwDbWnIAgLsaF6Wd9x6AH
jy4FCU4FLfwOaMBx/TSzu5hL0auH24y6L/8DrQ6Y3vGy0bmlhNwZ12JMNtnKzgNMaLp+SZ4DNQv2
hXpijYUL1yqJPJoDJpyJDH0RbTh5cZ/AiYp/0x1aCJsnzUrwYLt1edlyhNs/aPEaL1dcE72lgwLc
4tXjJjxtVCxw+wD89LJiLb9/pMD+Ke3UfJDur+dkWx7Y20jKDCivQHBHEvzNEgc13DpYXTlww3KN
6lnv2XPpQjz4Kb9sqlHMMCCu+eaoExkt+mfqLkZYkbXaChGItXs2skvoMdeVP+HCQPE5b2zHWHiU
3Mg/ioAX5ZL68SPpUS4eW4Hw51mE7wuhydYn/eoMNvVIhmu6NYTJAK6iwDNDZZQKV/QT81Ebs59i
SxxuF8es5P26rPVgv1G0RX8U+nV/NrbGYtOj+s79MmYpeTlqruP3iU1YYlsqPOV6b/x59jlwBLzH
yXwmiL5z+tVWM2O53GwQf3n0nNja6B7DtnSl/a3YbcmDhxVXOhjmDK0fLh7ENd8lzXx+ATXJUKB4
NqMj9PaGIEjOId6v/HTRHX3IfbEjHLbKA58N60uIMjTM61GJw9rEWYZa7x3E4qFufjKcTTY6REf/
IxsGBTRmeRgjYkqbWlRIYH27ifrZFYJcEnqTu02VWxxYmgGK6blEMYwwVtbIM3NFTa4Ebi760DlV
5KlX/LqcW/PGlxc3WBJWHfhAwJSNXqARRvxAkPObfBTE5J8ycgQGsRbyomL1VETEyiEEEGsH5ham
r3PA7iEgQBmYNbzMADOO7mihES+Lr3cyZW4TArk8hZnw8eCNJIM7jIaQ24PAu0m86c7pOmJWGD9a
T9raxLwe4Z4il/3b49U2rSeRay4Gj9ITSmDmjUNo+lxvvpxNRrLAf5gPGdAUlhm6hXSNeXpgzjPB
Ckak/cJunAxE0l2dw+tDxgh35Poz9e13rLS2FyS67fntACpCOu/so8uGaC3/h0N97ILiePQvBM/9
JEBvuqWSZ0tQv7hniYz4AD1tlzulMnnQOmiSrbCLfiJYGEEIPktQFzAL13HQm7Sp+C5EAwB/kYef
ouT8gdXQLOUkbFUfzzx3M+vconbJJ5GG1aGkkf8Jw9zISTEE3tSnbTyMhn5SlEtqDbQO+wPZkna+
uxzWiBJZ4oxuovB5XQPC30BnMbsiFx7n5sA847rLPEyW5Is3uOorSE+wP39M2IwIAJIvzFwEMH5Q
ISV18cwD2N9kP18sDkYcU45Zuzd9HdZVjPnYWWRznzW9UNvRXLaynUg+pPfD8zhvUO/gRC+1Lv2h
aLLVUh1p6F6/cPER1gJ0fR8xVvY/NjW/M0S1lQ/ucQeiz0DzSL+vkzTEbzI462/dz5aQL6wmjfL+
7dtZ6Ihg8GcxQkyw3EmQYthVCU2X7u1CaVXLTMmPN8Y4RMWv7n2bXBrtXk47lG5O5xR/BnSyJy7Q
WBW8FJzMdGHYti5eqb+5L06xko1vkCFu1k5pGfgF2fHNwE/KYzKNDqtegahUcuD6KrnV23uSq6rx
NtUF8JLOH3Cc7A5SS9hz/Pxq8UJYPuu1KNzaJ1wmh0tohlKCAS6N6TSb4gg5P4/CVKZ+Fg1Q7DCM
74J59T+Ya6Uo6Ffiaq6zR4rcW+BAnQQ5Dfrkn68eHcN7lC6TQoQ6cF4l/tm4ebmRhAksDak/wenR
JNhU0XwOzJZ3En7UCP1yQvEuZ/IOO++CPt5lfzXI2ZMttD7xQHC+SSM28iUDNhUmTXnmwIKfi5QI
TJqtfTWWouo/FcdtbyoLdVXT3Ca7pdVhCdN2jMbUDbUm1KOM+LPYzpfrijtH66do3stPVMDnOvvO
h1s1OOH6QscgpLrQfO7oRajKUlKvO3POG3a51mP/FZr/VpcCZfXpHF7yRun+mhfvlrxTrnZBW3Vy
XVtlVCaG+RfxtN94DdYmoGVE9mHprqAA0WkuAMAGfmDOgCXjmLwvU45fTU7UZoy6Pco8wujRFiOD
T25jKsHCTY9wZfBqFWRMZPk99Y5yiatg94WLVHGPgUPARmoSvB8HyZG5mlDPyYW1PCvyoZxiGyC6
yGoCYfoD1BLQLF5O27qC8V9cs2jm/E0NgFO2lIHEUbxGexuq24C/2KuP78oNoL/NQIOQsJyTytqm
d9XMkG4xx/RuQdh+dYk5XzZ72udLuWmkE5woaaEKlxf9ufmkyyXsvYj2nnh6G25nTWvWAzcA+cYi
+3+6dA8tMBReDWoXNMz6Ni5ccfBHcW3P9VjqZfN4xMgi3utBUHrAwO1L/lfGrJKQWNS1sYbmSDgf
P7trjoNxi/VQHPWGeVMMonNRcm+M92ZPC5NejtDT9AXYVS1IEWe6qZ/RlYEEE9EoEH9V2BkIgkQ5
sOL2LygUgeLxRRFnGfK5Wc1HRXih4OWhY8mmKglavVvxsaxSs2Rx7opJcUQ2RlFpdg9SnIuRBJRu
LDTxNj71phnUCw1Qjct8RpHVt2QQR8JNtGBe4o081QgKAfYTvim7zzBXpr9kv+WDjnAsMo/ieeP9
AIu8vyIY4pL80xH7lGW8zPJ+J7cV3UbTwkN68oLzep2Iaqe86tsyw6kYUpt5oSID+bGYOHqLgLzQ
2w7NtUlrt3DwqVTPKESGQMoTR656nLLQFpjHMQm9PQWmNbYNN/yHD2pj9hw4Pr4BIx2nylez8g3c
3d5eF+LSCSlzPTMI2xky9yeK178lwr+ZPYSo95DrD31FH+hEWWnJ2VB5kWVw1g8lEiRBY82wfzF4
6fyUQBJFMQOrnOu8zAFL2a/OCuOrzNhwFp8TIUvKP4Sqi5x87zmy2u1XyyKiYobylopy6Jalxm4W
QMxJLWc63H7JDcYGil5uovkqDFS/fEkz7C4FabbPB9WlCGKiYKMDaGmw8hduKSUd4FGBo07U//KU
vMM0nu8dc8YS5Ja3hfira29fHzouCYU+cftvXbfn7lhVkm7jdhFc5t7tvs44ZrnUiPe/cEhBepMz
hS/C+HEQ+ZsJ7cSIdAOZvE1vR+xzf0+OT6H2qBvUYQna/dcLqfo+sN+/1gWzKiUK2zW1Oe2ajGRx
5UGPLJnY+xqIXoctNN2i7Lz1ViJS3Ij/kjAMkOzHzKTRn5qeLO7N2ZSsl03vT2pEhYPonX/yHZmI
I5g9e2ipQGYNKtSjbt72UKFAFp8qhY22/Gzm65ce8jgUGpy9/3S1EL/nr+0o7mwOF7X1Xb6LejU1
OWc2GBUlvGy0raYgg2f4k7Nar8TyfWt7m376eJ+crQVrlQzBOfPeaDC0qhw4LesBUkwIdkb7MTMw
KvuZ3CTiOklLicqHNKx+o93X7iNIJ71hqIHjYaAIh79c74Ad9oSr7b5w0zgOlsA8Cg3zPmscEk4d
jW1Zbxtc5KqkyaQux4/g0cuDrfWvxl1Bg4VHFXb7zwZrOmPR+CX3RDTFvrH/0p8mCm0SGpwyPbjV
hJrRrLddY/cW2w4+rJO34djHIG1Ss9l9Tw3PnFMUfZxsu2VKRq/QhmLMZEcmlKVvB4fCxbT7tjkp
EjTjZV3rs5cOvIJunzZv8r8bSlxtQl2Tbb0AblfUm+dG62ADZFklc0nJxuVr5ZeVclznpaCnRtg3
OuL8SgkWSYZv5x5n02WQzGwcEWDYHHwekTi/ryJYpJb2MPZawKwzB9UVZP1TCsCWMXwSQBvXRqrL
qa5PJAhN4z+icLQKPxyh1kLd/XXSbJvlMRcYZCevmR7kvlj0JEWMeqjrWlagNXVGtFMwr6gpScaM
pNOaWiH6YX3Zmo3ZX2OujOuwieqrHnLlrC2ybJ+xQmavGqVeAREIjLQkFs5gvNqmoxJF4ihHV9QD
cRjaWp9iOaUvN48NM/+GQ/C+SXw7k5hG466juJ9IHPcAWhkltXxxRMTIEIP1KRMxudBULTSUJc3l
7sieF7vISF1oT4nO8XfuIlf1hQWSD3sFYzFjIwtjcHzj4on3mKgOyvoRuyS4+DJjn9LF0giwE+lf
rHfyR+DD/TteSZ+TLDMR5onRKEYrFK5u9KIcoKfTmX4GkTbCHZ14uxAENCf4tIom81GTh6Xekpa4
B1rRPHvhWZjZbhZShngUUiEWQNEmLrRoIOAduKjvifVEXhqeIOlKe+LNjlnGWxlHxOAmPYHB/wiL
1WEIru3K3qIkIvqfaOVuCK0Ulyt61LRvrCrcxv48Oqe4NXplmPbAlvI21NK04dHOqi50REv8gvhV
elBxaOeKSK1WGk7ThYa/fRFn0dJzjTXQyBrc/URUDIVvSewnMafAqCSJz2NLunv7dPfK7TYDA+v0
kYB/EUhCQJO1ePROs4iy0sMMve0aab45vU3AZtHjkyb+9qyhn42/NAW5fbtXBg0Hesu9D+fD/Im7
bsK+SeLvYI+6OHTzL78P6HFY180Vrqa+RHGPkyjiE27JkQ+GtYUUMJKI4bP9P2Bll/Xh2/vTCqaq
6YK4Twg72sM28fkjYkMlAcGS3izkYyheOZpWzhxn6knd21sRIU/++kGom42vkdtXQLxnaWE+c4bY
4BIrQ2OwGy2CwSYv8izzwrnh6djuqscRXf9vuiO0FR/cn8yoYuEn4LFL+w9+Ebf/dNNhI1vfArIo
7/3cXo6i9KRC5KN+lOsiS4/M6V3c5FdnqhECw08Kx1Jh22VuG0AVbEn99FCzF0lgxNiA1oEj+Dwj
o6oDBz1jHogR0YbdwXkZQefK+ZDwFwDIob0qX9X1PsoD2R+FzRhPLHIIXLOWTOmdEWafIVseWB5p
tnl6Owu+CaSFYMduPmby8Yg2FZBjJTFVm5XNzvcPybze403SKedgk01ktn9HT88fcR67VtTFwTjk
JwUKHg1LRon7HMwUOfMXRNUTXKGzul1zksDbhxBrlxyfHwnbnMCVRpFPvdAeekUO+oRxnHEZITKR
W3aXN5B1eBNUvujn/71XfJELy+DbD56QOogIykx8mZca9pKUs5OjOtuC1+wj4ZJK1heRQrhfz7nU
Upv6Y8mPhxQRubxbrVz1qZhIdTAf4Yw22AhVXjFdljR88Ymfra1kx0P/EP7MCJ3Qezeu0K695xTa
8cZHveHiillgtdS536vMJlewONveglr8VWvtrCcK5jlNAe38avgdTOJUAw1Z4h/fGKNXsHtvOEud
v4qfHKJdajzASbK1ocbNCtsuzkyO5c+qGmcuvG/in5iwcoRy+zqDCrL5Dk3PFzQNCsL2CCLkEqCR
R+PerwKsxgsnL9kxf4XSgPNjgpaM3wHjJG/QbG+PYf0WxY/za8iq57iZQhshJal+kygW+CqVDWdB
wqTsPACHrstLutB/NVogX6LOjJlnVoub/mn5EN48rJdy8mRVoCCaAtZe/BpSZdmlHULLnbDfAZB3
7xTXdJATd3PRnTDRWRBeJ14JNx9H2A2c16hg+NqUXh3nHKRvyY693BtaLPhvBH+5aHmaC0m5FTDy
4bS3JAePesIYdUa82wNiXevZypH3Gc/EoYJdhett/rr1eD1/nQyv/9l84SwbSVKBa0+XxDFCynGS
ZuF+LgJ9KlGgjLcHwSGgcXtwSz5TWCkSigYSuMC7DDs9C7jRrJO+fT3brmeIIfm7usEtMx69Uz4u
bU0GDG0bbRuTtKnv3zanAxRWF0tFwm4B1LPhK0rP4vCzbEFPfNG8XhLE0r+RLWjqr/30FWRYCKoO
VzjjNFzMsFMDciALClZTAqnYqR9YOcHdf6PmIqKKDmuNWLDcLjWaVbge0GikBgewDvtK1PtEWNLe
vtVApkMhJuyg2jruzluI6uQI5hckSBTWcLHLUS7pzWvlytZrOuBOUtO8yui/ENlI6zrc/D73sx5W
ajBbnUsew05XjmsBV5C8nOGe9uPF0bHldupm8AFnTXGFDnVe2R3bMsB5WA5BhyziTD9Z5l6CZMT1
XUu2vs7ZdtEQEQZXXqrz0n72GYZKPm/72Git4ER9Ak+wekVrgwUtkIhou/uyMAykU9JX6lxcpFMB
xEz9sZ/2EtadI2KBtngLipTXlCwXj+sOgNvy6mcDnQH/G6fvX/14aTHgG3wq2CszRhF0gLclrO5S
rRWH/OEZS9VA0YTBcEnoQzSFCxiCok6MWgCN8Gc1hqr2qpbgV9YnEgGyEkvnmd91lhXDY20+E6TC
G8ELASiORazE+0W8x+SL26AxHqHz+y48phGT5sFkNtD0jkfjojO+ISZeMBv6pQ2yPX9ry9CK2+aW
dC3vO8ZhdGrZbVbdJkxZSSThCyjRLp5pbdx4OeNxj62CqH9fJnLHxO/kKcMScUHozKwzcRVQzwcp
8vTUVtg/32URwvUd1t6wiqS4ChqVkRswGZj22Kh60TTZny/7po+vKcOLMufEIOp8Fy3UZCApZdqB
o3w36MSr8EapXJR2aO+TJsjeHvK6Wua4CUqZz9/1Cju1eCSzhoosJgvF4uzht0qsgrRxfx/NQfWj
JI3NLfj5pc/ZA81d2BFrkVakTLkBJtPxHwTDfz4icM9IdRCH9+wOLkrw3aOKRTBmW11uT8URSJlv
+l65IK+YRy4KIW3p/kwvbxBITCY6+yNVgC79OreNvn4HtqIZ7REffjgmYrWVaCfJHkfz34SckZwr
W6rv9YdZ+K2o49+vudwJtstNHLJXiK2VZp5Mr19xj+roe9EaR9nD6gM7pAPtdkTINWRnW98bW+h8
8XDqqJs5ziLjMYJp0ad5qgv8CYaxGpMAEhh7r2fyH/6GrQb0+4qPfvOU1vSref/TeYEJSzOYQTy8
SCesdeL6FIcx0p+1qUaZZQFjyLaRS7hqQLKS4ThijXr7YgAtBlUsXDeQEgiEuu+waBUzmfbMEkck
KPp0kjoWUfDCXdN4kqzsRVd/G487z1ciF0x7NK9GSCNzsGbsg5z2cbhPhAtIAn5hJdjlLfu/OIB5
gW5SStq9SLafqwmYyT5HZbrvGRYkWh7BuGV3/H1jFnurp1vRvHp5XXvsZ+pNWOK115ncUVEuXEoD
QubBtrjHdo5GLV2TcxDTry2SJ2+uBijCBoM0V1jmYSlk9NiA+74OhtYbTe2vfi0XpdcGV7sSZp2w
ufm9wNwR9yUBiq31zaYlSIpYOl6fxTowOlIlt0Vi8Gys5Bwjvfvd7f0wPLjZcJRkqvtlL6YDj7t5
n7WNdBxymU5oQMdyPBjqPR2mPDtznOKfo7PB+ZXgBouHPLBG54vZ9qx5S4rxb0QOu6ednc2VJrUm
DvGqCR2lVdV/XKXyeRmoRGSOt8d+KZDC9RwCljI4UbSnD31xe68U8Yai/mY6NfcZ5z7KW/oSSDzD
H/WSql4a99oyhCkceXngs5LIYcE+11+ITxncTdwI6ZUwIgAbrCeeyFpBMHdR7Cj/L/VcCAH8PgiE
+2fQaauovRd07gIla2KLnT78Ro/bxuxyqU637V84iD3fRSswX0Wn+8VjFd3PRg0me3BDd0x6PCIk
o4yQ9DOKWMQLrAQPZ6+SSZQZdR8Ov+yqkjT3ADTE9wxYOI+vnOq1lH0Z8F7Pp+KLttwCp5goxdqd
l2b9Tn7M84aCatJevEAaJ+8MMOG9AIa0Lg7FTs++Dk+XbySvOnAa7x3AvLAy1EIDpSVqXaDR6Wg2
ti718yd4pCdnuf6hgJBaIRLXUcxA5ufu6X27+zyPfAxfYz8CeX4NK9+JCZg1p9eGcV0yaZqJfDff
OnyYoVqSe72qiQk/7IHTBqo2qdwTIclGbZMGYtU08e/T9PLvOY4OAOZc5osRFiXHvhYgt7vJT6L0
ZJlZl+7ZoL3zt/rAvAG1ZUNC0VmEA3aOSoNApRbmev0W3snyXvXww8ggH5KepGgYjeWK/B3J8RFq
XDLvvtmwgYLqgIZX+IFZGYwRP+B7dOuYuagBiuU2Kx5vpcNnIHRgsGWaWIbhOvtKcUXEfw5a8yRA
6Cb4VoUVAGVrXWvbwXHlo7dEwFxlktJDxM4yqBgWN+gPtaUJ/2MuJ73b62WZQ3RpLLhtk7RIPudK
omwCmTVWEoBY/NTY8mFcMrSOFNw53fVyxP8x4ZwlO4znqmiH2nQD65j6LPpcOQbOdIkGM01QSNoS
uA2DsBWk0bWb144GbEazXLcmi2j8M+3aiETDLVy9LiTJIHdZAKdGEWOqUBucEzty+6x9bNgcMq4r
z3EgX9nrxrLQYbOqBHeLVvR5O4Y9RMMC9t8NzbOIUS+SXfH0r3d4VxUOP/l88OpHpFCn81vMk7tp
7x7ltJI3dPC/z1bvUmXrQddYp+tPubmRLJ/x6FUPFN9els8XwfprO+1Bw67zQDrHIHWyUZc/KX+3
xlvbn6x1Keqst9Akk4htGZOLoNA5cT5YyXb3jeA4LucRbRoCBW/DzdSyuilrdXhNY7ev+KLH8v/G
DSR478bZxuz/bLuWyObD/AmM3wihtzY8wXbH5h2wQF/ZEnUQNoJcxRvPDlyjr6vYHvHhKavgceaJ
SIl45O5leRJqRIbvboW8hRvZyMI5Aju2dD3eLGWHngcuCLxX9jAw+qwH9SFfF5bnghRE7/kLAS84
DCG3ZSrPJYI40P8xC9g6pOx5pXuPu7boGPGuZwyMiPmSOl3p3wD/vUtPZHYWAMiBLRyahutRTnQW
/sH9uH9ufgHvC7zFWN0e5eEdAyWij816fsqBhqCXd8aV7SoeoEGo2pSTP4+TCqR0B32jvrMpdAIV
ZkH8eP6KC5jlwBHV5jBRPijWh7dMD4kQUNxIh/IXhDhz7JWSSocGA1tRdmPQsPNCiFM5dIuKKM/d
2Oyg0b8k96qNhznZzXh/p0FaMSc59FTOoWKvHUZmCmcqperU2l0CcWK3kJUfhHLMdQ6OK/OxgKGl
Pi2E8rNYrwC/7kizN8gK37S4PyRrdgmtsIf3YnNvMdxCpKve9UnBnTUmhrA13wcZ4iuNwisPPtCk
ninxIrvFnpVdhbno1MOLkzxnn4j/ZL8eVE2QL4Tz1ATP0h/RZC6hsNKOzGlaKioSLLEMGiTr8MFW
vKujxkd4BOYNNIPw9kGwKA8WMyk8EQb7BD7P+A9rEMmf7uIMsrFvkOFSYhIvZOSIW4V9n+VyIBqD
Cvjzccjf9G8ZLrlx+9eCz5Y07eeRznXtDMA+kQymDLpBxGUW50v2rlvDVHYFLkedCFBz03w2j7GH
sAcd92qspn6g1M/tnTeyW6Yxz0WL9P59H8yX82g8CmtoNAMvJj+EOz1AvXpkhzhhXOz9+6NqoJBA
Ie6GSneV+0p3AojIDJis7lDJL1hc5BxkAlGHPismUbm7QsC4bhh/eEV8n2I7vRgs2mh98eT+RPER
bgZjEQZgh9o6VbJeXuPXB4XvCym0h6p0K3mqScMHTHSL3797Av6HROU8GVQBWxaw2fdkJsSX2cge
yUlVeO8UcWVXNFYpj9yhNjFV5px4/IEDIH8MDlDk2P4/DPozIS+CvumPaBv878naGOtPJpJA26Cn
pAv4FI+EpX6wNWjT50gd9xY+RTCoZXzD/dKsf3cN0L6qPWDZeKOjnmyiOoOZUq3HVNVV+D1638YS
/czN1zi2/gVOoN8VdbCS7K21lrDTIGSsWJJ3CMPrqSGCx5h1U0ope9xT+v4B3sS5VZnJFW8bfX5l
ahWBvEMfg+q7mekIfVRG0NIlggajHqlgIz78wLwZhWAnRmDxrjWLrwNzTgAygScu/F6WaGrio70E
e4hY2IOPhbAmTZ1kdkth4K3vdo62ZPJN+zPXF6PvhotUe6qgBfBpVSm1Tn1NoVPdQfyBVbcRFddo
NA1g0U6X0J/FKf7p4Yrm8dQCLrjB0AHFO+fVtDnXF7rg0GKf/TBgGKGm1Bua/cH9he56fxKmjgrg
qfvnaGM2nn7LxvHDF6aiwNOyU6p+6HRIUVNF/ExS4SG/bIrqzKibrPMv0QtkCR81jc9Jo4IIWhGp
5zy4lQsK4TgkWS3P3aZXusKtZ9XwdLh101LW0xhJqpgRNaKO4ieGWn7/rFqaaYRByMc4Aq1nGXmO
yyvElX543wJOeTqI0NkuHpd55uqwCOnVhVBDOlzkcqw/g9/ZbBpo1RntAyVh/G5z2nQnm/B2QaIS
LAydDUEkDiiMWU/jhBwuIcwVvTBeSFtOTRARVeNFxpdqvFc3MyvNl5dlhuhGzs469+ggM2a9MSWa
N7pT8yAQAygrGh+Kdlmcoufzwh3J0O0mrjyX4ivtOXsSy7FNh5CRjLI+m5486nBQKBzr2RYr3JKm
xI+DLhX/NwNYAaM3ZkVEViPxFeERvE5YeOB9C8Jz7NnD94IQa4S5VkZFbBfUFrcUuHCNej06qk1y
boUgcMi8Kcuor+KbwL1OSxRkjsc+8DiUIgPh8fMZ+krlJbvyOZQkky4fxHzh/zyRcROdBpbyy8v4
6MrpdZ4tPxpMhRz3xdD/9zYmCpxdl2i0A1CAmLSz/4b2vgCaB9/QBGkKyxHqZ3hdtU7/gM8nMQQd
BXtbBHGZFyx/4Qms9y5SzqDdXMrYXuFKA+CoAFADEy63MB6jcCwydU3wFeH7fSXFeZZkQTIoVznn
Xyuw8g6ptyoLamw+TEsfVfXoA1z0sOzjOIatOiGVKMd6YWnX+fMDX6zEDNejn0EnoxhAeP7r/59I
yYg+BOR63zM3GbmiPXLxL7oyps0O/0M31jgSHw6bYvFJagcJJUxRaIzz5eAiBlMbA+B4ukIxb9lB
c9iMtiPa/5zHuUfXjwkH7d51moWa1I7YXTiv58Lt/b7Tz468X+JRHSmAdEfV59h5Ectc5rYWwyCx
hnBIISRfqyiem1MYKB/qI2IEHO2uwTfkgVWESwvSrALbx8f+97jdx6lP0LBvmUth37sxwNHHmFU6
P5IBRRFtMWpXSTx6XMYT2OuhM+evjzQCUge0e8o9yFYC3pMDwxZmCltRBpOJGh/WVpnS1SOvE15B
YmNi0Yu0yVy0Q91h7000T77X9q0mPbNYu1/y0iEMf0ewEadt0/+MAC4hjpvIXPtDdj3juYEBqhnA
REzQ8GrXZf4nszhuS5fFGj8p2dZ/XqQ+vQVd55K7O8QK0Bk50iZYItYTG1B8ExnHbBXWCOmYkC9y
/vJL0hdQho5AMdbbEAhXWFiuR7ZqVWwQgr7aXb+m/kHjrMTjWs/DgZxHW2/LmbQ5PShzaxFtYJIT
FaftuiNd50ddmBzuYjYsWoBlOQ8sidndQnybmGFVdxRXemOoOevk7YmmE31m3MFQEYmZ2iMlTLFP
6E6lCeI94l7UXxnyuk43vZkktMI7KOwyDFnBTmANHuGiqDHDfwQYJ5oQvSHNl0KJv+AIZq0oNvz7
/6nlRq5aIARmQZNaxrIxr7aMrkEOfYngA2pdTOr0NB5bR0tGc7bYuN5sjd3bRqOQZ1W/0TjtNn7a
iVE8GyD5VDpZ6DMIde269IE1OhjfQYEzhg9x94CjwubHMpm4+8vsHb0mVeDt1T5Nji5Kf+yqHhGr
RBrKszj0h1DmLgGYxJ0DsPLFnl3aIMpi/hHFThvZPRGYqeOqzM+YZE1pfn3gE/sfyCDh8b8iGDeP
YGTYjXeUSQhpQEu/nsJm0iJnwCeh+Rsl2sX75TUYzoYqEFJtcRmrBdbc3CL39wdb2PSEwmTy97em
G1lUP8wc0SrNXDuUyTiEQbZTANm2mrMFU2c2UOS3C9OPv0KFSNUVX0pptLBo8yfgjqGzxbjCh4jZ
RnlD7OOlmd36WKYWn9jN3vktuPg+qUAIvJ+z61846zyRmFmW15patCWrm+hBRIo87V8yvZwGJ8Ko
7qdd3p5AMAIAggUiQYeTp57FF6mzfBsfqUNxYBVfm34fbYAkpYCEjzWpLnNi6JYXuYa6MwY/CP69
ccp3raU64UsR0r3kPMpnJQcTunlBsspV/prS/Ma/Uuiwfm0rlZRjoncCnTV9J/JdXZ4++vkfhxH/
eBDoj7xcgpAk9dZfA7+Jhg913Z3LQieBd0DdA59fVKkIxP6f5bMQl5TxpU30UV/SVdzjvCxCxVlJ
GL1ESPIydN/k5/TO8SI0UZaGiVqYcBMYKumc6JigwJUrU9aT0CB6bo5Z8tQ3+18veX2e+pGon4hy
yilS4IHUXeAjkjJcIQ6yviXB/F1CNUPbCXvO3wIfnXxE7EFxY7KlBuoga1HxEELOAcybUVJphguK
w9IAiOlXIy2Oxp/DRV9+BL65d+TcDnUqgIUjvA/KV3Avmc1VEd3Cz4A4eA0eiQn9VMfm+KLvbIiY
VuWFPxdsMBoU2VB9fXH73VZkp7DQ0AJXCt5uQ6c19dbvEYak+aE0fuz64URxvPoELPv3X2kheV8A
3s9zxqqL1K9Z1n1TmnuyV8XLD/BPAGY15YBjNN1FO0FFu1CtThPjuLL85KtRBEPKaliEgStHkfmu
FopdeEGlim0VoS5XSUbQljSn7nMU17SAYPJuEThQppjEReIwOQJJJ0yisxxXdcp7jUDFzbql/00V
4WxjRErlzVdDE3+2psZruk3I48onMw5xSqaKiHJ5IcQcncPKNCVi1SIUvIPyrF5QxmPo9JkpJq92
2B7M+InvaoMm9/4D64H/FUPxGaKC0f8KNzTZfsur0Vj0WvmgNTpAm1lCgxRspUyH0B8ZVnLLTZsN
fTOFOCftwkXJyoc9Cvn/qtdZpjVt8LNOD8wcP0lfvEacbmJyWinVhGxOuV0yEm9leLOwWm1HF/2h
1XIJJ1mcoBFEzW8YY/zvduUuR55KcGtmjb0ejSmIwgdTSBUYhvgVIeQG9hy8q5DgyHv4JU8QMemu
TY30yKDs4q1LQvWaX8bIt1uSbpIQp9/3O2sTnEuNAR561rY2f6h02lM9DFzf7nMuDlLXeMoiIOi4
wQECGEqdZRWE1Dkw3vmfVr91La9MGcwt0VTLAt1Uvk39PfbQso12ycmI2jwCvPF+ivMjMwtl8d/f
jtt8VVVYwh/evnrRBy4mHJmkBU/snPEDRHazXb/SJ/SoOmTtbZOPVKEu/cpsDvT2X3TI8OjgD61J
c5uv6zXIC6upAyuMoV38+49L1IOoKPK2XLTdfI7nzyzrmcUHI8LnrLzb//P6shoKJCvEAW6hEf4O
ukMHr2aSfb0t1gtNNMm84gJUwm2YXqqqba+PVdiPF+R3ucw4YJa2xL3n2P4U46z5OU0qadPRYADj
uqjP47pC3V8X5GbqWErQ+WykTGHSNwk82rfofnkX2iWJltgouF3j2/d79QuDGeCYPkAvSMhq+Hdk
b0kLG5WWuj80Yv7hmLkvFjCEEymc6/pNtaSb8cvCRVxKdOjMIQLdyLTdr3NSkxpG4LQcDBg8ESpI
ut8eQsEjTnwRRhp0cqsSEbY0CxMi6yqd654hYUw6I5EVNTjkdlDk03Nvnq4hTzcris7ihEdXV3+n
lFsqu40WM0z3TU3yhMvupcg6f8hTxPlY3U+FM6OTHPZFezXutO3bX1sI12eAtINl2RMSaHs3BcUV
RISj9TdKjU/k6v6HbvhILEI/YLjDtqK394QjL2v9CYudoUBl7pZn0I//NkihO/KBeFPY3rDBMeBG
E8zIRUtt1L756t6Bh1o9P1OTHv/PceLgpeiFym8cPOGmtLzxuf7AtvWTov4WNbR2jyXWoZiuqoiH
JpNUPiEv8Aav+q+H1qRpbCRg40ZUGZyYGuhCpxxQ+1hLd2pg7s3rH/8RHx35SiyYsuE6mhxj4Ahh
IRjr0Ucg1fJ6dDe5dxhYH1o57XSBWJFkKHJWUgcdhqudPLNhhgcYpu8IsbJ0DXm9Z0hu/jsMD+Fa
hPXvagsk3+XdY1BnYIKVoxDbAOJClbowl7EjvGTM7/qTJZFdJlZCFd0yxu4AnLBivEkRv+N06Z3M
tGzbn4mZfnIeLT7KUdU6W+Q57N/+aHL6IEx+Nr2l8hRGVLxTU/Oty69HEOzQD9VYqWabe1hWhwhv
zc3YjOgx1erCuW1/6THSWJ+n+nRVlemawpGzECUy5xWPrpI9vMeE2rcSq5yILpBDP2XjKSSsTr0V
dedD8PQIHpnrgvbhXH8qVbjJA9N9437qOx0sX6Ob32I/cSQY+8/GQIXXNntU5seRwVMHyLqiet0S
jMu+l9zNeL6cvrf8RJnxXi9DjvQDDpgefK0LVPuA6wPz+mVSbcYjNjrFnnXA8olq7NqPuIHug1hP
iqON3jlEZ1XoydQtt1kgOLpYQv3sYbvMOeUWuhqVY4KWS6RqHbxd8n4oqf90wOprL9pCIS1Lg8Q1
9vb88luYAd+z6oQWe/S8OhqJ+/JZJS6/37ImAPil5yLFLj3E8o6rQrLV+rHY1pgzGcFDWtxjF4fw
O5KFGBjieEnLS6NFJpOQa02waUwOckaqMvFMQdu/B5uKnvVYRUO67bWsri/P/trscN5RrsPXX+pL
xO/l6q2/yPhK4amHIgDjFI4b7buZevUUIk9IVIcqnkyYU1hPx73BT/PqaPXegaE8lKS39EoKaWLm
0vTzDu6fhoAO/kiINSXgkrE4N8UAbrvAD6SRiDW/ptcBSxlnDB0Ty0gm9/2BqwFDQMQ8DUQthUum
q0u42wUBqF/JxjzMkXKxAXKovXMiZu++kCyEUwHcGx7i/nuDaDNqASwM8JDy72jfnMRK2ias5AAq
X/WagKD9K1N2/3mTcy28qezTQEZimRAEKX9iJ0AewqTYwCzs3Xz9etq9BXF5tq+ro7g2/egg8W2J
Wkk93IdgrTmP38/FXoXqFy6B+ECQrZA50CVKUA43WIGnAx1OA3Q97B6imUKePceV4FFarCnnm9Jq
KZxguBVIfrcxnp2GT/aJJ3NVPpoR79x1fkcI/inGwJEyME616PTGtsBGzRtuiKCSp4ZmbusJ2v6s
u/mGeeOGSLk21neXi3ZqZpeZhi53lJfiSluWlIZN35chOrqJqW5fYqN6egBugGteftdVJ810JNHP
ni0tqY5Q8emahIGRv1gMIhrcd8PXvzWKSMW+B2QmpcLBRdTd/wkkKhZz7O1PCMx/DsAjgNHoZLFS
ONoPKPmd147AJjnRsp/O9XclxO+/f83F4wI0n7AJpyUBi5df/nvrA18YmZvEAL6P1KLu+yao4wgv
gKfHScHisSjvo8kl1RJ41mwzwFE1jivLhQ5c+YO7+ygeNY1eerSbsdnfsipfWKIsl5bTNXRFfuJr
/c0LP1vvZQwa1/77NybVZyU668DmoT1u7nBxHEEPLokWmk5ea0+a+Q8l3KU309SwN70c2ocwWolL
OlgmSptR/O8xh5e+pHlHPtVIq94MJjXAJFGQ0e+hhFvQ60ErMDUEtRQKhkcIhmnLijTnP5sbNqF4
yb8FJgOBU0j1I0FWKVMnjN0L3sO79Ee5La1LREWe+q2+9t0K8REq/3vPZru3ReW8jEgc/QkHr3yN
ro/v9sgqowGTpplMp5FxbimfIAFdl0DNwHkDyWPGE3SSvZe3K1Y3ghKgUWX2N6t4VWhsX8gr665v
p9v0EAxgit+maHRj7mXCUGpqw+Ly0D+T0iG+wWQHHNVVLINWz1mIkofYFDL5RLRXGZ8IxnvtQzJd
WPpsI3SV82JW+ZotHjEfEdUAFpEiJUWDbkRKcEPQ6Qo4W4ZDmAEtAs8iurQjsijL2fLUIUmJ+AZH
caTk820LhvC1H9eU6SLvJjPZuYXXDq8d1MdxcnhQ9P9FLOtc+6kCo4LB6/K5QJeCCEs3RD3Sju5r
4t9Y52XveriMRNLY709YYk8cVW5imb/YM0/zYlzZIJv+8nXM2r6B4sAYa9y3TX0hrEkEwIyy7zJT
9ZRJcSj9JvquXJNtWiqY8fbm/su1oj8N6HLoVVGezkGBXsvoLDwHg6lYjufokxMG11QJw1CT4dAN
48SIz4DvBwzgKelk/bOb+ZzkPkZpwmR2wWWnz2FoqBp4jekJMNd+2O6Ug+oZuZh6ahg+cb5D59HY
OkFWZPc+0Y601zd/wpKJtexHoXTaT6rbiKl8H9NOjCkLfGY+j4VP/NuuGXw24oAy7xn43p9AY7Av
G1xcLewlHxkVf/dn28/LiI6Q77xoiSvQHyDL0o6vTcpBajj68jhyoU/Yaf6usQYoOLM96hJkatTn
MTJX5a5s8RY1BgYQ8fipi6tGcIvT6v/lBldm/rOvJp/z/eMGDuda77yTrwT4lIHFW/0D3lCi8djM
aK1LejJ3Xc/j02Wc3S6xLN1Z2Fkyjy/bdR2Mr1BVztGCWhUQDYk11vifBjkzxN+cHEOgNBjDX1BD
7F1GUI43OQambk6OoOm8kwJzvfTuiq70AVGamn9ZegeAmIqiMYSjzpqIavW/85g3KqILc23rS33w
3y7aELi5IpLT5oOVzUirxGhjonJl11WHjcpxh+pbG1PsKzCRLuupKQyWrgD/pNaCxwn9C2n+sa//
7kAgmb9Ysay5fAD5GOWw3/9KedKI6kBilsQD8A144rzzier+2pXJEALnnPReYG7x+7CNb3biYblj
/JGKQF7sPMOCUiNlaZpZ+6yWjJg3EnrU1VJvf0mqYYMYwTZlTzn10nztZPNUKgfg0jdQBDaq0Alx
UxnDcmeslwQj7b+d4BbSBdQ5sUc8C21BoNJUiL3TJNQxYAmGfvyIZ6bcgMK0N7/5lQphf5PAbKmt
OrRFked8v9ulkhCflQZ56FMb07VIkq6JV9B9o3JxK7Sx67a66a5Z450qdsT0//2x07688y+aju+w
ngJY+DRHwkx8pCjqnjNbzmFzmshNOAHHJ0iFwfBfA4xi9eiVxqh9VR8wyCk6UpA5OfXmOyipN3TX
dV+OHItJwe64v/SDYbsFpPo0XjELgJPmlpeOawlcda/yXRYGrZ3nd1lVOqJOC+SZYR/qQFT/Esy2
Upng1JYX7IVCqmeUp9P0heyJPe53GaffpoM+MMZIH2AukekJXAx5taVAkhwR3UT1WrkhV89GeSZt
YJ0Nt9rV4KAVhP/yf1J6iRz7B0PXMHPCUWjm87yEiboAKFKYfazTaDteTv2gKfCzIRhU0iuqVNKv
3YAlb5JNCKFXWIPdH77i61CpcBrCMxsf09mefc416wXXRT5l+8p6DYptEUue+PhLxV778GnWAvP4
AhtrQePEkg+4GWqUMLYcRrV/pdPmZu/9YaT1HehjazWkeWIh4miwmZVVkPvYo0FQSDVeqzxGBS9U
kf8gIGi1xXefVPFXgLMz8hidghzjhF/idFRWpTk666X8LIiVZzixORi1s6oTMVqESdHJO2zzoOFt
eq5DbPNu66u64Y/ZbY2MmKZYUxLvSOF3xOfweot2977CE+aS4jOuboRwlOXrhfovF0FWsSxzECgm
xnW/y95otNKCz7fyvmIHHYCqYOZ+wSaqTqyNg88TaCYgsZV1v0FbtVbEvZAw1NUnJd9qhza4s8nb
virB4xGUDLPZDHehS5QPido5tMJJK4UxftGKqYZoKfvwrjoLJVKfjJpHjMN/Ep7euMegoxOH3BuK
QEo9nDBnEb702OFw3xzQeVWC++scaXogaiH5sAfU/53uhd0OkE/dcBdsWeUt/+WYiydNCWuRM74t
q9Dz+9IBFgJ2U8PAZpu7MLPenwhBcfZbj4TsPGBeoF4Sp8+YT+5MiZAfzATQj0/3VBUrOnKZA+Hd
tzGGrI1/JEaXJlHHSE8rpmL6+In+sDbS7ijD370sXC8RwndFLUWaqDLJo6MAijiZzRGi/fBolSrM
I/mwBvx9KE8I/jo90UIOqXtAtZH9tNSDES1WIg13p/fVoPIynhAZqpW2gRnjku0tFMwzK2G0JvP9
uPJsyNLYCBY6/bcHBpghhwquXyXDxb+eEi5mGpRUIc5IYFqB6J7ZMlLrzaadyO64g7xgVzZMRVT7
sN7CyAEiIBlmRHXI3DXOk19f+3EGU7VzjbJb5g2elPAHIRW3v6hmTY36Iab4CGrSE5p0P9isRzDa
wTOvhHEfXfGxcpwd5S+wvO5SFuBO7tTT8d3n21Efw0uCfsWZXSax0nkuwG82V80PiYIdAFjfw3sr
KLpsfVl3EakMocNDASZl51vOlw35PdReRekVaTN+Bt3J0Q3hz+xiApr0w1i6s6eYIf+CEMXe1YRf
MpwS5iJcojwefCV3hillT/nzl9MKCZfjFoPCsPXH8+o8RiYLmL7BhYXicKt6yUzzeeT1xtfJ+8Vr
3/jShJzuUMoe7V7eDniVNlHSYRZ3myTjbukWmAqpxvOI+pUkFz55VsepwTzzVUesvuF2g3UtlIHJ
Y3friPM+T4mnzfbiw/Wi3/iTHYqJnUNPqnMNWurChLpUBy+Dt8Zpd1LOIF1OY5T4lneVZi+nY2/U
K/UnrbyKZ6aw2Il6GruLJe3duZ3/hVw7A1jvm21H0Js2E8nCXtKHriT4JtW7YSLm9+EwOShAoldF
YPpSSxo0PMMhKfL5Ryv36rfep9474ZyAeEjiJWOFdjBhu2oZ4ZVAetlofJqy8bmfwfjkj9Id6oVv
MdiKAhXf4dJswYYSYgvYrFnMLzqH/tB64+raQ9ijEGZCqOaXWNLrsZ1CFX+8JHnKIBB1QuePTyWA
XIZD+zjaNK55bI+z1M9tZOKW2fQxRhs6I1YfebMYb/qJU+v5baq+P2gm04i7WxfOhupz8wMlBJfC
hD73eKuktMqrVVjbKuodERJh/WyXvBKZZLa+2dGPZndSCZX66FOIru+s5etEuEOwQSQNomMNIgJq
WgIm45muxOf1pKDw4dSPbeML9PirKJw0eGEC21SCo9ba38ApvfJacd77NfyzoDQ8QgKlTlPK0LZA
2CWbk9KYudx20JiG0RP7g6cI6DzM6IwoSa+g9TVFJWm9xM5fJsPOPcjnVzxqt96vOyRh/7Zwb6pX
hs9w1iF/8xvOtFPLo9EMsWenZl/Wr2QPLB12hxDZ2Ki18Gu539wiT5k1/3EM4Q4RPFPlE5qKHJW8
kQF4RRw66vr0kWMMyRZbW/02Ms0B4WDnWvSuiqLd4zo8BfLo4tI4d5iVmvRYYWiRj6jfX5Dv8XCC
JMtiOWkw1CmKJD8SG+I/wunhqTb+A5YxiQc5LM3npI3vazTMkpgPxHJ5JwfON1aHV3qPcZ+G6sFB
pCAFFJ+FMneDbZVQXRzFw3l2ABR1MCAvobgxgqPUvkhxyMq0WRmL8AEzO6R1mWDlumN6QlTavduE
DmBS3C6w6rfy61PaSLqUDFvvqKqJ1LouVDHUqtk594BWw8YSdzRHOVjic4SdDXltI4LkpEo896dF
ZFn7l7YDsQ69A1euqOxXvnHF64G16oXGB24r+8PEXuRfsmJsbqtTT+SxGz6HzgxOcFWWu3eOjqKP
ROTr1o2kZxfj0xARsStz5TNsYTi4V+PUcq92hVP/xVJQCCF/aCXAm8GQN+nAs7n4q8vP0KDTXyku
AE0lFOUgrep975segRIO/zzWBxu137Yqfw0nGGWaZ44OE3V6I4EyYo7l/tBxsRV/Bw4Hfh+wjTgC
P+szSabCmE3mVzLI7z8/VUgEwdynCmfCt8RDUCdBWatY/ktQ8qE/H5D80Ff43rUYL/1NBzMG1C9z
LHtXe22IHLlnU9QaH45Iao6evSh8HfgXHD3RXUpCCbXcVjzeHXvWasykgashHwjaAozkABXxw28k
GO4U+KB/FIXHj4Jdg0TOrfjijofGuNRc5ByPj4ige/VmWJF3aQS4vqPjIBUzWXgzvvFsi3BkiSaS
AULdC2eylgIBHu8MyxYfRzMeCyHAyQppOx7CB8tY+guqZhqmRugqf735FuquamcwZikcA2sUOP4m
oE2/0N/YgiTS6hyqIRKz6rJ2lHXrvwKv5ZIN4RrNxC7OV7LVbhds9sucQQYVgOQnt2xbt60rXNTo
wIgL/QkA/vp+UneTZ1FHaTVzIcGbpaKJ6IoAzhGg/0IfUTH+3UMs2bUI6XpJKFWvi/MFAXLmPjBR
ebH0W+SfNbMAQr0aor06Nhc1QHH3ySzn0f4mbJsOBwrjh5+6v7VgJvfTuVKkl6a0U8r28RQeqpZX
WubPil732fm0b4iKgGn54O7QjiiB/mSLGbH7d61KVQO52+t1yl7bhPqydZeOdmNZxNYyIIkdplg3
PLvf+d2wbRLe4hpVD0DHCfKyb47PSl14dTskWYhcUsO2bPvtRJDUD2TBa/3WfGpUKLlWhTdzOqRT
tMV8VEz44fPe2DFsaQLg4d0/9mkzVDQMoCnlLXJAZ+0FD+OytDHWoAb2uy/ee1wqDdWi918WFMLZ
HhJwOruEYjAZLLnnTvylPJV0INfyuQYBd+KqOYpIDvmWmDePJkNIzA2X1zhdqq5nxrsyhwriWNM3
e0MjzpbEpj9cSbxDTzsSdzILeeFTFAJUTWv/96JyvvVz8UeBxpUvn7G09x4gUqCO1o9cUKKIzGHk
cudUutF3623QLX+kP2gkuw+MZdjMljT9tR1rI9tnSY+bIKa6oKfFIm2enTqetHhQkj/MPRLnwnXf
C3ia85ARIa2kbWMOmUjz6fX8TPSjAHGRSNZ9pIt4kxOXbDI1z5JVBQ7vOPtdlTIvxlaZZFAsAj9t
cfZY+SYL4IU3bYp4yZagHS6y1wdsBJYsqH0mlTAqvjQm4mhtvkQfch5Prfq2aEMNKaIBhGdce19y
rErv4BEygUjIN5LM31AdCEVq99jssJiKNpXZfn4Y24JsL/xHr0mjol/Kpmw9ll3vwCnG2dRlFuQf
Ui7D0T17JuUjXfE1l46VfQ15SVYTGh5UqTKTTMOljUDnP/9iTxS0LgDN8sevVEiPmAyC6ivVhORq
hfaavEhZOZQbEyasZSx2insJpGw0TJ5Yr5oDldp1VqnOKxLBO5epRFAVNW+l+MCP7lnCHEf/gqut
pHm7dwduP/7FyYwr+0MQOQBwBLr7ORvpE7Yk/NOzyaE0SZEnJnkRe4QA0dblMNBgOvfBrvEuTNJc
npIPOdQ1NlSinVj3Zq9ziOb6MMqeYUlYxjG9JJ9xynXr6emVeuCwK8iHwGD0yYvEPk8CT3nL9OAv
61IM+Hq0diHiFOcoY8NFmaXI9xaLkdNg9khPb8YcRLY+m55P+AFmnfIful1biBPRTMExn1eUVHq7
kZP5RschvmkHpCEA3gDBbCZzXAL7HCbl8I/jPOkVS3RYOFVEvx6Y6G19PCRDRt0IdJATu4pe9N8j
qMAZ8fs+/8Wkvs/anQFnSwbECxNPUijDMLm2L/X4dz14G7epTcC+jpK6YFh3hbugQUsrRYkj3OOR
2KLkOaopLtQpGIGGsjIVhBgOLDdNOH7x8LYUbxU86gxsHOSTOcCOUHEQYWFuEYyVRZeTIDVUEiLg
rhTRaz34sBSPhMPVOW1lbjr1tGzvT5gJXFBSWMirVIn/r0SkY7jPtcjG7wyLllqBDoM7ZSz3bs0J
KT18YqmzR8KLg24EHGmds71HWMxOcZs3k1S6PnXQyudc/UZEz+AnPGAqsul5h6sYXU07uuTM5uoV
AGQlAJmHMhcs60m2ZLztt0RNoDVi6CjCWzhdPf/9XcU49/5aytR9x0F9WujP2qCTL4vwwKMZTYs6
mnWTiTsL3obIPcA94zTEmQR6Kb43hqJ9Idtj9Mt8hLyX/MDyaF8RRiOP393nRcnVTbUI5AZ+Uacz
RP2Ho/aDJZlSNPl4ssV771dHr6hXaIsy19PiQa3ZVwvmXvivLH6JGjWcvt3o/k5ddYCw36MiF+dO
u5RhIbZS5Dxx02uXED0ZKpobAiClxZpAA7hYeYP4MxZ8Fq5kFJ16uknmj6v955/z6hZfEJKJVqgq
2hryBzHmVqcHwwEXspe/GJL/cNSvYuHLnMydOUsaLenXmeeEWko9T7Pg5Ssk/Tqw2FoZ68L4WGZt
2Zqo3LeuBkY8xt05A3ASi871PLUox60J67KmXioRfVOHswW/1bPsfYipw6gOPEFT5VKoQYg5hg6N
8OK1o8OKyi9AxfeW90i3vVLgoyde73R8FnVhJibVxtsfsUAGq+4LPyx8CDW8b3v2N9tvoD29T0mG
yNnhOq4pfghZSyIcckoiifTPOb+lSNK57G/WJGTyC189Ch1gvfjBcMCYV7W09YGda71BIOH8od38
K4aCmadSUI8/vw9la70iyHCAf0XsqxVHVjWnjbZV2MyMVNKQk+IVbW8KVIAulbFC7LWfE1KnXVP7
gYdHBqRKd7DY6OjEtQAlYVcq8rB9gYrezpoMfYMsRcd9bvf6UWE7cWZn9/+jn6q+iVJ/HmI4fOHv
fGntcgRu1VMMz787KEwLJpEfCY/3c1tf807q4GhDQUmJLY1NlUH8A+CtNI2/lch4gA1zLp+b0WW2
LQncqptDCUMc696f74Yznx7HzXqenU3SodhcKyG4beVkBtvDaxxHjFV303usUBvCotsG0OeSPYXp
nyNu8UYPst5cExlhidf4RB1H/mLFtOg4WeaLZlGupwk26z5pISZn+ako/et4bK3uJqJwUKWmFmw3
5k6ag8Jb4LjjAvV35A+ph6cAKhzwBQ+Y2wK5St6pmLAjK7PV3EuUr2qRSyxy132sRUWYkfY5K1/g
2ClkaS3ho54gxae9XGvyB/e7f3K8UWmCKy+Zd6paDcjWcpovvYz9cYXpgd1v0JDczy9uvhh8yeOE
DVRwp8IsiUu6I6ETmxH+V11wg8Vftec0pckhb3L/dqcZW+bVbuVJSGttVxObdhzY2Pbmpd9+XLC5
NAZLd8rIzAmuZrDubBml3yIjJrRTDOqtfIdWewkgXZDA0M7dPvXs9NX5jH4m7rKxqjA7owmyqVtY
C//r0cnVF0YmfntuKAVPWbuKVC7ahfxjob5ppDWJGMe290L2TcECPfZi2BA/1vz/+WbPOuaoYR2I
lx34HY/v6YH8cuXUFzQicIFaiSXACv6rmsZQl0fRlA0NjUvdXza4n2CPXG/64Zs5Udsc2dQTHXYd
KGPBdJ7AbPlorPiDf35EyJ0xHSP6APGTTv+KM79/y9CFG660rTbTJQ2LXSUt1ul7nq6yQ8GysBKW
cH22Fxs2qvCwbuNAKBUIwBZdH+Zxw/Z4JREqAtWD598Y5OXfm1+QOh8eTVSjzUPUzqvVHs698U9i
vJAUgDYH9leTiolpTTT2uTQk/KMvxEkZ4H+XDoLtXMKwnO6iXetmTy+bX2HlTasmcGWGCh0Sk2Zb
7HkHBq7XX8Q5BcNPOZ22TxTVjX83i+iVtlGsaTLx75tOnrwbYho41kkYxGJW4uQq1gBDs7eaHsMT
qnVXfE+6ahEwPBcOdLtO5IhLH4SmfAXSH6GX6quw6okgTnNJFMjbtnQYxlgnzQjKlK9RDuv6vCq1
YEW+SbIcSwfWEJitCFk2Jq1KmAuvutCMZp2xGbYJgpasYjcdMnUIElUG7f/0/jwwl9FiumfZ1qiG
EFcKagrDsBUOoviiG1rmuXOcphbqIKXxijNe/a0v84hsV3jedTSo9WbEizqJXu14Rzid1+A7a1NC
LmbCpSNU2kUa/9LM/PdbKAm5ESkOthDQdU2fBwCtSdXwjaqJOAoo2q7mFqA9U0AZmRIBiSVyV6Zo
WqmCWjM/YG7Nad7MbjEhO8Ns2GDGSi7DX0DIhxCjfnesPGJasFK2v6ZARX/pRUuE+HqyJParoXn8
tWsOCGHGonA0PmMNT9gL17bwVAUk3M6WnY8SswTFx5iSXDccJaJtimX1eHvGIKvv3yosgNnu1DOg
kuTq9uH1oQOKPMTWtnTVeHMRXnMyd1tJeekZPTHOYvhaboh5MaaTGiwYiyyFMo/VMHFnbz2NklWT
lIWt7LN/l8DoeNnhFVMKBKgnFKWTyAxVgh3xKKI6OEqWGUhAbmkyGzPBg/5WuEdHRKLzzGa4pkkC
uTdvxClwzTxm6Z2HTMVzvrfCcyqknXzMwcgb+PPEDj9ZGrGSTeEMxKC9O08Y5h4K59OkLpAJjTml
i95WgCBQDgp2jPcKVPGFjkgosIrGLuj+BDYNv16MjqipVauYsvWKu6mbX4Z3pJeG2wcHudh4Kx9j
YMcfLhahLRfWmzf3LhpuoYIL8f/k9XsQagz8FUuKXu4oTFTTQnnHLzgaDls+IE8gYRPa0CLY5AIt
quXoVKdKhJvJD2Zq8/DMo8UqyxOG1J0c4McqxCfLDXfADdmp5g/XUe6KQrmQex/kwyuGZF2Jw+eT
DU0EcWjYAHnp2YKO4asOhnJetBw0jNTGl343xMvnW116Skq7tyWjfLPol6S/d985rRFQkk2gFQt1
TqfMDjKNz5U/qrUMk0DGgS3Rd5ftdcFTz4ZiAdc5BYhh2ylWyIEFVcSnKfvv74TT9MvRlyD/dAXb
tesWAUOHQu/5dHKKL7WPgIugNklj3YaMnYIrrD1c4wvXjGKEOikKZSZ+R0sFw502z3Ww8SFHvTL7
9wrHE+D7Zx4QkZQmWHBWdfTDNcb75obGSxAjrHBFcafE+aMKLATcEjRNfO69gX79D+B5BZniv6Ax
NPz2zO2uyYWnYye94VSgseVw6rRr2t9ikvohwi0s3xXCBWYa7xVRccsNLoMRCYyucVjqXaih7c6n
6D2dYVTyfMt9vGG4ySoiD335oCmKwWDDrzmfHPP8HddK5aGjT8sApJ59nul6mBLLi17bOTLDbQ8+
2jW5wsug9y59qbDjhi6Wt43dxCKSpMFonP2s5X/4UHr/TeZeHUfkzpuQUJln+PDoBI1jmJkEXo7G
ofKefN/JGrwfjunN5++v6UcJPz06w9rTev9Iz+9SUSWViiwhfqEc/kPBRX4JT5HJL+xn7hy32j/h
Su7taemvFXXKdiiijvOXPCIqp0Ks1IFss5XpbGRd6Mgcj6pkFWos6BW3o9eUSbnJvJaadcHHzCw8
uAMejauQTLoNBqzd4TmC3C9Fj8JyE+/WLxa+QyXIZQAHJAafpfREPK0azQfl3poCT0AeBGmA+CTK
8/OFSJbCnrIigrLIRiTaO74UlYNlFNBKl5v+lle6gphbgI3HCihd3cxZhNwcyYHe0zhDBP4l7EGW
yCX6nUQUBoXuf48C8Pl133xofeBCZYkso8mH0jAWxHwgcJOqNzEbKONNDVBlyEa9h8Wy+TGj9q9n
RTMda5KkCgppThVG2+5/48Z6zd/Catqlp5wEGHx2RSOlR42f9gYE7y+JSuAaBwJ7WtSjHznjmzOk
zSvYPZPqcbrbj30V2venqVwlFq1u6syvUazagW1nY+wD9EpnAEeowyRR1rEVzpIEeZCnJp0miuHN
R9yGqzH3d2zt0Ww5U4BBT/WE1bi5dB3GG1TdW+/FAD7BHV32IVjQuViSdakFuyP1VxkFu0TvJXN/
Uzjapj+IL5w3mA8FR2G3jrRKxcNHk9Z0RBb6+xzZiKVZm3633HHSZ2F3Gkb2VWpf3cUju42S0RpG
JnmXZvVoeonJvsAqbrJLIikbnRJXZ8jj4ahxaVuMr1h4286OXE0fDZyNhVggbCgJaMZ0HImtDENN
SZAHXN+ifyxYW5ZBraB+5UydF7dMq27ckyZkh8KO6Z+SqLKMyVFOO8pi/Bg/NH8wJa0gLkpWKut2
r2qmfgFJtyYj1H/MK5VARte8q/w0ka3Q4Z9qybMRG1wv1xe7qMKrtUuepjWpeyFv0Mp9SSO3jQTQ
76gY4Ju79gPEguQUSHgCmhWaGH6OYaaAXThLMBe+bpa+ijdKSgvYGaS8fw9gHgvL/AozwhyUTSJY
X9kya+DvNGzHbTNc7pBn55AQPdHJX6W31ZjygT9Z33WkzIYtDNuGhfdGs/bOxs3I+tzFnEUHsgvX
EE+uTwIxIyGr0YwtP8kDPDq5xxQbW1rsoqTQn7AJ4pxurhjM3ODKCpXYNb6MUQLCMlVxzsxj4EQq
OqcZmpOQHWqsgMQMBnMIGOe5Vsu/uFFKfLj89fdKvDSq8oHgR5HqQx/Aml5Dqv4rjCQcmNhtNMwA
pwti9hs8iBVZebWujdtI925xhOsiItwh7rRdgf1GjE9zsmv9ySXVxFlwf6PqrdcDroW6bmSAjikd
g9I44Zl1L2VjaRMKceXAtavfG3LfLzlzIC/XjdMO5s7pTwkVe/amae6vOVNQVJzoMNtkzvKqbcS5
qvkrfVZj4B667YbdIItd1UpOSgQHjIR42rrdv7SE57Iwt7ujmn8jNLwY96gXPAiG5tE43/lomlYF
PXmvm0mQWV2bPmwGT7h9wrKJ39DkRnQ90jmjI13apJkHYabyPi7EWzajvWf7s6mPFMt4hQDD0rL0
Mc+wuciU+fLTW1D2Sz10zrNEhS8U+cRnCLZK/k3/xxfUkvrk4dGim64EgsQ788+735zxa13jzQqk
xRiXusUiH/UNn/TBGsyqAoOuoPL5lhGGnPDLzVQysxcnc/IfAbcN8YpGAzX1Mx+DHJbXnTRohGAB
EoO4eLAV+IhN6U4w8BKdmDNF1k7WNSUzHo/fa6i3xyKehulSxGmXYUDmkGeocR4trNz9+QHm3Ap7
A0dIhzfJWuHA10RfUmeBht5ub/qtUxLeWumlwl7sCOoIXjPNYr/GZcANrTI2//l96vtIw0aa7VQV
2Cy6/7NVRiZpfvooKiNgL6RG5tDK5cHNbdEcSrPePSPUWxSyCZtD+GvWIC3LZ+GwzaPd3g7JDJJh
NGM/CXlp5XZ5SvdXolHaw3SjQ7Qd8L1wZckej/37JAOl6XQtoBZUs3WEnjhCCe4RKHQnuBWlHAN+
q3EDod27AP2CklCyemlXMUa37QhfMHLCYE72O/UUNIuWPrbSCOJ1/dmjXakShEVeQh2QQ6xa5ngP
lENpMA4sZlwJo8YEDX6sDlcuikczNsX0VY8mL6nwyVwtsihzgc1Th6a92vF7JvyP+oOLMTs3U1GW
HNif1XEpWPF5pjkyjw4zFJzlgFU6MPse2xjYz12lXd5nNL7pfVfJpxDOVglRMNX8Ap7Cj+MnJ4uM
UonraWCq8sKbTCCydpPIX6n8CYEY2RNJ7ZOciDRk4W2aaJJcpukbTurNl7dIBOhWhNEo1zqdv6Y3
WC4zXQG2qnlARgEWkN5ggUv6+5XvcnDnNgAFnTMuJ/FXjtB/5xRl1eVq03nzXeAqm5JltSk0iQgn
an4njFDtkDFl84rv3rPORiaxtHvv7RTMA7ypG40xt/r4fblWqGBaa9MRQz0uyQUaXKp98t8S3DSq
IXMHcAQfiGlUxvII/tTOPl/Px9CT5/nwQIV6sfz1dGfnS+KOS7aO4XX/yTQYRFDkLC15+Ldzw5cq
n17UKjfBCkdh1deTMdXCTwRzjgB0ZxibZZ4iv7pgA47qG+o8Kztr/5SlCjoVZBaNYAELIftoGBZi
4I+7QYq/Mznjo+C6UXLB3FWV+W1unWnuzfn+W8gZ9dP/anH7mOxKpm8WWemhq8GPCx8j9rnkoWRZ
pt33NszqWG4sxRuow4P5dAmhAT7HXxIe39UPrjxWo9vUBpAYVfP9WnElGvnD/zDOmKXk46ZGeKuv
j5jSI0cJc5Yb8M113onpw0aTt/XXVtRz72+ns+5NytoaNVUWQOv0Mbu6+BmMWMkH+5+HypePeu2v
UHuRPobx8OUxm9S9J1AULKdRdiyZ79R6mLzKiVSJZ5tX/7m5NfI5+DF5OTRYb8f69R453g9dsQ5L
eGHTvOSj3tSH20aJNieBlmdRMi5tFFnH5mF9rk0HwX9dRJDL0foYfB2/dw+FsaX+t0/udVASmAtU
/rnGuuj26wSlheXzNSwzyEENMlKppeJdPcCR5/hlsbQr2G6tlNcdJpv7MewmLR7mZjfHVztXLwNZ
5yr0qDJDjEiiQrTSMC7Y2bSKrH9hfosR+cB3tT0fhZQbdsmxmy4HUAZxIWaCgX5k6+cBWTrjSOuW
arJQVmbhiacqtSVE5EoleToSY+x0pqnmsrnbEHjYQB7wtU2SOQ1KE1bxNnRXRRuTfseJutoAPzd6
bOkOZXm0pFgyXq7qljOc2gux8Tqr2jJhXeINOLcdbeVGK3inVJZCFGNXO8sjGr3DQJmUdokd22CH
0AZdgI9wJcsDbpXgtPttIM+orlY/3JaU/6tVRrBdQb80B61xLROeIDeeb47q3rJVbsfg21wwDwIx
tj6lxgrxunVXG6i9O18Eam0Ng0oCTXUilsxNzJMuYvE0XfnrAigiN44a8Kz7FL8Hiys93AkrZmUQ
Hyv7ZmIfH9qZSd1n1977R/BFG7v54JG/NjP9zDhXjERip0buhDgoQakA9SnNohwNeEKk7krTIE5L
WGUjg91edzmnLAbZr9NcgsQwPQP2RTkSRdY5Yek65m0t3gFGP8vjD8YgCk0bfRzq4OjvAfMwn9I4
iM+GbshvpXVF7L7+/AmqlaMKOXvzNdLYpSdnigcLw54z6hgpF6f7wgLS8QddiKYUp65BUQjAa5yU
U69Zdhv0iZ1r7szZLPIeU0NP/tfXeQ6qehuHgD+8poJFCyI0l/ocM9LfHg4Uh0zogO2HuYryDw+6
ab/Amj/KDLTF4WJH1QeQEB9iyOMtrZwNXh62FjYW0rGcMoJ6WFJbr4Hm3QObrNyrFG27tvSgikfg
cO1tobwDs5XC6LgL5FGGpJMKQALbU9waNADQtIP+ITNmA+Ob1E7RQ39GMpK03vVtFknZerxcfWdQ
qp5uODtCKmb3fOAisSMNQy0GJqDPl3CRzGYIXyqSpwC27q9mh2vXO0WqMhTbgEEqemo1DDkYfgjk
b+3kIVdY9UO0P4qk2+9Y4q73Sz8Rbi4iORwpiaX00LQ1xyC0EeypJB7YGvpZ6Ye6CxhcmHvCn8ka
RwhbkF1J10/ZzbsHe36iZY4disLLvuz329drmkFw907ArSLpbtprTNZbgM28n262IirbGGj9HK03
vqzsLIwrnqHVNkPD+xDxmxrdBBpef+E9QfQz1kF2FQZbUsmnWIu7+n4m8MqSwH3G9UaiAzLrwcuE
FixNR5P7Yyl7jteg3BO2/ChOO+QfPV7o0O1pzWfb6VGWK99M2wXeFkeE3ZvlBT3HuyNIkJnW6y8t
1AgTYerT/BlqHjfJN7DS9KLGCi/ixRxLg3KLtPBqt0IRe2Zz9aGrRY23DIHFhZet62N7Gxmo3FW+
JBWbcZgziC0SrxqDgxsKiTaVw/2wfaumiE06s+wr1NDvtSYe8u0fjnrbic+iwOJJ50JoglnNJf6l
X8gTpTG+5y3pEHjghBepktDQE5eaaDoYqPCfXcn/5iqDY+HX53aJn2cFvrGx6+WFix9hhJ+uK3d2
a9QKD+koydd7D8Ts9z0aTSRqSXFZP5YeLAkwoTAjWOW3I7kf0z5rOTsK88gwEeqlba4hFwV9/cYL
b6f+LbDfKXnEbsYImTuoBqNUCl4X5/sEVgJd3bmmGqr6bt8vryS7xSygG3ZKPtNIcvMLh55Bz9ji
aQ9aZRlGR/yrgO7qXIoZK8LJNLdaaVXr0chmuq8gmBBbr9B/9EggQfS3zVJAZIlhR6FiXPCgPR5A
7Kl7NBv0jaDpGZ+wU68NEpKU4BrQ6eRwIg+Ee5rkelcM8DNfwIT7bpsYnVqC/3zwYYzHuQggrmkp
jB4JitBfvhmkeeGFta6ov2dU/chEdx7bYrgGXGNFyvS0l5AFCKGAHotcDaY0NJk1gI4eB1vCHfMy
KGgdfnW/AyJzRIG1QR1GabCzF0Ga6uzhf+8uxSgGsKk0rMD+UsqCfUdg7YsxcpCG5Xch6KsnghGZ
twn0k6kaDT6LfPHimWmUxg20hIL4YlY7gKaaD59EhYNO5FHCpemB75pwj0NPJx+walwf8xyD0vg1
TL7TgW8XFYbia27Aa8a40PDFnOG0Dn8hO69EL6w2eJDbRD5aeej0kDsB/n+k/hbpvEryte73n6oN
AggUUOli/xybhORZItRh3zl+AlUlA8bHmUXaA6TFhZoh37iohRR/xtEHfewhYWFnLqTB4eXchl0F
8JRQINHw4oaawOm8ZW3Jt+IXX3kIBhzoajE0JN2MVTGbB7PWUWmMZGAbR0tk25uIo9fN+ddhRYxv
O3bNSgDcByetmf0e8iss33ctNdIsJxgHeFXXC6i6TGR468MjQmtkqc7aGBrE/t52Xs8vf3X1IOTb
hXrV7h/N77qmL0lNbBY9AfSyBKV1v+ZUwzgzJ7dZIZZoHYvvVAwBGZQpm3mqdbYtcKQZD+4vFeBq
7Hd+p98i9vP//xVUeh8p+HVMtQnYk6ziEDVgJSKegzp/cHpS506MmKZT2I1G0daFVfc+TpMHjSe0
t5i4znAblvWnp4IjvFxMiPo3UASRs9Nnq3rRi+kimY0WNvorD7RMNDtIrg8waYcGDqVoCeEgumyv
gaiHOnfkMBbDKjuMchLtvAma44R/eXVvSNk1dDeYQG2kk0Q7drrhe6ccRRiipPRKdblNfRBBiOhE
ByApww7cNXNDeQ9GptLph5WfJ5qJeYN/LCjpZ+xulTogkhZex7k182kENXy5FfU/rr7JrjygWw4N
G6nFLvxaR2Dkk9Sr5RJ5YHiPRd3YmaBWKxhF3/SQjXSgSkS5yeYktgIlrJ44GSK+LWgR0QFimMhy
4seMTWsye7Dja+jZurnUxzASLBTdW9Ra03qveGIYULHYREpPVvZQeYTEYDlFx4GIHetZj8DneXpV
ZGm1AnHd3kL5kxEFA3Ry9m2Q7M3OXlFHuCHsLdY721//GNX+zBvLY2Sa49QKwF+Jk6NDo1r+S0WP
51skMid/WeBGNrIZG1tHt9HzmNmynYdhcC3xrJ4gF5KQrdDSUhyWKM+Q/shEDC3Zz6Y4Od+JYuGg
GugQjg8cpVMFnZ4jbLAIaSBIXvuYK8CrigiMZsF3YNCn1+DBWCEgFc4okTrUIKXjIG8d+7kui8vb
s0KdgX90fHjeItBV+EcmvShVdLxHuySCgUz2Yd75oy+Bbmute0nj8pk4RQG0WCB9qhCN/n433nwL
Fxw2inXiFdJ7XqCkV6OxBMbnOIV+W8CKeE0EfUxf2RGwIiDuhQUsB+o5QKyru17Ouj+ottpQ08C5
lq0g49KBBMFfNwUm3j5MfDc/AORqekbocDbRamQLLZU8eASWbbhGzTp6e9baV6X79Nu86iwBkVRO
P2ckgW24GCvpK5B0swBgorHPL2A3KRAIldGOMwTGvwm1LYfK8x8i3+C7tbcZD+7ILPxV5Sd/2akw
6ci+catc99yPbOIMSa5wxsPp2Hh2EJWbv9YtDXum0H4oHvIgqRpAv5BcsdpQ2zYjUX+A58Gps9KT
HAQFLckGElc99KKl51Kif+O1UQYJX6RGL3s70wGqCVA+kXSTM6OmHIqvxsp1MCH8/OeaKugT5Cib
f1BADEBx/cCy9MFnTLn1XyMii2Oeuf3pGfozHEGWTFWRMpaKWlM/m5ZBr5yEPyRHoDGSdb65R0Xw
ebNUL5VUI1bVhTNLaI2x5Ml7pOeapOzVIbxh80yRp4rh0W/EJdpvMpBJtOgbB0XlcTra1FEiBNpU
HdyQ9mwYsBx7WUegdxE3WlEB/92VfcLrBOkFTXwMfCq4SdiWbJkjsrjbDLuXU9fwvJBM8UQvqGbg
KRGCMOhLLVjOrvlSx/w95NOWkMwc5DRQMlciAQekkANnn53kcMeWCuQpBxR3WoICtVJuCCRnhKWn
gS/ltkDEMZhOMu/iS/klNeg7PhGA1/Ry65bMbFe63Ln3PH4ree2PM6LoyxCfNmKJ5AJxovq9R8jb
zp0EDlTHv9ynC2CYUO3bQENBSb/UYWTm6pLDGbFYHwnu1HCpx8Is1c1xVq5jKSX1Vf7i56ZZuOhs
voWD3xny9UqNf83V2miqBRuQkgl+aAJJsEt6LiIdbolI5PSwNlO8Q5OGFat6FHSRpsSPGWNJbxr5
rNG71yavmgWFzLCbEDYRvFwXm/TwuH1C/wYx3LlTbLE1FSjtEeBi73XBB7iY6sEeq1NnvSlsvaCZ
RtU1gaGj9lwLzc1MV2QEPRog90FcxhM/HZCvmWqwg7XVxOSEVCx0lp5I7Nf/+Ah3T8IkMzW9jAJF
HKG0NmWggDjbV0DHDSSbicqryh2FPS+TpInT/Zjmv9ofSGWnFwZKYqWEhgyxD9cxhigZTOshxmjx
IuwTZhSB1LYR6fI07mr1MT+ETUcOXPFUN16eXdI36rGQ6E4NntjAi17u0LdwBGrQGOc3K/o6cPB5
8WNOlZKK9q09y2hZNCmknN+wmo5pu7vvzD0ra3YOkmdWhXXMhfNB3PvqYuw02Vm6MNyzNA1WVReO
gxapxFVIHN0xF04XNv+Wqh9CUrjoZOy6dh1Bp1CzsEAl573zASpCexOaW0Wbfha5H9Be+8z8/3PK
fZPTl8Yh0BpFjfNXlZ97lQUJ8oPUu6+fiM17YrefK703638E12wjT8jL/IyS5sasy5HxPVZd5C7q
Z1PIVTPLY2KKXkDSwUek7w5DOj86UCoKCHkqyGe5GATb0bbZYSFyfSaF2yxFtOiMExprdx6liEtt
WJm83Lox8+KgA7Oz/hFR2nBFjgMRO8HBSXb7Cy1m5nt4QESEE2H6LKlc2bTCrakF8ZeJEbjYw7uK
nzX9SBrnW35HjA6HX/ggDT0n86tYc6EKJd+sHjtF1oEzPw61jHk9sp+cvUXT9cSotHwIhJ0kzxFs
7wUWDu4EvEDusLGXTt+h24vHYlqiX00ck/XlWtNjbi5ieseLdC58tZ7KS/TWuSCZdOj0PedSsH1S
78qoF7IybbO37DtvqWhH+2RISYLnsgDiT+EyaZcQBbjCfvIy/61AJhQUYfcYCb8TTaKHh8Z4oJAp
qIwRMGrE+hPi1KaMBEcDgyv9ojGRewsJgd4a6KnhAXMW5o3g0uKlzYy7g06WO0Xb//lYVju4W51S
An248lRkNd5jBBZ+qFgkOKidGseZU2NlrsECwf6kjT1UZJx7OvQw6Ftbyh43ACaSwk6y9Yag1JM5
PT96OVNQrT1iBVy/Rj8mpSu29uYqcaq9FNwne/Xvcd80MMl0DyvwxT8mdncKTnTa337b4NHTsZ42
vt340UpFcbL48x3zvmIQU6WYSfGTmFY7Qf6QFIp1Wr0u67c1Aevkf6/DtdKUncIVklEZl2YxmNcz
xbEQr/MIe8tir7O8Eo5GhECC1OhlaWUtHE0jUQyzsOs8svH4HggrN1B6n2qyfXn7N90JXviyW1+p
Bn+Z8RdotjoVsm/a8Ha90Fyz1OGAiycS2SiGCu4J9Gax3sV/Vjsb3h1qtsEWHThbbOqaLMBohB9a
uKA3bOFtb4bjfspKTWxQBVenDU0eYzFEcfl/KkhKh4pYZe8pgMqPt55J66w/z1ME5g3gzIMepVXn
LbwNv14ruXh96tIXj5JHD1NI8KNI59IZBKgA19HLxyV5jxtjaM2kZopcHp30L/9ts52FWs8u2esr
XPEzaSlCrzCoUoL3hdlL3K3vMRJeXYL140ofbU/np3UiMezb4j/LO5L+0JDFII/R1SOOi1m0uxE3
qKmrwr/AFUoftAIIUMb6YoDB2VkRRUKVIGYngKmDNpFQGd/tnROKmM29Uybuvj20R0joyQVfJg0U
UzhfTRAzGqp1v7HsaPrXDpJgLhfMo+krsIks2TsO5M1/8puoqirukgpnjuz2sPo7tji85QAQzaPN
G3EpmPqyrh6XrIwFV9//gOLJjjzLVrXlcd2GNQhz2m5VtncKbCufdCO/+aFumHUYFebNCvWhdO5X
/VIDoGY5vg2DDBGKYo3PWqqAtJDr5ViAn6feP39+RW5YjembplkgYlQyKZ+oP3sEvkQf3lcrXRhW
UvRGWgOnxV6bbVLsElJXB1gW8V9RhA2FVAjLVb5s2et3Jlu0wXwWyrCwKDWo9glmGenyZBnTaeWo
wjhqkgzl/KkSrK14ug/lNIoXgcA5ga+PgAHszuujSSyhJYbAHAOVTKxgxj/SLy38ze3VB5ZAEiVo
Zu5T/KbI47ibRCjiJ6sjPxGuMnJAJOcHV44+du/FuF2wOSwxnVRIyT7GiSNrLwl9aOnldZ72Zp0r
F+uyudWGoWMtxJYUZGEKDUDWTbgcKdy711hy38MrdQJbA6oMFF6VvTtE4CN53TImDenDFQMK8E40
t4tcXpBRFEtMJYH9u7jfSNKPZEKEeRHiR2fzZKpWEB+SEI9VGLojfYUyi6AOMeFoe+bve6uUMUEm
hofSlil73qROsAB6OHS4x+Zf6JFMoM/AJpNfl7MaD84Ni3Yv7SKPn21w57MOm1dADerDZ/P5GMQR
rDT7Y9zWBmHV32rNf28BW9G1X2l73jpJmt4z+u7xNEYeF4NU00uyNPT4zy1OqGeRXVFozlWXE7FR
ctV0ejXYWyWCxKoH1ogUoEdyl3B1TGmjoisrY5md3IXGTMM7e41Nd6m/TeUuk4u55hEEhyDDAj6a
JwPAUbltIAlqFeXD3/BeAQwhAoy3Khc9ArqykxG/+a9qyoojGla9wyLFSd1p7N5dy1csmL8FBrKz
r4QIdQldw9BXAlfwKXWDFImtjyWafmsAWjU1nk4fiHGKPoLVUqXbMEBrzHUHpm/ejD6qFFzlHCa5
kBYX4QjaNad33QUpF3/6T9eK40iZ1pAWgV74XwU5J2+v8LYbR0tOTd6jIlFkXKPsMQAuDVKV5b1S
nRIkkcJHCbJT+nXW8d2kFJM/q6tmLJsz5DG9fPCiKc3vjXlW/E3V972E74aXwLpf6txgsJiMjLo3
4PRGwjMGaF5ShtxMHGgORyW4Co8thJHut+r3iRj77iTHcBrmR2+CDrt5ofRouBBbh/qLj2/mJO4C
LYGMM5hR2pBW5UxshNtK3hTfs1To3SKFxdIDLquwFc/3FYK/mr+Byw4zV9RJip2DlLQ4HmXbZLbz
+0HrQeWWz1QYJxCPL+sPTfHw+ZazmBPowRliZaqZt5NilV7BSWSUufNLaGFiXcwKv1uT/8zMPjaJ
KmFExQTVKUlva6ejJWvYBap2xf9G+2BXInW6Iv3Rb3HaT66USY9D4Q1z+AbCUhHAMgH4d40sTT2p
GNpVyw1DEk+db/qDpQJM0x2MV9XZ1b+ooGqEXLQ8fJJMYl+tjjNBpvKzWrcozRP4z1VhFCWbhW8y
PGIYwIwPYJXayw09pDg35K8xFBjN3qrO+zbiiMwkhGGrdLfaFOQefnkpJuueKmLqEUIPks7J0NSt
22RGjSvzBCRiMaaEYlGsi7TPx/SIm5CkIHaaRHAkVMea0QHHdOLcREWfPvc6iinxQFBq/WTtpdvh
bf7UY2PfQRS9Y8dFeAP6ZARdzdQFAGfNVq5Bnfdigb3HW5t0b06ZuzhxmfBcvIp1dBjFHi43ueOG
Jmjf5VEPFhpX+dCznehJpsMLpN9zbN1YtMwEpZel9VUXqMS3qqgyngvYWBSeRZDGXxu4lAJcXyD3
J5zKR+wut/kRNgG5FXXXWrLVlfuPJ/sjwhE0X23ogCon9AqHOHGzQAi+LyNB0Z8/5AEfALH8/kVs
BjrzWrS19ZTRRe3VT4TPeVtds1oy+VwAg4dIv4LeDT66M6i6XHuW4luBjEOCj5b2NBBb2Bt7WyT6
OTxyKdk1+UdJ9pGu5E8AKuoKLPUusDyAizW3tE4GSnE2Rdk3AUSLupiCnuXhEnnOtdgLIioUgNnB
nRNce7505p1ft4n1GrPfN/WS8Jbaj8BQOl6dn9cnxA7Zm5YMmLx7AMknrZQI8QAqrPqQcLQWEtl+
p8ZHm8tbUTjAsNzb2oiTTr5oNyY33mYUr/BBMZsN+2Cdp5m1o4Qrz1G3ye/BNvF8edE5rLMATuaM
RKcy1V6OOtEAuzNy3DKcQ4ONyhkMUM2ELgkCM+uK7hbS/iAnbt89BwCwpoPuIqSFzPbCIofU0BRQ
P3JxfTSqbleGOHZ5jGA0LikDy6QMZan3mRZQxIbgyRhsTjikK6fJlmcTjRc46mESzaUafVuPsutb
4G5O+A+i1XUfB1zO8qFUG6WnmJ/7bSwmk0o0qIDphOfDuFXpzmPIXjptQOUOgTY6nSmGHpCpcD7M
+h3oGnGOlOFsnyyTS4sg5nXncOLGflJ92V15A60H/GmFzAjWeZ56/IwOD2OTZzbcynBfrcmbAyIX
mgYMiyqPeyL1RMzNiO0daXLYHMI4eMuiP4qN4LH9q86Wpuw05QUnY1ZB5jRp/1GDCImnFhswNHPA
DntBdhDNsyHuBupJ7gf/WppVBL8wlDkX6t3IkaKgBqacGa/NI01ZeafAA3jkgH7G1I2lzFVNQRVw
J8Q7Oshk5+g93mfJIMZrVe9/j22faH/o2Cp8xqgEfsYUt5To51trItmfkztw2q69DT9XaBv/mBee
r5td2xBCDS7Ab9jZ388yLk6jL9C5p9M3sYSyIUrXJC7r0PKVmgwyKfNavo6CnsvksOLVSrbBvF0h
1AOBZrRc7LWRx/FXWfVIoJ80Hkboy8J4RjMNF4BN9EmdAoxUEJccdBYBKsQSO9WeUE4OIKcSKx6S
UXTR6IF930CaSfYOczV1LAsvUJ2JUpeQVbdg0IjUgnmtq3FpGlFzuV3SUS3KOq9Cgv77PytqNXeX
LD+7OFeEA42TMODqpOnoJi3cXgHEYN9hfQhFOjK52hnytJ6twiuOk54p9DOCV9S6yCTaOUjUE14o
Rwdlnyc5OCo2f51IZ67rRdLIHRSBcQvZTu6fBttDHI8OH52blS7bj+Nqk3qmZNWhO6Xg3PzPogKq
5XEXItrxL05hfWNVpH3ik5QRZVycAsfbv9x/dRf0+Nd0yANOhilrVRsoymwqVDq47G0xTCtc+2KO
8Qp509q1Q2qG5G8yA2SH0/efLhjfeWezCkHCq4TXfq3thyqAV/s3sHnZ+4UfORWkM+5AqgPL7vW9
KOGUDkQQX+VCgXj2q6y3pHRQczjjHMhvkFl5sBCLBN3IDfyNtPlEA8Ly2ZNY7G1pGjkBkUOjwUxo
PJaFSUkLkKZQfKeF8tC7q5x9eQ2TFew/chpBJQIndWXmBg81TjnLjeYfR+ZOFC19vdsLuSIXhXUZ
PKS6bdiBkTunmsKwqsef9AIkY1NAuL8K8yWL02CcdH24NoRJSFW2DQXKJBIR0H9WtAZkhhZf9AF4
O9il6fiayA2VX60hXl1RcdkszV39IEmYJzqNkzwQkfmI0HcYxhKmuVPSNufOuf0AxEGv0+UkMHp4
lYYTrmDfd+8LvuvMusFaWjkbgoQVoFZVmX+gA5UcliSKDh3u4IpjBTTTGt8qD3922X4tc/PFEFk/
1lQu0Jt8l4EERPVPBN24aTlqlsON0nXGkaXhtxOponvwmbp3wn5Rz6nhPsQgS/6xAI8Gn4rspBNV
dfi5wr6chW2Y1JJqfv+JVEoXzYMWTAiC8OWI77TCsNhD/S5ZAReLlesIQt6T05tOcjnXav4RbCfp
PrIlEOK4nCCB4RTsmismVvvnYalBxs0YFZa5ToKA/n2lsVRPk7Fuo/49qVSQx7W3Z2vUqcPgH8H6
USaPpBG4vJNNNzDvNo7dGt7HBM9GFM6gilONC0bIT7oFnPC9MQ3GrFMsXn27maZKBJwI4Udc8cKZ
8HRivYkZkhtfWcATFb+3ldz20OC/gqDBdhjSODXXtf5cV8azQQT0a+2gv5YHUPfjkBuuVZkYmeyx
ga0s2yn3gcqPA5f/oga3L7CpIu7RFKfIFflQC5AesbF+8hUQPH7h9Y7LxooQSXHw3bbX6TfZAexw
0Cn/gfhsZ3c+hf1OWkpT25VYuFTNAwGkHcprIZpw1HWqEjxWE1M2mSZ9lTkHwrGKYgtfaoLUkwp9
FEzss8UWdp5xwH8OKmIsD4ldNEJ17VNU7eqfSn4k0U+sIAaSY0IIkevk7dnAqQYy3gtcpCR2XkfR
hbDb841o9M7I4nuLCzeP9pFsG20UAwgFx1ip2jQv2skAAZPM5MGLUIHehURn7oGyQdzb5mDJQnrU
uSC7onuNCp7Momto5SgAwvG9kKlc99jkU3ZS6WnwCyb//ERIzPG4JnkOyCnoOABq4EBalzLve1Xs
AXpPv6Of7oqz+cpDIp1HVrmURurPp4bPz9ukbvlFxStZHb4tKCVMDDIJB/1QBNXSu7weshtjaBv6
Oxuet88sHinub3TmyVnS4s1M69nLbIHo0Ybl7hHZhYrKspsj19JtJr/zClO5CksqGElDgPypDX6W
ip84tIp6eqenHQIupk55kosznxxOB5JYBF/olFIleOEUTLJ9650uRv4NuFZ1GiJok5LwqO/cUKvD
yzI+YwNP+FUXVSQcrUz7zcMIk8FLx2YExSrN2hYkKx7Jkl+DJMe/HwWdbkejI7NbyWtggMldocjI
H2qe8DrRi+KaD2hV5/LdBQ6SsQtaU3psL/UIe45w/Jqw88weSxEqn32CDKyKdHlOVEPf98HaAJ5I
wX7CQKtBDlJuXNTM/kHwoYTf7UbzV9P846h6ZwHaUW+y+VDggSuExx/5355ehCrsxA0yPMPAKIVE
LYSHaQ+xGjl+9WZnzYjXCZh3Al1x0n3qzKIpApuG58zLtH83mkL3tYm9/xFQ7SP+lnmMECLaVKPp
ZriYog1iX8IBf7VocW98kvgr0ifZzj6NHPXY155y1zqykc+9qPTfd6rEQQzWQ+GXAiQf9d9Utakj
J5oQjMGmC5dBNJcB3CWIGjR26PeuHS2tXdXGVYBUTRkZ+0NFgwxJ3dB6fovGMfnAo4v9bT3UR/39
DetcswD1CIofYkHKkeX4Gx3GbVFzoir/MLkazxlLGlCuhw+x6IrI6N/5dzDtAYNjl4hwPkzZ+ySM
MkrZw4qPsLPiIhLO0DpK9ZyBIKfMfM3lrRiDn9Q8hZC9H0siLCZ2lHwcSRpuzq+kiH6D4ZhsAW0R
j3nZ6w5rHFN9Tjz704sbWh5twjg5UUXg4ep8gPOg7fCNEw9gIU+j1s3pUnTbGD77oZxazU3YD9cL
zVQtQodqL+v8W9NSt6Oo6B0Y0kIm9564wsB+LNGlVuPKPh+AxY/SQFM8+O0OxrKTaNWrG6NBRqHG
tp4LwdiK3KTmgoKvrc6VNgDYtQn+OC2lR+1XPsKITQVGkrpruHCS+ScRZx9GSCjwToA9SbH+iKEJ
3A5/PH8JMe05pkVZ5Jk0FR194nS0bjHwYeKRRB51ZAB8LYuaj/i2vKsnr5audTAkOmdtt2MBy1Ug
fPFnshcWK0AetoCu+L1cgTXhHnWCxZHhaG0ikcotGZ7/XfTiwIEB0lkjKlHfbfngs0LVrvW469Bv
LwgFEsndaP+F7dY6P8qpHNMpT7188n0KtbU9NJkldxvGhoWn1/MjtOxtFS//INx7dax37WJUrW+m
EYvKlJFHTBoDmFi5bP8lVoJKWQx/TbaVgsApWlF24M2EULdu7wXPzzRJF3PsrF50K8v1ZLUgcwlE
S1/E1gDOoyOMuiW8+ueQC340epdB2fmmNEon5qs4mQZ2FDWmfTWTvSI8DYJDRNrC0zS5sf6mznHW
Ti/xxiBQ/w2jn8CYCYQvT35FzwB2Zued4SicK7BoxsPAXzxCXFFzjgjUpzSA3cx9+x3EozVIlYXz
Wctn1wZmU5GdXPucTJd0b0P9CtoPR08Il/3HNdhqi6+1DCsIxVbTKdmbBSnt//syWm/dyqzg2lNi
Ju7QWY0e6rVkvlBzCrky1XI8iHVPLd1QPg6nbs7fL+nZRCb7+d5rVsHyyceS8NZjTW2Wcvf6nYQB
dBBCo5/qJg9Wp553pMiJkNvDujhNfzactRR7cB3U6Zs9En2eLvM7AsQLTTo9oSRFkEKWpSVBd2NN
jvlwMKJRN73ijHZAwSPUpGQmwtSGv/+V5nyYwBOQap5HhDAHqjzibhKtGo11bqBV+BvgzngTlQ/T
uzVnDkJyK+hXmF393kTeHQ31DHpV58AJYgzi4ppYc+FdvPhKPCveAHyZEMyVrF9+PujR1BDXw0/P
GpVQ+wzDUsnv5BLGVEsWcUgMAuOm38TY7sELciW4x7WRwYJClERkqqKGPC/ctuc6ZA2UlckyJQX4
Ua7Gsgl6FuxbbZ6krS7WhCVPjacaViQ3hvZvdci16TC3SIp4fo49OdYwIk4Tz8vIsyddBRssZXrD
srsTbwWjkzr91miCoL3p4Hi6lHmH5glMu3yZBPq7PxCnBXRgGElhFTVpE+t31WF+U+Mt2i/mg+rk
28iIc/z4jr4M6aEzVBoIwTE2eniRIQxOpHV7p3DBdM2Z55mG/Pyvgyuv/ujh9sDsHZ+rPcsUuFJS
hB4YXpAQPUGG22S5AOF5x/JYt+hGH3+YMnIH+Lx/WdgrcmYjA6RiHWBaodVGOLIvfAF1DKLv2jPs
+t3QnO04vpV0tQ/FeIJxcUD2ECywnXjo5ocRngJw6r4bOQoe/8Chub8S3KwzfItUyebjvq5OA4wO
2oS5r+EaOe4EIXZgnf9NkZ0ZwzZKzVwwr0bAEoFPmC3Fs7AnGeJMmn+w7uY2CFZ03ow/AFMODWIk
PO0iT1V0mgzCSGCpwiqLu5RQgR8Xp/IJvg+G/HOo53wdZkFjkXcMwGTfTkk+lgKVGNM/SqAkbGRh
J4OnmN/5r2U9nhOCeerCHYdPHMlecoMu1A57slOgpp6PTyPPYkkbBEhbVXlzg9XZSN4aHjZ4bmir
RY1L3tcwkICBanbtnYJmUeNsQ2vLxFPmqxpzwQqK93YKuef85XwmQaYJjhn1KtIpBltyK+6dyqmt
VjmP7+kxAWR+0BYH7rZ/52PnQTLLwW/ROl7jiU1FXFB4sHjaK3Jr6aHgfmuOjtpBXhmfYpU3nFFr
AWBRm87GYSDr4u+j9jV0Ukdz27FoUsdn4GZa3Oxdh1wUuZwuqVTTwt+cotqix3nYPvuoX6hv6PTG
wl7Lke/mKCjFof/2B7R4oQEGFcGTC4vyVUWDvoGj74UtlbAdE3Trdy6o6N0TUqGXSXtYOS/t2CAb
4SZtl5VOJ1eayOGWpYE/2aNIayR8MR9SM/LJOmJjnCsgL5tDDu5oCDNni5PSWPdaf2hCjWXkacUi
hToQYEFYt89BgWBpufcFTi0EYgqAqu3LlMvWGUNeUUmoh9Pu0cYozwOvQ8v2FMo20JvefB3AQtOn
KrkwTqzp/gJihr2CaoMG1yWWEbZ5ea1U+pWt34lVRaWsTebC+ddJ8PP8AMzacLn/8p3OkUDj1Ufw
5oanWtkuZfZi898gQA3cqa7fCMWMrz9oGBqwrE/z9LjjZj9zHx+x31YvwcFwE2O57wW8P3uMO20G
t6xwpSrZayig4ojsnoD/eJrLbK1XbjX5U118099WONYjtfzN0pH+PctFg/sg2YMxjaHXo1+KQBeg
jcjKMVzxFhCcd0kgnAjO7ZKHcFUXkqYd2IbDmQj7+nkayqBuHCK7cHlPhn4sCY6A4CYs+xRuuit9
ijRYCPnJczlSN/1hR05+4XgcmER52t5NOFZa/z1NqFlrfUQac+Lnz2jNOippPrWEe9/uo8lt85+I
WUYLT1xDsvsK5qb0rIylEl85JENoZ/TkA0QirJiTPzSpCyXmZVqmJL2fwEizky0yvbMg9N+M6MYK
CDe9fSD2KBmlj2qv65IhymU5MlI3u0u4+8ySfzfA0smhyKLC7tFs/2wI4BPg2Z7kAU74rxRaRGJB
EuPrDedDKHRO8aZ2clzvyuJlXMSxYb6WP0zckYFzTe41QjelF759cJ5b5VOEoqHEm/Shw/JR9wJk
x0987rtHML8Km9PLVRUCyN2VnXSXUJYDAfBw0F5xhIlp0+hD/5DiARWI5NOiFHGJUVY36yywvuIK
WMiX2qPH1Iz22x97Icy0wvkSBv6KGFP10fG8fLOLgZcyT8LeWgldY+V56krcN51Kztg4fuuQoQ+v
zhSlOeuVVsp8/PGn4NSuxJq2Bn0pHPj7YA2f9KDE3a5Inu4CtzLuC9KPywE50FbhrPkwFWVZVv6I
Cso2i277sMu4Kba/3ILZ7tgTF4WkoOCnE1VUYqnZohUV4Wd/ziwKRbIyM/A/Bsbrw7Mpx7D3F8BK
eygeUDpISElF7OYNiIX6VOlat42/F0zqXRJjEGnkm6jgdNR3TNgEs7XGUgYsNaa2OSEDHFQSRvnM
s+PsiNcPGFzeoUAS7vXwvSdcqU71M/DXwzdgXpzjL8vnVm8vv6YpiotewYeJJ7Q4ZIpT+6a7vkva
nESXjFJb4uog+SRsdbVVja96xG/6LqFP5Gb9cEPg/yDSwsxJffBOl6ydldHKfgJqpZBicE7Ms66T
FE7wQc+qbQ++aZo9Ka8MJB9O9fJLG/eAc3gTAHY4m4FB6wVOKZQo2F84Ek1qVdq+fD/pBMgxRKjf
6qcrGDIRqvvETfGRwhXdKRTGW4tONKTLmSovX8QceiPEjZg7q73BwOUn/cqGcsVJiXUPBdpcwrIt
dwn3bt2Av7W33jpvvrZU4kvf/QByyovLJVcgWJLHeBz6iupih5yW097Ev3IF1taRuGJfoE1iw0eW
OyTQ/TTZExxXopcaqMbrKJA4aWxfuYX+xBwoL5Q4dhkhyLePhOR68d2ixw4IoLz8BtNF/LH/mzIp
BzdWlPsed7zwN8WMPINs81etugLQKT9+pdjXM+zcyO9q38DJHRnh0gchpQi+bLKBszxxTNwL25Zz
6apVI4NIN9sH2QBs74kru9roBYHAXr31NBLTbgq7p/VdNXqfJySIJu5ANuS5Ovd5y9WvHvvOTtE1
34J5BNrlWJ5ZLrISM6llrNNjp9OCjEc5sKSv2tTQ+/xovhIBW/eLEi18ZkobEmx6jQ8PNf1mJmEe
Kf5+6sUa8NN6Mr5NSnKc6hv1OFX8oGjmw1ClEG3E3T06itIKLuzi5fY7mXFrSk7bSjTo01bEWVC5
QmlaohMExFHb28l61xHp/0WZPiHUPDffIeYI+IGzwko05pVL4BUGcubOZU3jj5dvp/wSCGK9NSNh
uLK76HgrwEYO23jlv8N5DIKFSsI8fP/3EM6RU5zTicW1jGxwNYHLTbUKUIL1wrhbvpAjNXLW8kIe
37jj5vsNOA46XNsFosUrqWZZEf8f7meLvAhSYqwW6KHsVLmz4cob9dHge6jRNMjF2uYl7BUXKcEE
n66xXmNiI75KTjz275j1VTNi7A5b3YBlxXuM2T/O5F4DTMnGoQXwLkr4mFI/P7v+GI4M2l0mCIBQ
+N0IYg+sD0Z0C6CjkM0oGJFkcFZGY8DSvhxijw71AV00Qv0qFdZ4t0vwPLj6IaifE+scb4FrICRD
6sm0Ml+hvfLRq61IZkw+mSkdGOhYPmC1sDKTpEaHaCQ3kx5sBA+gCLIX+5lHMNYlSma0U/B1WtwN
lhg4Y/7K/U739x7efEuh5ODg+8yMeKgnWyo3ja5D/b7FDln5RLi0xX14RdR++wPHDjKn+F4e1Elg
CcKBrjaWMUoirQFfnbZtHJ5kxDQRzpvqHy4YN5MBcohhAGM4mNTdVZdvj2CyqjS/ILpXUbPXnXAb
ninFcJ50iUnTr7mBdnETtBBBmmey+IrR72g52uO2vYOOa7Wfin7wWbi4NPleU6VFLzMqEK8OtBMx
N1N1tJDPsqTvcsrHLEGfJ5+cGIQAqbySHxDaBcn8JJZgKteJR9InXhzd9QlZitvvU0MG16ovfrGq
n/6rVhoj9XUtb+DiHRhb7S6pPcS7ftnO6P2Psp33wEF4CTNlyeg/ebEvJD8z/k9G44H7qVpW75T1
8FfRa0d3BBY3/4whJMNJI8g370mUBV1eVA+QtsviQ7mUCk50F5YNv1ATzvhD2hlZANbJzUC0ROpe
69zhEj2JS7B26rRuSIcpdqAPQMgADvQbniRx+Os8yKXv8s6kLWxMSno9onE82HHc+vQ3n2dA0eU9
vAJc3qrasJ3eY4oxx51MGnDZDNk8tZXm+rNg1bW8iSJOYtTU6UNTyOk/pY1hVnVJpuiR6l9oP6Xw
3c66cTEQsl29NrjIVD+Xksgzft/K56KiN3CGnmttBhNJx1I0WD10nmwa0Gqu9A6g8ENVmYdJP9G/
pbKqMyHyzCCG83ewvO63EQy6MpM2qJMvWQ16+rQZPki/pXh+HO3XgZip7e1vr9d+3QBxO1FUThgT
j1K2i7ndmIWUZRxjH0EvYNPzsfM2ky8HjKtzLtKG/ZXsxeQzZZB2yyW02+9e/wFijljb8EqMljjv
yIu83gKU1hJWvbw/aMd3xv15813jA7L0UpoiC13Ise46TBnETDo7/KqUOYKSXUz0mge8bo8NUNoF
k9aL//NhQFnvuD4XN0f9/OOEJnp+b+2W12dJpwm4So4vlwx6AqvO0PpBPeuK7NwyRqFHJSGxH88P
wYAppjvSq/o59V8NRiRBNOA+r7ucnCGVB4BBUY7UPTvg8SCcHAdTWxv4LEQr+3L815OV9VviCBRh
bXCG61A1qoEtvUQunjZTYewKBkjZaDav9my4RuraNlbL51ZHnLYD6swTaYLyPl/jyPaXsN+YttXe
T+gZcOJTvTCG3HYrwcuKoG+8HaN9Wjic2fs7YqV+g557V+w/IlX7vq9ta6zMRW25w27S3LnI7CdG
FL6QsV8AsmHsn6WDzTR9CSysoid3O2HADPK7fLPrh2UFkjQH7pxYranLxow+qL/0Tp7d0alUSgs2
27zozgJVuc9C5bflVEiqfnQi6Zb8fGat7IxooxiJ9mDDzWQtKYFqkRJeUUiVvU+lnVau1CzoQ6Qm
cI/chkfiU7TKEWRQVj1RtmcJv7cIroQtJdp/OMIsovUfclOHHrFwoyVJZfttz3ZYjCRMDlEmE1im
n73jI2NJ/kQyEmgxde1hakznT7iMBk8ofSlZdDYgNsz4shr5qQNJYG6jA5AfbXY0KQ3Cja4e+yWF
11thK4QtE6cr42pkgnPGAshDlM+FxWP3tpp9EsHXkqW81A1On6rmtgKWU7cAOxYDqFsjKqQDH9ok
arh6i1qV2zfMf1qMAIzhJFvwX+DgZPK53mMGjw8zZBmpYnENTujoCI7BHRCbCloIsuzg/J/lG9xp
ESicodQQTT35VNTo0j83LAGcqZuzX+ez9aQbvOfTQI6TAVuaNYXqrpB2hkBAe+5ZMbI7ROD93rD7
uYbp55CfVcnM4XOBBvJnz7VKEJ0VYN5Sb3UHo7nIN9m/sqMtqVwO2Au0O/8auL9e+i78ZfUsnZv/
0MDK+LrNHkn3SwGWgvR5S+O/mw1UwSiwoSZ0VyY6QXagH9H8TR6squ6mZvWOzHd6PQmuCr7LRqbF
Q/uJeA+GJGr3gPmse3VPQTZUz2f4qKI3xKyj9Du6jjWKh5GYGhavyM2wIApkm7Djqgg4vcK9gjmw
LYU61LwGDBXeJJlS0q4CUH7FWJTqTvCoXtvcp1eOq/ANppcQbNjgS450ifOeCb44id9PaZjiOgrJ
Ci5WyPT48J/dJRyHAvuN10YGPjpBUKvtZ2QXoWy9cLg62hMoVFE1xD1p67vB27Yz5eZkOHFSeU7j
DJ3rkD2KI0hXbKxLycqSqvvbtFLElwhx5/99xSuMFbf1qyTdGDMD1/O4TxWrMcV5tu1WYFOI3AO+
dSzO22Efn61ypHt8BbqRDjfL1FKluv7VqM8/4l3s54v3xjXOEdJia7+eBtUs6aNrK36yaKqG30kE
sj8cLVpr7w1il9jPKpf0Y9PN7eYR3ooxpKuQnPhIPqGiluP4Qt0XcrNC/Z+Uz2nw/xCUdNJDWb5R
t7/SiV8Mau2B6ndiiG4i3He6Ss+wQb8dQY7IwvPS+mA2N8absw5nhlslNaVWUIzCTf8bsqWE846C
Z1DHw87iuJePIQmmP27L+uV3IDdT2n+SgcKwvnvZqdePhmxFFw3CfU8u5aU08uQqXsVxIEHS/UNC
HyNKqH0G4K3kKhuyBjJCIZVgBmMwc2ySy2mIjGBbYwhFfpV/afFKV5qkQxAHblbQLuZxl9Hq8XQl
JqRUtCdkACHv64H41vi9CE7sw5P2ClSWdEZaYqHhDCgdRBPDtPaXVMsheN9RZDvF8toB2c+DqKSa
gvvSUg9yZquoXgb1VPLsLHXuNXWwk+is7MNunfifEWl0wPzecrUlERya9sVtU/5h0ysyiW4AFkuw
sr+wf/fswdCNfUYpt1mJM4veuF26LpB/IC8mOOylwzZo3ZBwccAFJqy/GnmGDC9ZObVWDeI3N/6A
TPpTp56FQyK92bhfvFj4Xn/pvuGRqz3m4uFAjXK++4J10yty5bleLyRD9gE5M3WYrsKq9OHfnFpx
bCKGWVAUuwbQjrX6bUkmw3reveiWKVGOnJWyQWLXQqWCi8U2TnHjDuLNzPv4F/HbJcvMFLrjapRJ
XrXOfOZlyKRju00kiUwMBhVbA+rkvvkNDfxfykrbAKyrUqAgB1XONl6iLoQwVuZWMLVi6OcrvfNi
J9dKVdbhRGfk5qAjFb99MpBYokUDNst90rFd62F1qZqEWfK2AmOfZcdjbEC8WW3H5L3IHuL1QvP0
CD+UTTej22zELWHrfGzA8Vy5vVx3NjV9AIM+Ss5xm908k4y1lxKIX0ptqxNlT2tkTturRjf8O73J
BO502wg841wDd5rb0NVJ0+DEx4ANwcU6R0x2Pwaspm4DlekllQp1oGDPGDCzO9E3/UIwbhivDQP+
YHtd5frqyuLigxD7ZRdDR1antwMYjA/5HHHZ2mDrEv1hx4WE0jKw+MQlnZ+dW9hurZ5ZZSzJoRD4
kxrEvmcSXNiUYMjhT4isYU3bVRzblNwz10sEhHiCRtUM6Lj/imIHoVKjEfaOtYR5u9gxkB1P4laW
0PR/MV4RGGDEDWBJQoewv+E2RovaqhCnGp86/IYhlZMAz3Pnzmdch92S2SsvfHIUXwGWAuuo1APY
9kqTWAEwLD0HhNYeVrOVym6D8AKek00eszVgAPQr7yfMtmQKX+bOvQJIKmT6Ah3KVyPssyDx68o9
Ymz4fSyUFBKL2XuqKlqgGegnN4GaI8B4ruHev++FAOByukWqP20Mym6O1zXr4eHlT53QB8c7gb1L
LjYj8G47YF3s7V1AxSBeh/sq4QgLrVrjPITAdJpW/UFOlU8j/V03FDVIjoYRvGcIej6M4J1/F69W
k5Do837rInJnvTWxWe3ak7RMiAtMyMsN4oTEROBVR2D6GiHOnvJo8lsm9uvnGZIwlElPrNjyVIFv
7u86zV/SXWaWNKcwaxQWMxuN9wLMBI/oOXBDIflEfwweSuuQkbUh3+OA5maHbWzgaoY3aMhhIMnx
856LyXnKRaiOZvX9925STs5r4DG2fyrsyUHRuauRh7neCquDEmOYCA5OnugLsTQVjIqrX8ispgQG
4Y//ArRdJQjbufrOdb8pw+D1p4tWfWIh4mJ0/26TyPLGpMsPZa/r5R1YcGbNlZ49X/svJwSXMO6K
9AK/ly7gS5wIPvHoJRLlUzydjwWkhwpf6invWcRDpmy9QkVGplupenNBk6BU2SKGA0EHsPEqMzZX
8AAzEHpGmWq3bXajMbzCG42YsehSeZDCFwa8RcQa5KKWJdz8Oyrnbo0vgQqJWnTLsAuvXcWQ8OOd
9Vp0eBpFnsoAG1MXNSuj68ZdHQvaFqXX28B7t3ESCA13yuXGLc3Xwl92UmMcu7sfVvZ6g0GUITNP
WwE4wBYbcsjp6Q30iJa8L+Rs62vtNIsIQkdfzzWh+Smm6iBAoG85NtiMuxkVoD2kig50jrWo3d/L
SlOZ9yHOk79vZRsdA2lzjckZiwhalCYrCOohrLp0EM/yEEUwuzKppySvFxRshHLwSQ1lJwNjNEBa
I2WH3cTjclVpIYAw1hKxl4K1iLRjj2q93+Ee6E8Rm4MuWBL+s2se0hOMfZjo8JKYFIFsvpP0SZMU
8RoebWVAoyCLgg124B4UoE5gCLWaov88cCz14D1bgcWhVs1lfivC8AmsUy9Espv1yNqiwURQHmFF
XyTA+eGY1z3H3TfvZ6Ix3XWGtF9XZcBmhTIe/6vm6Hx1/i0ELyCBVS36T66nqFZauhZ+X8KAI2B4
YC7yuoj1XulSv+tKZo9XTeC4PMIwd8xiNJPQLxOB/45SPkGfJCwnYXZndQV0THaYf+LTx/KF17ej
DmKbO8UZshmRGdbYJbDygXSPdzaa38a+O3BGwMFGvM7Ya5QDeAwWc5tRPxnkNEpfPeThw4ht6S3m
Saf+z3eNzgB2kc0JFidwLAQ8cQ7JHrRtjizNvPTaqY0ZpvZDrPRteerGeMzglRbKELUrr7ShqHD3
DyuwR1HaOItJku58IR0QJC2XDi77NCY1aChywLJWQG+1LkzHORsWNiHGRsBBftRKLQ5kJ84vV8g3
yu35ToetulA2pixmegbZrA9SyEzuNdxX7VHyKB5vuVydF+5AgEgnsUrGso/iBaQsHuE16nmki6jn
JVWSoHX+J4kS3X9AV3gQQZA7Mf5IeA5yfbASIl24nwOEr2b/PRHRWU2b4Vfyubio6L9/K3XoKsGe
cI19sZgvFkQz8UMGetffnckAi7BqymUQ+FVnXpZBBS3zYJHpVmWp/Owcxj58y/mDMUNaFeNd/EwZ
amCHRWFsItgkv422sUpAyl/YJhWerlzfXtf4OGccExhqhUj096EjQxq3QMsGc/81KWnBEcfnb485
qBWvbhuAejTwyj1K8hxTk9oLQ+KJs0eDj97QEnJpFAZTXnc0C779mKG97Oz/ElaRKDxAhVZzDb00
bI/caY0DeIhu811BoN2kkGwR+2+NheqBq2nGE1ErUauBOB52R+pQkRJmVI5O6tFjr6N4uXJS4D6l
lAnzmfidhNJCvNOVq2pFYxRvCNKIwfVsq1BO4MiQIJfwMfY8sOu0v5W8pT9cfTcGOxWrT48+ZaAb
LMPrfZgDNwg6r9APhzn0xjjgLbnJABbuQXMPFS6Dx4qLdcjU+64VRlcWjdSlc1T/rE8CrOXR/Yut
hZ6x2gpxZma4g/IaruMGvFqT0PgUJfEor/6Gmp62rsrdJ7oU+iIN7nwZSXlbaMK+sZxBX+1DiZZb
kJxRDuZZtIBpX/vHHF+c8WVWMyEVvkvc9I5lbND2GS1oFP4lbfSFvpqN31kHmTm7MHvyiA5nZt/a
d6lAEqefTBgosTxjI3XpZ8MqzhOR6vR45v+HzJl7hBm4p9tZ5t3ssFYWFgQ41o6dm3o74DOz+R4V
rTHLySocN+zcaH6ees9u3e+8WeFZP+DUgIJuaS/YiOzO9AKB6PAyb2hSclRGgcLTObC595HjTxPv
ZOjJKABXiZ1TSbjXm7I9sg/Ki1xfllR18fbM7nVSxKP+Sc/7Rcj4uWpEbL0TkmMXBxo8SaiGMRzl
RjqL1typPA40qujEHoNPQRo2/OPrqNTQh/t68NZrg5WRuhlQUG3bEZSRyzbK9wiL8IdwA1EAbNNR
7UwpntbN16uyLiAAECY5vpAzDkhX9UNkG5ChzQTfqh61Ugk3fJX7zveO+uqRcr/cNXcmbib2LVTE
yFT8P8KtlMiMgc8mb623YprnmeTSfhOJ4qFON2IjP654o7oX5jdd3T6C1PBciDN9lrR4lgrWl4zT
M8q6WzsyMsRftxDSSxJ1Rn/9ldXrkD/D+jCf31b+iEets8ApKCHZG0BYmCjTlcuvmCjrNWdopGE7
OvXFlxYF1LvvKoWCAdVQtM12+lUgkxIo3Z4DI+Smm+KK3RwJ1zw7C0SG02eOsdD3ESwRqrjHl0NL
jQAqAFayW0hDBNz/XHUnFDNblnhOTN13X6Eypzte6CKMOxvBzzRRpENSygORTFEqKHlCxW6S4QCt
7N/Vy+ms5NNimgsvXPN0qZJOtMHvCg1CuA+rYx0F3VeqMl6otehsT4udsERIbuPmn3iZH9ydprYo
PSznHDRiSMr4iLZxvLtVGqMMRgDbuGfr54HH83TySAbkzjAcviB8jUWg3zp5ECvpU/x1JmLTugk8
glTKHaGRZb7+gv9nMPRTrpAhxmFI5K5MO1i5MrjZmGdSDeEPuB+L4/la/fCji4dSSOy/mb7fhvTF
Yh+RXnLxqmyLm5hlkJlO5IdWZkbwtMSU3SdivXalCWGJZhOm7fd4RQ9qb/08oEtZ2OXQMX0jYNGR
0tNpOKNWBwgeGG/CBk6LBh0P8xf+VXaQV2hxrJcXQ/fmlpljcjHGmAvMZLmwGtTdJeuCCZdqm3cy
Uh+nHJA8YpAd5VE/o7NvkbeZzbfPLhUvAlQWni6vjPmxj/yCNnTr3IuIU9scuktZiMZSj43FqHB6
b2+idU7odbizb0PHtHso3ssuoZSblXbgPDL0Jhs3+akL8SxLomkfjEZMUdEYbEiMsLrYwmRxukxR
mkYGJbPkNXtnywD8kQACO+9nPRXmYl0miAcRz5/tCQDUfOdWGo2SKnH6a/hITocwyVOr0HujSsh7
fb2iy2AI5OWaZs5HPZmlBjMTn9N0x4tvsydYSrsw4m8jK86i1k5DfvMv3pcP2wgjyZpokwNbyuh7
Mz67c8jZHQkPDtsV5OK/GJafYzY/6oFnJ1xtAhKBqKy5LdsbGPvwlZBOjKVjWUm1Oyyi0AucdDvM
KKPW6S3cM7FBHbXWmYG7tSNdVsEH96/GTiEPa+8LXcdlVAh/lHTMd8jj7aglWk6huF5u4DUzqEug
3Uv9fdMpfmhsC/A62P5sJWoh0ErbDA+3H+ZjwxPkg3+/Ja3jMZe170dpC5X95XWf2atuNGlDN+Y+
hax468bO9GMbpk49rPpwkXJy2uc3ruxQLfRFnbzSBd3vUu2JrP6DXN29W+8BcX8/MzSsmXecTdF3
V1O0J+3WEAbIMwDiyXXdsbIWncftVc2vLOt+IeWfGe5fiWCqkM2MDmI3LuFWAkzibBl6b0Zt6DFU
zJoSjH75FgASDzSiwFENDgeSDlQ2vDeyvbZYVKWlxq7PD4WCFVXGTKzUktktmeAPErLFyh01VdeZ
+LrypGz+nP1/BPgNjgPBH/zUbiJhX+rxscs4nXxZi14kgrPoK3ij6jg18mCPTaDowdhAKXXwnI5n
Xd0foqOtkOrUxIvjqcRnW356LD0+oeIOirs0fT/fGMjWTRdgvIzJgGlpZOYc9MV29KRq1QC5Bity
T+t1HHCgResAGXK9iPV431vntRMNyzsdTvQ31ABuknWPt6RIcde52et+qJTvpfVzi57TYXKn2RGf
raEBUh2DoOR7sD2hFgTErjeJEweLI34517ftQATrcfunhRngyx5CpEP0HnbSIQLqDBV9mbpIhVNO
W52htxGe1Pk4//Bp1cw1TsstKAkIQ5S/Ler42X+4oY4Lj9T5ZtekeiDw2EgMWGnRutlWl7Oe6oUo
xgRcpz8G0qAO3XXTlbneuPXEfMitqUPmwRpDmI1nc/qu3E5L4ZEna0LQxGFz+Bbl5mwJPttUdnmr
j5C9N5jSmN47Zb/3MGeM5jk/qNsyf6wZ0w6duQ0T1eKkaXHyD/L8BeUXz4xvFMF+Z7qdaMyGFtDu
ZCirCXbqquvsXO3WdxiTkwX9Q8bXCkGhOFGGnq35lWg1r7dpPISa98NQSX5cMTrC2oLso25FNaUR
KQYVe71+mP3d3uOaAJdrOa09BjbaPKNa4NbEvYVnqgf//46w4C0bXJX+e45oIIJnv5RS5S9jhw/j
W2aiPDtmSIK+DwpaoMo7j+Kh47ZVNBfXHYCt91zJnohalLb/69fME3b6ALnWdKLLZH6gKkkJNTSi
gohlZHWLUT6FsIJidLXKvd5j+4L9ZS+xvwiFXC1JgpcaepA6MnDxlb8kRC0+u9EcTPFHQDTAGZzY
EO9ygRqPhO1g4A6gtnYbeehefEX0KSEHdtNwDN4JWrPhXf9J02xn6o1uey/+RpUu3gTHjqz3Xap4
VpMTfl4CYJmQvCmo77OiBg5TDeg5KZijkKTnvcnmHfJNPlFxcUDLEoHrF5AtGSQ4IP8OKbdzXqXg
iDTndjtNDwd9y0YPh9HTRvzFeF4kwt1V0vRabkwaHVkhToFftg4lrpbWxtvGhoz86g3UjqFzvScp
ZGpC/BteQ0i1mQz3MKHFSnMKA+ahufy4dsJhvxZBBWteMUkqqF2oKSvaeY1y4tpG6nsiRIl6rM/C
LNlBbUugDyJ6SN4RaDg5yfTp+A4D4ogiyD/Invsv+xI48bB+OZiTGqp4GnBcKnAWxJ8/eDUe6YY+
j3y+9x8kP/C5ZAZIUWitit6Nq/ya7xUcJAq2f2iwqeMWTlGsnU2i5sgzUHkwtDcm7uhyDmf7n8Ht
ic3LsgSqFszP5vHkfptwti47AOY8SLmr4aUfkTmWXs+PUmQmcCg4kG+WnmVGbKHlCHsCFuiik94n
8vikMfzrQ2kmbOssfpJ2yo/mD9sUVKAAvSfcwRLb5NJcKJWCsadCb13NXlUM8EeZrKJWTGNeNNNF
15xoFYzTNuO86fAsUvQD1hgp9hXOw5DpcSxZjHlZ5wdwYIKaVS7In3AD4kv7ybFWNxGxtf8aCnnP
hlIJfSpBqWGHibdPjEoyCQxH5Y3CRqAOEWuAuV5tpYW0s/npl+JHR43yJyTj7obAQk1Or6JADtuD
G4BEXVT8DqnITvzvqi84DtgTpuD10wURdLKsW1EtptRyPb2oFiPqAHvDDOu7eSp7ajUdFY6Iad8p
G5aZOuze9JKXxkjUF0Fp44fS5cMXDKpCWETV1ypQ/l5MrPI23ef1eoqjDAoZ+dOqscQEUzEAR1BV
HXyoXTRhpeeIGKZkp6ECWke56xvXXxMN2DAhbtIwdccSgEm9K4EB4Rz5VRT/OTBwpLvJv9wV/+3F
OWr5inKLJZaQwOfFBQL6aMspU9FaPKFWOfbjhjuB7jx/Mb8tPbCGtAQCvKdWLiQ5Mj3XfdSfq8Tu
pMO4hk96u+4Nfr2jHEYtNyYLM0EH6yMMWy5Ux+/OkTe0FD0THxHSrZkBj9up4NlMj9PRBGPUT9a2
mcsjq2ihL678rv3Txxtz/K4jfD8JmVxyWQsqSOqiuiOUsoLNvX9z1lTPFRdRMck9EOBtAnHfrQxD
G/7rMFlCp+WnO2eTWCNn8jQM0cElo6KR8dsLfE4o8YDd4CKUzBiaPkxay1EmnVCFqHPQA22ULP1f
oUm82Uk56y5b/Vv5lWBk9x10mKIFX6elNyCz9t6bEsCkH5i/LMYJ/q8oyo+K6MgF/lKSB+ahGUrd
ehC9PWClmcpXUS+WT3+wLXJ24RxTWEO4mqnV+lyjmIHgbjV6mNlAQGId+50mq83CJpT8wLUPtxSd
f/uPMGQRE4NmcQVO60ROhYZgERXdpVAo8Hj39j+B2Co/CbcA1K515JxbZ6kj4rCuXF+rwK6NWm25
ZXifPqUFsfKMghcHW7hJcT0dzj+KFIb8w91ZGKHONCdVb/+CZWNxAdjRIeX8InQsroK/2yunPPTv
FymVl48lGcqZXT+CDFiDu+EWym3ln9xIaw9vZCn8R8UV0RfMrHi449KOhJtDIlalScnjdJ/Gn28f
swvbeg/dYGGrcD1Mi4V/KzBodtwkGYVK9Idt3Vf2AMCTDHmNMJnsGXbMhH11u44SJ/qCgRuqmUMf
19cxWDS/XBcSV+a1jcOr7IvluhB0+JsfQ1iJcPSETp1igPaGHMBnRUNXYaLHsvtVzF/ZALKUQ/44
Xcc/YeG7p0BqUmMjBBIutSdA+j3vEM1KLs5ISD988hqUy+j+94UA7FuM+JPFUrFXuwdrpvpuF0Nq
fCAE0UbdhRV8cJV2zk8ra/9OGY+vdUSt+HXdvbCvkm5P51FmcAevwSElhx7kSioiKi3FRB71rkfc
zvtXmODst81yxoPEfoXbsN8vD5NQnp8EYOLxUjCp9RJ7NfgYbrcKj5WE2kNiHWFXsdCz8rBNnDBY
OWYt43QK2mFwZWE4+k2ESQJITdPz3pFcy942oZ6xsv5yKg8+5bYLCMAVt/NVLLB4ZTHw/hVlHY9j
Ce3eIFhPriQBHt/lUFDaOWYC4gpH3qjyv6vP5OV+eg6T4BkRg0g2LXRSRURyKC45g2qmWjHi++Hc
3U0vVVBDqC8lGbqOfu5khlapyNho4WkfmUwvs9aaqmHUKKmy7Tcwd6U4WTUsTPurk0uFvxgOOsnj
DVS4KzQ1r32wJaNY+eiqk62oALdLNZZXNi1Y8aDKErJ7ZeXHm6o6Y1Uac0E7IaX5cZ0Yv6hbH2rl
FC8bHe9QdsyGDbyBf4WaFLEDNcoRW3ZjdfJdxF22ITVrirT1MOlaguSeKV7BYbWgqwT74O3QsoQC
/2iLl5rv23BXZeRotLOmCFBjCpRbAU50pwrd0OiCgcrPlcNon/vPHp8IzmhRJDDHd42/ij8UWqMU
fa2vpvFkTEexcFY3F2mQpBQPb1U9DuoqDapdK2N5wl0S2luGBaK1Ew3VvUTlJin5zoUGpDg+tKCx
eClfOyWXDohqeRvnHXKuJkMkm9v3bCWcArJZZ5xLnZ+yin6Ei+9g+SjNrIRUDe2rpUblYJKO+9BM
+EvCKBeKCs2upvgEA5pb61Zfa+yUBVMhMgs0yGQDLcqCuIsuP/9FI+Oop/cTvO4w8xFnKdYDLpOy
2trdeGANLOmcmKlRLuEKKJdyFHKZrpn0j73JczdMEshUcjdvXQXb/ebj23lHf5lK3T4Wh61mET6C
J6Q+FETCDY5SwZ78t+5gegQ0Zw/KBCEPCMUZ5q2MvIHBNZx2ETYO9whzybJmvJIBDTOzQNoA1WXW
mNylwkMZeHpGCpArZaRTMgpDTL26ZgMy8P0h/6d6pJbKb3xhEFTTgL+MP7ONJrjZ/uryyiPIF5M3
scZDDshCVAYBmp5SJS0PMjx7tJlXemoM9cee7zO3pmnETDupQ05UElxHPGXSYb+ZUzCd8QAr1+Fx
+ZeGQav3RtqK85lnDx+Dyox8C77DDUpojh2CxNKnKVPwLBW6d+qrwEIOtx4Qcvg9S4MqzF3Olkvj
4I28r8wswDnmeBrMOvQ5ve2FRjqEzPX6ZSTEPxZd22KxzNc90eKaVKSMG1qMzFJFkgUjzaUv64GU
zc4sbEaXUsVMoSxGWJjX86kEkgSaLuNNrR/BXtLe5QvtIqHMwYLMez3mfisA2G6YOtlceeDlw3LD
5pvtKJ3nhyXhiREHt1gkl2xLfyFdF7YJC2UzZKwQWLCf820zPJt9tF0yc4x2TKOJ0O64hphU0tBK
iBRoMj7HBPVb0aVDoO6gKAn9iRqYDR+xdE/zFG7dvTylCG4j5jQMCV3qT5jLWOLzVZqNwhRg7BI1
V1xCKrF5/tqn39irw1XE6D7LRZss1gnHre9gdXL/owvet9rwnWUDFc1qtaRmu+ELaIU9u0i0ToOU
7q4Tni3nw85qk3EyeAZqM4bDy+B6e9BxWN6rRHfC3dpsPHJmEUQbrs0jj/5BkHgVpbLWItsS6eQ8
Gif+rXptwlakqvWhlFYG/UH00HRm63IF7J8maO4DGnJP364ytmMbEjtZvXGZxor1Rh2cdG1Ylev8
yvHg/3QJKNjQIQLJXKi0CcgGrg/+pQpwt3XWPfc7kI0DVGtzWqvIjSKVF7hOdmDYZX0VgJRVChW9
crWLeuanl8PEvPXzfEqZ+vImIc0rrU9IMwTZNa2M8l7uULTS/S5cZdueB1I6EBYlKiy1g6rBCXQz
pYkGcPpDemw4Juew5fXOnKGQupBcqFHbaUiDt60A6APTotN4V5LSpOuECMMD8peeRFORldxSPKTj
KurDhF3V6guaytwW1TFKRLbrPzGHzAdwUvpfPB4tPEJ6kENzMalWbP0u9hIUZ0CrQX2DclYU3Ni8
4S6WEiwppIdKcUvMpZBLPrsqImqu3m6autSgzB6Tx0p4lrBxCCjEZz1OBRxoQ6KREqoY3vBeyjSz
kTl5Fb4BzZMLZSbcLRTXP6iVKvpT9GVrSghdSr0nDDyLi15yUCe8JUoIY00s8TqKEI1LSNWJImbl
VlICYzbMAAIEukHsr5vGPP8L2bCOHcc03QtFM57lV8OPWUgzMewncj5974x3kAwCCAs6mENHisKx
PixxRSu9UErGww5/KYZwEBEs9G56GpeyGJ8Icl+shQIVbT3osd2w56B49zAophrarujHBWYkMqB2
s+7yOUs04W61Tlp13DhfRbFezvW98xOmWrpKt0gkv73AyZwty/0PcoQDd8LSroJVFufOWGC4yySH
QyPU87a+L7rRJIrUjxT5+YgZOqoOlBrOZkA/XU/MSeSnFz6fYDV3wh5va6QH42AWd5QtfyFn8wEE
duQhfTd9+zyBNtGw37dm90v0EGQRXL2AuSRAmclMKk1K8x8lDIh1mVEFoomo8WL802XseKHEeqhz
1haHYdyUK5AS6vBl3jMxS2W0/y4FRmLqaXQ42oBzZmJ2OHUKQky9Q4LtFuNpTIQh7sg7sOdX9c0i
9hDi+IvKZaL0DwAqEAc1wREaQhV5JHUzUaFAAViUAW4JuiwC85zL4jnVtV8UGNJiljclPNSdvEMM
GFsqu7CnbST5lTlCzLuNuymwY0OSFNPRi8GYUeHHhYIxdzd5lXb/e4zREj+Bcs+kiBdMtu8oT0ax
UTx0GJ7E67dubOtckaDjIm276O3JQZaHhoOgyKb/dxd1eRzuJUvHDuLgaT2L9eaQW1JQCN5gcYSE
ywyZu7aWYoUXgeFY779KfBn9t/8DMzTyIACkVFKYl6fcwPOs9Em5AxQTE5bIyHiDzFRm0zNGIHUm
Qnh4gqZfbzYRSepUJlZBIURHMO7nah38SUgF9NYCxfMuVP4bCK0dPYrH5a5+aeUZapfhc+0dzHTj
pfSSRG+hmaeLD/+CGNoZpJOk7VzzB0i8VcHrKpYY+PQvxoQApJgo1w2ZI9e29hMBzS2nk9SGhGAs
5Ih1I2S+TM7DaRblKA0R44f6ypzO9dJOEjSRQ9lb+RXd68yF6AzRq0m4KVDSjZLc2VfcU8DMxgwW
vN0qsOkRVxcVchtnJn7Hp779S9IKkBVTAIsvoB1jYvJqp/1+N+GOSNB+bINDEpsANqZBM9FNUOBW
+3QGmNvGIV66Pbug+T2LjEw9zSdbpUPhZNfPq7xEdP+gAm2IHuA5rCd8WVqlYyTvxT8jsJqZzM6d
oHj2JhpGn0SXsUQjLMKsgNpziHuHwQu0gNOCshY0KiwM+z0WGcX5p8N5q4Njc38Bzcf2tNXyHSim
0uX5mNWPzDFbzIS/K2CiU+uDEZxoRs/MYhKtVI0VUVyQhztE1tQ5YBRDUBazh8X2EdoxCDrpxgmz
3g8vcHb2nekqa+8X6fJ0qDqi0GE7QLZLq5Gl3gTyaRvGV+vLFyMVskbRLhvr44S94uO9J/D2ezM5
x7SkcH+m67BTrQJD6c1KkL1lLqd7m+60OMtpNdo8ZvNxO47ZkrSp0yheTYjpY9qhe4oQpfChWFR3
DcXbO2dcU985cr8FruIs5379WMoMfoxg525Sv+TP68ZVK6/kI1y0EnKaUh69zZJ3u0h2CwqG5C/M
QB1zeXj3u7n9EPGITioWCHHTIy5k7xprvfygzWwTlU/hyuNxnfgY1aHkW8ckm6FZZLR9X77bK5bG
XmQzaQj31KuF/IMtFevNUSa54eMXbJhfeG1fQ4W/6BZTYGxauwR4XqYKa4ZM3qTvuXZ6t77YBPMe
cWg+90Kxud/RV1bIED/i4QVBZgXLdMQ4Y9AR+8xnf83cbcWTg70jl3RQALwhuKWU1R9JO6CdDztt
Wb6zaZJVEu8gzeaJBi3ZhyecQxblTUyyRJWj2Nim6q6OOeqHCl1aRe98VvjuZEpKgpBsBRWS75d2
a5rsF7UDhcC6Ng186oP0VJanXDkLi8MhUPNWE7llpQXvguGA/D2kixSE75YDkgDpZviPTzq45Jcp
50foLXJ5JFE3wqpaa3OrLXRrW1L/LV4SR/Yt7KWyK5GkUQAWmqg8Pbuq3QO62GyJWTZMRSeeDkja
S6RZ4oLlo8ZznRM6jXWNRdMlNEIpmms9tiaoBQmbaaqcgQJkood+8wXkqd89KG7+o2hbC9DaIiHH
5HepHLg/rjLb6LGHyAJsS5OM9vnP33IMTocvC5p2H+C0wlW5V0a6MX0YA1T+Pah9y854qiGv/1xU
yMX8jOioxE7DWUV+hWrhwKU2DAOPxB4SHgcghs+attMfiDjHZqHztpiqEXxgWHxFRhFg5gaqsGBZ
xQhb7EqEg4IzHEWxmqTjfm/KIh4wmlr1zqHydwWfLMDJAXLmENLf9VmduGsZ9yc5nvHkh/EisOQo
tIrYZ6sNH0+XnovuETsKHi8j381CUX7YXOHQgGPhKFb1yWyF+ckiNoKfaMKu4U/g94YCWgxQYs/U
PXt3w10K2G8/cTl7w4Z6D0hjmhZa29cZF0jlrV4uCi32cEjyMRfeSCS+2Yxdh2RR/pDWJGwnJHFn
hZfbYNEd0G9I9JH4JEZQK7C8Vq9YyvR00Kf5eZgXQEOPUQfPblvLRaD0DtZSU4nO2eePwF/GEt3J
+QsNFbq6k2r7VnQ51qjrXq3K5CorFPHQ42xOn8vUVWpOWk+pf4YtavX1SosYCbi3pdbWuG41RqhR
16i4wswwRobdJVJFaSzszpslkg4xHM4/yOrzzKDGMoDMJjJ3+xwhaBvCdnd5tJpBSfvG4TDqkZNW
SSjWb2gQkMxkZygH7N28UjcobZPv9qp+jJJ17+4d/3BrXOigRLnq10ao66yCJU0Bi7/DpzSRD/KL
Dvt0nhUauF/bgduzqC/zaYwNT9qY8cASoEahWQZX4rBwYDi2m+d6waHd4JZDaf0XOvn6eqQ4Lwpd
cJYQ0tlHUI+LY54lkJHrgPBLzbJ0GbTGvJMbiuakwSg2Afp2yadIUXXFKUbAaCJJp9Ac5DoxYP0S
sZi499LbUxOMjyduO2eGtIcJAhQGVcIfd4dbaATxt6BuvJeEyt0llvy/rA8e10Fqm/8j2ikd4Gyj
hZd1N/i431Aq7dHU8h6qzO/x/f5Bfs68ntcrMB0nbKATSlPbti/dlTBbIjWEUSie+W9Swc0Cz1+D
HX3I0UoMf6Tc1CjfXcBqv5J4FKybC+Cr3zHV/8zErxg0DbVb/ADnIBJN23bAUVr0TklfFzkRhfAw
R0lE5pUz633EKgYKN9JCO/wseQWobs+fkapW0XodgUSgDGDznmQqiBbHc24tu3l3s+Qz5oarZV4N
aMo5ZYQDXu3XZloifG/c4tQe50EH/soqWMWK2mH+AXluyjvvfXAOfFFAHWxFICZgfvDokgX2M8U1
FB3XVta9V7QcN+xAQMspnvPi3Oz5Zr2T+ea2ZhfHsIgWj3/58oDCSdT2GJ/DQdTy/8B0vCY3piAu
wul9DnFL+IJ3ctHAN9wicI+oyc9KPS3Y0pJWrnKLd+fYiqgfwHRGf/TinlEuZshNiBaK6BTOUxDA
QKOpCkGpn+bXTVUeCMC+pLFckyI/i9vR/e3Si2/PcqcC9XDbouFNwztUBQcko3vtuoadAC4oqvQG
KI8aWMNsVTOaUZiiWBmXQ5nOpasv/wpdj8rantoM84sOSWEhSTYF93dhgAlYSYfQvmyelFnRl/8l
uBSmRh2X5rJLP2n1iA5mir7Qi8Rh0fg6vRnNCkD1fxZZz/RtEcKcm978f5oPdWgW0tht7O63Ygqt
gfLsMouhZ19H/gb9Itxgo3VC/7nhRojiDjFHmA8iAYLu9S9aM97wN0XjBRGZ4R+dLQKweb72zDr5
jEyXA3nXgxgIxsnnoDOkNqgWZD6BY98Ij+G958f8EAELqEkW36CsdAi+DWBZ+YJaQbJt/w2asR2f
npPQh0QVDqmg2ZMhZPfMnQa8zZHZu+RZTmf7fPX5qTkz4+YoJY1Cvvf3PcRKKucriexS5H/O2ruW
9Uv5Ms8usb+JsJuAB8kPs7SoIN9tX4OWY8obpQOzbudy4Kk5iAPZ5gZQUIgne9trr04zUYvRUiEw
XvOwPzwtUHblpn91IgbClnM2zyELHI6qi83MT90oqHCrkRtSZEOg0vOV6+xN2hqSlWZAKtRP7Q8B
rGhS0DV5EwCwac2XUAzkRqY+0qhvxLzaPKKMLjy8W4NxQS8wcCRrYUqwGE1C3xLeDL0SogYSPfIw
MpoQ2FyFZ2U2/yhejhDp3/gwFyzyhggGU5yaJzRoEiQJe4Li1VsEBL7HOp3bf1zgi53Y05ln+xJe
nzwsyJU/o5G4O5mJvPVtoV1ih1Z4iNG+VCQW96MErzs4VlaTqb0IMFsl/jlM3Xp0lmgNMyveiEBe
BGbAOBbQ0vTsVZe8lxH5ctE0VR0GLuogHR5Xg7cU3qua4Bf1Y8yRFr94nYC0Dcg4QZITjiEQMNBY
9aNBpW7sAQu889Alnc1aiRMswWYbwndGHAnK5LyP2KHyBsCGoiMG2d5rD/29EQTuqlqxqhbwCaS+
V67T5j4hZH40mlcm8/rs6We5zc1gEbLW2KzzbGkNKleG2KKX2DKKhAN5HB+PbePnZhVFD7T7C3mm
GRyA7yF0u8I7Rj1eMOdTZJ3hiPcobjQKhq+8s/urFFri/C5QVrQpZJB2Lb0dosFRX/00xfb6XWaW
lLlsBxyR0UFXQT3pn9GMYxqi2OgbG72HR6gdQUswAUzR6ywFI/0T5eqWMOxFiUsSR0TxEbZolry0
m2axLgAfVR6vsbsIIk7GAQ0nMhGbRkfkLFPs1HrDIAlc/zI2web3tvHV6DTZAui8j+zrtoNbfvLw
dEVaR8Iv20aP1VTLD/VO5FvK+fLTFC12K7zvbJ/sE9+VobiLINdxBweyt8H6dMJrE1615iF1jHG3
Bt8aq8BiStPbmTiyxOda72ho5s2LaB8atq4pR+w8OeG0r8voK7J8rsQzQlcrVM/Fl7box8wHbLWd
EMM7dF8s3Yt8EfYAh9umSrXYoOKM6LJGFGbS/b8UIeIsVm11WXq2+im/WJMi80udsyvzYjgnDgBH
dqGBWlsO/EFwVZtmp5vvruR7zPz9/coyg06t/eBV1R/gr1Z7o+hrHRIwhSI8la/PCYZ2EJl72I1n
4AgSI5DqacB/nSXpls9x03QRiFdgCBs7UZeaS9lteycivI16FrFrMAUDpJ+2eGq8yk89X5oABqeg
s6LePJSuCfs9L1uv/ReMQCGxf7F7REw+OPEMOgJWfzBK4QdTfwCYE1v4xAKUFA+JLDV4+/sRpVMt
ij08IkvXB+3sKWudv7GqDF76nHSlEoHbQwsVVC5NzEXXrGFygWaIRK9G8tyTrv1o++YJDTOykeAV
WsjYGd7sRCTW38/Oq+MyoWVBcCbW4nA9j/gtgIdvpuQrND9KE4O+ta/hmdG/r/bDcOV04OKVB/cJ
fT4uEKOzbMlFjKOH9mIGYZvr9Opi0IUhGd+MuMDStkWG8/qljw8Ul3oJNdy91AmOA6+71xsLKZW8
vOUiXEkNHMY4RtwAOS5c9ia6XfwmAbYrXyRvIZSyKAf1xUAVCVukRSbnPXPeLT7nBevjoiEudYtH
WwM4V8NhqkPrP1vLmv1C8Xu/FwF3Lwg+u2GlFPKdQuenWAjV+1kdrQfgFvCzn66eU25f8rJzsRVs
PFpBFmkRYOmqEaZHcbLQdEXoge4e8w4yhQHqWMeWkfEZncmXPe6Grat9T72ozqCwP+3YHhK2q2/D
ALUmvYwlhBZlIHaDbizj+bEPb6gjwVHWLs9LvUfz2Q5h0vwuHHTIwnKIEf+FdyQzr/gDd41xuEYQ
Pwm1aeI9DZzlv7MrPSgUGOLmi7tmgyprNGNtpULeQjNrp6syaar2kZDkvrwCNkkE9sEfO6FmXUY6
gOmNlNSoSWFRFqVCWHOxrtxigQ8+e1o3uMDqkizLV01SNOy9f9snOp9JeWL/lO01V5zn++QzEGJz
rweBb7xsyUeH3h1A9mKAgfKRnXf0MkPi5y/mfGz9wRVeC7KMN2zFrhOg7m7l4UDbsRERtfd12Cny
TbTlGsdQUnZusrfFqOj/RmlqNU/E19TGsXI3gEg+Bm4+uZVF3jwAQzkDh0/M0US7asJ0hq19FFZj
oTzTogJMZ8O5np+jiDEJLboGc2hpDzDY0AO7HirajxaSlBmxE2UgMsEGm5nAbZKqAfII2JGJWoB3
uQxI2/5YNG5jAWFiRpczFShnw91mh7yLMoa10HAt+gcEWZr5HqYumM6i6dDh59oRmLg87t+kaeO/
wwPfPtDWkeClhchbSD/ZZ86ZsEUJIXbLM5fdugUHh26yP5ZsD9ZYP/kUXhM9eGDcTTJYsJvsnwSw
KNTJ4BxUFiVB8W5JyzWmdpS1xT8ytfSXY9PCEjZDVxrRh6RFAIvgBVkg90pkp9iNaBfaB8r2NJ2l
gskxrvGFLRrP37eebGO9iVD73yE2I88jJAaASAGxKSGCP1KgKZ+dk4J8pxKNJXBoHYQbYWOY0YQk
uv5rG5gu9Ms4TCKST3EMSF7imilq46XwrwyjRga3wTiSLO2/mBrJlUsz/g4uhFdK5vKqpfVHV+vC
PwRmt653KYs5uy/OXJMugU3rISUFDWnCAmxz01lMyiwGu4mBnVT8bCndNgy7ST8XXMjt4/2y9xrN
64aqFDAwdxvqc0qbIN9TJoEwDwndEfnrE1HhPnQX7lweO96DexSRrk4rvGEQDLfjFmOtlUIT7xso
mx8cFl6xYB/Rug52LbXlcxSi6AR59z6VeGh5sNgENDSTDJ9C3DClCVxIbNzmoW0EpvGZts1W8xEj
WqE2DmSFgNERNzwEyaQ9JrT25pxaBWMhoioWguPuNfj/jqwOLS1igfkQdXgWt2syihw4DqMi+6a1
wF+ROGI/I92u5V0rkaY3Z2ZyhfaH8H+h8h8xJKAlgxoEs7ccd5EPpG8X1IzOLqNEdPUq/ACsO8r/
2u+UR4j4tyI3faGdRRhA8tbAiNoSRqWNXLhnNGnPJESGHpPEq8VBmE1gAzbxcTGe6vq8JguNilQ9
5rQlW3IXP+ei3++j5ap+yI7GuiZCpTGWV+F7bjn8+mlR/im+RN9IgKwqxoDVhRiT1iz4rOHeyD1+
0d0nExNlMTZ/dW7XzG47m1FgU/LWtlkPT/NgcyrK/1V1OPFfPBTue24CCY1jDkK0N8QtHeJvO1zr
qfaeSWZUKc+PrBORkM3X+uQ5Ab6JgTklKNas+mVMg0IbVL0J+P3/Fwmm1UTC23qF/Nz/M6YIQAMa
GszpeDOmo236hDteAAAZtto1LUALLq1yAHNfoItIiwexAiCRiZN+sytOwxthuTc7JT78HzF2tTre
7G39a9Bm7JFw1wsv1Xndd6pDoEDXHJIWONf966vu/0cE98I41LZtw0KFF1/HFqafPrdMekW/tSv6
ie8kK22RNsR3M7oF8Q2/SqDyXRUeXYZXz96Gt4JS7U/gdgYUbA/wL0NA08XGL7sDXlkmO7aV594M
fl1chc6LzyWKIwTgTzNMPjqwuXAVm2Gxp8/mUGzTYKkYOGJdhE9pX5bPuD6CLSNBJ8GAequVdhZy
PvQD/6khx0a/koWl4HsNAZXCVbvLp/NaD2+4DLbZlj69IrKNOjol+hWPG2ETAdyuZRm+Mx/iQ/j7
n+UMxZe+/y4bs63UIGbaKJHzaabkgCMYFmBFIXHHFBnKJhPD54BIS7Ar3zYOxiwQ5cdnW7PGoNfn
mpHvwR/tj7eeJ1sjOzfwHZyPj836xwI/40Eazq47Ror3acJYjmpIO2wOXBThav3iPvvJ7+0k9xrU
t0RmplB6vd3bhu36PdGRth/gsIRmO+KLGK3BgLTnVnwIKh7NSCosjZ/rbjzH+gad4SwrDRJGQEXW
7DIE/UkYWf3LQRhBNwN1mCyvnmA2fOD/ErUGyyRIQBKUGFrC/EHG6PjBkJV6t1Mr4uiI7cSLiIpR
tm3+Ju+z4Gjv+RYP/BYwIXYh7JHdNQCqCYNIa7AaMI08NFF3o4B5ouJMFgUkJQfmiGw5zneOqkbp
QF9ILar40pD6ii3OUPWTB/zVuNZQPzrvpivm95AFKYWWDEFi+MNseXRnLWXXg+UI3dB9BTZfJtAK
Ko0HqI7q0Gokbp/woBXBv1L9dAq1y9ydfg5nOXHvP0TTq2hRnDOjyfqWB9h8sL6zxoXW3IwPmA8V
2hRl2yxEkRo3vUdOWTXfUOZh5s4Je+WJn0zig44rIOvX/xMLhwlgPLcgQCjDvr+zKMs12y3WSxxZ
/mrz1ihyNy5o9bbH7BQkv+4rsYUK6rOrC+EDMCEAJLXkGppDc4OdfxcRKSf91dzLIpvNZo9iffmc
4SdTnrfOhuaAhWWohwMmzMAYvQM5yfJGoF2YeQsexWX33E1FcdEFbPIndbgMZVE0ZR0ow+0qQIgo
a5Hp83SHLEcG/efjfpxsAUOZJlsCasCMJ8o7ezjHPIUt9ecSSEqUVCKvP1d660p2HRzh3C2IJYAW
6czISqQPTVlTNet/dvGkAZCMHHgcSfbhBwdqN3q6MTc45t8HZR+t4+T1po+cnHAKPU64pKCuEuSG
/MBSHFJpst2GRqca85Bx7+2qZMioD/+UO5KPB+dCZJf+GelzMJeALu3zopr+TscmGIAsMwEW7GBx
XoT7H6OmmwRYHnUXq8gpH3uKdAjBm+4NoX50DN3n+Y6Z47DMiC5NLv5Ukp+PGYBG/3DcDuaCtg5r
WG/TAy25N8RQcFcYe5vTTBxH/oA8AHbq9FHVJ+6gx94/ADM0CGH0o37EFagzNF6+rp3ONjfyXZtR
UcRkoiJS1Xs+7y3Fgxvx93o6CLVaER/PCAm3rS1b18eAsfkvdWuhjCJqSzH2R5yDDGXQH9Aszxbo
OUQ+GXsu4Yh7HtrGz5OdnsX9LiJDLXqFZLrvXws0cNkPiWhTjneXk0+Teov0DJNi+Fry64F6evye
nhMcKxdP5ebwNs7+7BXrt5ZsBaGT1xsBBDT2Ko1QBA6XdkJf+eAvr+MXh/yxU09qegMsSzMbvm0B
dln5D4oQsQOI6w8u/BSqEqNzGL/Yy5HNbISw0PW8TVZaZfNWIH+VFm2jXFvif+lzFrjPUOYfSgV8
LQXt+uiQsV+aNEDv9RQyCN2brQtmE26B4+roLMkeXNG+iSV/4/xjIJf4EFpE5rd+YeiVTGVofyaD
KnlGycz6U4XvND99Dc47KxIJyeE1Xg2Ck4a+CqPgyXqAfTy/AoHcB3PZpKmtgNiHqI/SOXH2/XeK
RjDisWkC1mK3iNcNlkYRqF86PWDz84sxzUUWL47cvLt/y62DAXVBgVJbOCHOfsjtL4QsKeu2DeUX
KH3znzXWDJ06QHnV5SP2HkrYFZrCDmzPH98hQ7c+rllmo3pPw/3DiTREDThpLNhNG1Qbm90/bbBP
2H2p6MLLp6rLCpZfUWQW+S2zKWG+wYFiYRoih6e2bws2/i5DgHHusdh8sL0F/MDyHkhyKBXj4WMH
Wl+S7+GqWIAmdsPNlXdNZNafWPWGeGfDYyz1fAWOb+HwmFQskUVjPm2xr93F3CVRIAQNKbMJLdIq
if7/yGB5+Khf6DLuN/hRJTF+rhVqKKsdK3k2/wLmLalUmBagbvBOvoAKF04fV/QtY2kbeHuH1gNP
d7d3PsHKGWz1BPfjdsHTX16odim1gUphWw/wSxchnejkZIfDy1unlPZaOCB++QwZOAlv5nB8xBQX
XBGRgFUNh6TCtHyI5ExL8AZoPY9i/ZS5WM/SSRJF1mys4H7F+Y+5w5uVU5AKQpDAf1vZfShKk/aJ
iCEK8xDOpyfAHSGrIHxDDb7XGTcNvGo1x5LeroazN/xjiGAYZpe947ewA5lmFE6Wv0CwI+2+4R+f
FTgdG4mEXpufFvRb74wFWYvP8Zl6va6StILMbRWQMwgc1FxGzrKJeDtlR8mixF1J3zgbGNrAFTkx
fmGBVISfKt8wQnA7KwwES6+mnJgHNe6ufRpzYb8cZe3xtMuOHv3Q/30OiFj/kz/gOiQoEfFTWe5w
CEbMoQHu5R0Q9OWLwKMbzRLyhY5qeIVtFe2lkYhIcArGt5UYPpRGP32FRagpVJqK4ymqHOxSeI4o
qHEDzUU6TccVBJE2L7UxkUhyzDNRs3bkv4mk2G67H2oZZX2pPlAKCr/AIsdngVd+3xGWvqMn6by+
3/MIMrOq0RLb802FL1A6Xt+3dh/KOtTU1PeEXhnT3vdWUzRX+tu9Q3NcMg3jSxY0HIcA2vNL4oim
XivUqhb+80lyFgm8yuFVbTGlzYiw5t4Hq8plHMJ6nYdZaSlbm2AVLfjqqm003d6pTh7XEM4JYcwp
KqDCr28haLzEwq8ZHIE1dHWv3zbAkr/cDFn58vJU1GGcUsaGUl7kCI/Hi0nu/SwT0U3KrJLuhial
o+YKy64ByaAhAc79L46jqIBRQPJFSa/Im+WzGZpps6ysr6BOoaWEIbUgfHziI6Y3608BHo98YgZ+
8v3OCouhEECUeRW230eMbQvh6tnjQrrqQjquxy4EyuM7oxavli5ENc2rFIFmhAvGElQgLtkooo57
q2hS1VBZW7oPvadt6DN1wfog1kizl3lVtWyQ5PIc9vnhlsGBtu8tFgCOfk+ijKe7NThRqkx2y6Eq
MyW7daJoQOLQ9ULsuHuz8PwA7Ao85wTtp2LyxG9zy2MqBAy6VXZ6jcFh9Jmk9/LgmWBcVFJuZBO7
2FkCqH4P6bATKJUUM/QxwMAt1v18fXrsXc32VHzq7RWAxPAnrWOL94LJVzDbb78QpWF4lA3IRFV7
kuKQ0V62I0VLF82DgKz3Nj5a4Rf/8AsI8RPOU6/pNJI20im9BMnr3Rn19L9vS4m0csP10UIzSUR/
UlLj3M/hSRvqDnLsT8gKHTYrrHCy2FKgqe88SyezK1avmc90wAWMpaLs1gAMCvfRBmbJk7BPnlV+
bPZg5c4qbwxU5/k5MV2mbBFzX4G3jwrrgjWbrxUQfgmlWaPXVEtlKynsdtaQ8spBK6DPKC1m7CJI
FgfPoZVVvj8ZJOVZLOLCL41VkkzRbal3Y0Cf2VaFjpkxrAIXTCeZlPyGQC3qoD4ML0SNQD4XmYgk
qZJHneDVcTRoNNTA0qbSXUe2fDeJ468uSUr2i+aS9nuHP+ovxWZAZ9SYhYWyYehlZ55nyk28x1q0
FZnLfSHtIOtiBblT0GCQ0QgrAuHk2I6cRmJZ47RgQOeE7IEuAuB/YKXggtU9HehJF1EJQCqCbImS
8GAXE1+ThfC4IjyApuE6bWUsWXfF/xU4+hCceepZ+RAEHfejIjdWkzkQrJqm8I/7O73MIIRm9XTA
EH1iUwsJKt64N+Eof2YNoZox6YomKtMtcQSzOyP3LPAFq1olM2Few6NJF6KeeScgkrmvHerIE/tk
1r0hdTKOVhFHZRbb3OhfBbXnuo/UFgZqyapVdVZr+wUyf38CiYYv0aXthUer/OSn71jn9Ybjz7Sh
NnU4KWhjyp6L9eiwkxJENVMxUom45HD9c+a3BvZ0ZAd/V0EtJB2f6iiM3FIo8kyqUmJEIULepgjE
epbBIBw1glMyYSONFyA7L4lZG5+0l0oFanoMujfcJ3dtamkk7uX/fv3/HpkPuHQbd7FvkigQgqNV
Hcsbim6TffSlDOYCPCRQqYQW4t6sWNX00XVAnqTZ/pUuu/n0N4r7sGFw/HPMY3mxwbh2fGR+1mX6
fR4ovYUUCIR0wF3Gdl24MAHXyxbsIOyvDphy/Tv8Vbr2dpeSnw9nXdNwJioGBa2u5l3RhA1J7mGW
cxBhQLWCafxihctxXcRiluKRNg0De523Zopean4VNs/Bwci8r9PQvWEMlPsDRGmnJwfg96T2QNvx
jVJOn4uFzYCHhmDijAqL9aHp68+UyYdrPEFQfAmTf8bADm4Jq14vjsHi6jgipvtiwvMLILqQsjgp
0srqqxrV1v2wwNrogp2cQegS5RfwMIwARh7snMoNv2GGcpMw68VPji5uaPA0vrAjAdAAaEkiuaBM
NG/R8SmLZuXnVKLJpGjb9V1xarBDcIldLuVosEMhlktFZeOatQMzSd1o7ngLXCc5nC8p8fq4AK8M
SsUsAYqtFFd1n1D8AX+whhCi7QD/bj5bxbLwNfXvxJlYnLgllB7QoFwwZylsh00/FrMf0WnLEQXE
1dbxiji6tO8LkeyR6RMyfDgYFwwPSL1+6+WdFoksAPXPQ1HNkK9PtZDFBsenFHXX4i49A7wwkq+g
M21mxw5HwOgTv/XFh6z/AWQeKCbtzSL82iU3j4wNQp7Z+MBRyWsbKh3fwpmAZDxCkrx9/SOrpiBF
KXsQyxjyoRpFtDOU9QePsuzHrkPfyxCZVjqsHICSJHZdSn1OHax9IMslGfs4E/9qYJkSC209vT3T
J6oL4B0D63psJKW/DHQQdwHIUQ8eAT6/yjW74RV7wOkoChClQfUqFwgYFMEVfr3pulidYwZt8I7L
k1nQe51CUSWYvJGXIB3JCbDaQbMiNqptlLazWMb80JBVxZmHAV4joCCO6ArA/XoSaSpyVYG1xnSw
fAUh/sUUGxKKukaYO1PPZZq9ryAA+pjMwP+d5+EchBk6womBHNmORuZVUdIjV/qjDFMLQY43k6mH
+PflKaWQZk0BxMIE4WhK4mrGd4wN+jxbOrJEtf7dUPpsIziVrkrV4pw1eO7OGsvrT5b84Gq5M4t0
kiH0TWY2a00BaxW3HGx3bpm9FbqBKw5yvI217TnbovncxmebnORovKGUBnRmlV2HDGWpg+Jm61y4
SjoRTELDHrA5mco6NyiRU4PAqzXz2q4xZaVgNgzfc96287S7sWcC43leFHhGkUoJ129pp4EqEcac
rW8g8xkmcnFg8BBHoWLZhXAh/I4Nm/NY9pEJKE3xAlTkYHmBkDlRA3ZMOd6Rl8BGULTLGrNyaIAG
0xOivltO3VCvV+f8jxl17vhjdX3N5p3gPqPk+Ra6YttDJXHAcXVCuQUcJT1p3MB2zjsnXKY/RN0C
iHEfjvCtc8fqRYSFLmY09HqrXt9Hdu6AhdFOFXNd9c2LoYVodpD7WJKv9+JQQ1s51FMsvYuYHUCe
rUtVpFrAVQbpWCb+uNqVPL9s/mfLjuxZSFy80NioviTI6LpWjr2H8xVnxtNA9MuGftWTqaOGPznO
41YkB+wySi1Jz0OQ26PXJIDLYjYDaDmvrdIJ94uA81c7s6Z+y8sFjZ90Jd5iW3T8QBxN0WuIcwbt
Vgcq374HMwPck4BHJ0ov1cVn5OvYy+i+9SXdkotCBzQ/nBVgvs/7lsEHHQh5QbNaF+LATkC00mJy
Ku1uyVE/I43/Xw9q34iASRGHib4NXXN20VHwmVsOWMHcyVsJXm5rxz2mRRn9as3/Crf8t0PG90RC
bnhjm5A4mC1h6znhr1jaFQjHJoHkWoqL30fPQZMz3BbvNy7gAaIzVgSxYg5m4EALmhDLOeITiSZp
KiL5PFpJlSeySMp1F8H8Ho1Seqze0tmADgqKIaBd/jwjI9ZFJQppofiyb1/AyfGF3hxN3/tM7Qll
qQqW9i5KbH4grJQq49We9o4CNx0xaJOwy2ZRoOOhwXL+BHPnPnOCWfuTpw/Nqf7b5GVFzhltKiT4
gzvAbVhHAuRQwkFAkw6mwgOq8Bkt2BYdTn4SpCuL9XbUPbSG4gxnVp8iq1l1pmCYf7vzG+KNaL8m
YltkfsTaOGa1HQDEm3FdlPZmAickQrlp5E1rRiBoAlBx7YrNhRq/c8tdKBMOW5DIUFhH70OT3oeG
gKRUMLdnAbAEGVLoNJ3HUJ7mQm+ZJ8nTezMYgGQSSbfeH1uL1sjVk1oHYPfX/H33HankeJv6BRc6
n5Q+WMkEBLbjwcLPyogbh7kHnMQJ+cPCPURom0mX9TobOCosNQB5OcqScKTifn2+8DpIhuoMN37v
WuyPZ2YKQ0ZDLIhTmkAHwUgVtl45ChkF591dsrg6lMTvHPDoBfztXfyUe2L7MttYBZlc27Y1prx/
r3BNvlQ1MJH6tx0uVNr6kXNUHpw8aLYsFjO+5HcMI4c2N0nCdM4q9sdOflPQ6QnK+4P+INSteb79
SDVR2HAEA7Bhx34ecuc7si89ZPRN4t+EBgKUbUQSzWool5qPLkLCCBNT3b7IEhIkMeEFcXmbhC38
sIh++KA9xmhf6K+sUzcGDyRz1rqyAzrbHCf82ICCZdv1EFQQhrrInpseJY+wr/2rfZUUrh93wxws
OhG38VzbvU8TfrfSONGwgQzD5BZunU3393G9n+14WEBd6Z170x0sg5cA1Z+nspl5EO9EQdZ16d6z
nFlr78ycxOMi10brgLzApoOBrwqgFUoXnDqGhmeZptudxODqxd2y8WDQZRKJIJprO08NzpMu5R0P
JwLHK7xIQfj7qfkWh7Y08YhhfSpPUPJs04wJJNOC1ITF8y+zIGpnIQC2GRzUC8rRMH8LUGewgIIA
u28Njzzd9cRnaujubM3OPaHCR//E45wHaE4iw8aJlZ5BgY2ThZMWZ/j6yIfrP3fHGSh8y4mhvm9b
IGOBiNF15VaLaot8aYiixhvnl4qoPUOqz2bdAKbJJwB5swj95FzTO1jwL5EgjTaJQHxad6sr37Ww
MKgLFXrdI8dBm0TcboxQ5eYoHMcMsCvPd59QBgtSycn7ZuJ9b96XXZC+oPSNRP4t80ZVyfTwqBLg
78MEOMY0F3iegL0dpvI9wdDLf/iPjJeTqBaqRa+cCYe1c27oKIa/YZp4NC63IyOh6QwjPVITw+8A
Kog2iGTubjtW4nnYS8FJft8dI0U8x4NvjryQX2D8LLZz5n2RJqIBroatxpPN87qhPbRUhtzKzY9r
AYpNfeYLp225aU/zZt4dc880Lvj1qBueuOPrsXQnpyJI3AmLxGjymmMtDiumpRGymdsaFql/Npoi
YIqYVg2kJS6ZO13DcAdeI87CwaCN0ujGY8MDitsOgkyCsMYpnoiU0wCkK7DNJHqOK20H86jcNS6z
K1Fd1komacCYyqV2pzu+22tCPXNTrGUalX+wT5hKVEQNcxORfV7ibpqVG9oZzKKkxEjJaoypVFKp
DTe/9CQwHheiuCVdga5U3Sr24hSr+cu0j5p37P07E4NqNyAzVKsL6LqKkhZz2IpqGIfxLMa0luyC
KgIl0HCgxguPg20SoC8x8lHDj5bBTZMEGKJbO/Ets8Jz8PxOPToSwY3MYXHgtJe8btDIW7CZZYwW
fwuvzhQgaVbbFciofPJIHcfBtaWTVfUKXGULVbWuU4bB1k/GUAqPkJYklJrIscj3em10+bMGbcP4
H+ka2CJojtbfLPTFeVRSEhv8uxQ0ZZ84E9/QYVYVpZXai5s6J4T2kAMQ0n+0pRp6WR3eMX2HIaMF
rSZVjOZNdGRbszS/m3xmIQ1VyEpmd54AJLcZAyi8AX9YOmVyEVwV0sFsnr/9cnU8CS8lBsFrnI0T
28wwFF4YzgTN9FBFYDeAo9UpjrkWzeW30uTmyuuSTff/BBLgLCB/QHDpuLGmw3J9H57t1B22Idi1
a4Rk2IhOGfahTn1/HbCbOIqLw/C/9wyguGmE3K/7aOrTcUEENP2DGz7xTsQT8jAMYgkhJk/uFWLC
LZz/++Ux+hcxFxvEXKglMlny6l6I8wy/HfHjxkgOuGuxh8534n1iXim3kdw1Zz0cZA0cVsddQM+S
EW6sqOCAbHGgxEa3lHr9VIYJb3caciGYhk58vKIMlb0BEV7akrkuEy63BvqsjJ2JZyGYkgZVzDws
KWR2kf4d1bEQjtpIY6LtmbdRuSUGU1Wv4JqOvnHAxpqf0Xw0TK4CWqCkcN571Ld8mSVb32qvocmx
2UFDoEhwTfbPJy4dtiDKtWfm7ERr/yoUmwknN8vh7w1y3p0fkt1+96swfSRFZPRu+2yeCYKTALhY
BM1ZyBgy/dlv3D+4UhxCQDODDEFYgqtmEoTigpkf5MxUa47aVclSXGvaCuYInLvFyk1LHaPTfIJ4
P4rwqe90OiRX7qlzxJKUy8EFnWIgxsymBC/Sq1YZfA0aI2LqTieRUXfxdKzyNdrOc1+vrsbwV213
ghgyLinRW88S8wx57mZ3WUhkLaSr3TbrsR4r/mZDqziZvLmwG0Y8M49aiNZ8EQpSbdnGhDZq7cen
5YKpC8yP367iPa6SZ3FybohKx6dGqY4anAhLCRjTpqSIJVZcjmahI7uJJaiQJAjrsytnyUwBCHr+
elcosQ5IDAkmA/nItSnRUcublwUpBInHXnnecac7zKDp0VmvoG6QnSWfcpHId5qQo3zqZTrHouJt
cnmxCS9TJOwL5wIC48C9F+GBy/1eJ/2KJ5VHBxPVboMH694d1z//2QD4nuJ6cO73+hBnDnFoBwve
Y6OKL4/SmPKuGiMi7+AkRGKUW4S2DUm53MaN3x7WVAvlkND6fZs+DsavciyBFSwbiYpXuFvDg8Sk
ZeBBST+x0nWskwvGVuhk3Qck+c5mVYBpUfCpbz28WTTatWursZI4DwTLsirHaBaDlPJXqrZc9JxV
wmR1urqiHrpvPqYwSXemAhuUFUNhx3udIt+ritMqJjUcbCf27aYVyuMzEOJj2HvpOQ11jUhgX/rV
nG1RSCR7G0ZcEvIVUvqT7s6T1kEax30bl1vJtQVFQys52eyXg72jx0QujZZ1uIBlbuzJeuzwohMQ
5MI//eLfe2ZjvM797V87O3xJjDcv5HFhA7AjmjbyWSsN/rmBE3R/2WU10ZCVznohlsulqKF5DU2G
zMpt4IjJIYN2oXF7FzKYDe+U2t2n158Po4Jwe0FhTQfLA0XHoC7Wo69g+BZoKb8GHcZS8GRRw/dd
u0CPVWpABfLpulP8g1WSK0mkAEYBfvBFcbhX8Q/abgUafV5gl1/4/HeddRl0MKXp4UkHHnc2SJcZ
Nnjf2RXKvW0jjUGSZAl+toSCa8T8owyJh8CjXoSwb2SAzylAOLe+UijD7PyRUULgMv+vuWE93Vl0
zfeNeC5d68adkJyDwXK/uVCkgDwFT1vKAsDzsrZimfpWl+A8o/Tc/lJHBJUoAabZYc+wJTKgW2sh
1IDAqXeqYGczfvP2JrVRPCTvgiikZIrR9V9XFQYiqWa7QBsxKmAOIsPnhpJhWiXKTswXhjRywTK+
bgfX7dRDDwpRLd4Sv8EcEmtFV3t5lcldd8ZGoUXvvleyLwoMugZ9mioKL2yBr9TqdxVm7A4xep3X
QmBHHaJMXJtv/zLGDZEpvWrg+XoKRu/OFwE24mD2002w7m2yHsV8Q5OWQjzJwfLPYEV1Vcvf4bXE
BLc1+DSHGmsRY7sCyyDlcgTBMv+NdJXgE3d33KATQDio4CROzO373aYs/8CmGacOoEFOy9K6/DEi
KyzumgaT1V2VVVyXnLNtYFJ5xqX635GNxRxkCbc0VASojNzoY6HQ7/ON0ZsWcL4wAV+5nnSCudYb
QUIng53K5nFKegklI4wYSGvKMVvmqjuxF/JohZF1Qx78F02+k69pgQJVVcrMFTX1ZTqU9bB4HV/H
qVCVhSWFfZUcbtj7xJMhnZsGah5Js/64QIkxQLtcnDmkCxxHRF4o6LgcQYEvgcXfs4c56gtt+HlU
NH1aYDt9HtTyMSpE5+d325CWDyz3CqJZO81lX9ryUgJVBvOFbNShurhKIszfeGoXlGARy8fAY/eH
md39UXi3ebH2sm/bmjMsKChNwI8riDT8TkBzUMdiZ9OBI9lerYhtdeTUHhD1PsNF4n1GVo7An4Ob
iYZs4v2lo/n28yRt5l5Ps/nH3HRemsNp7JjKKa23BEhL/yDmy7Cb3/RZWXRHRMsql/96RTcgOwZB
AexIBzFXZf8sua8+v7qVSSYAnlpM5xXmvrdIsXDuiAllX4ZBlbLGCf4zGEN+kPQnammNs2PN50kC
nssT7NIManPJO79UkfelUvT5IFis5KVcMlh37haULdwJ+AetcfQ0tomkHZSiwe19jaxE3V/z6umc
kQLMKLsEDO2YNySzrkho0hb0Y8E9svZN2fCMcYTvqX0CEiR/IdwbQYXiZmiltCI0kQNUAyI6LBTi
P0csLdcDLokMzrGBaGkerGXPUOZmLMyhwfVS08zjY78jhRm753aDUcPWTNeOrCfnHb7y8/pq1Wqp
NsghcJL3o2VO2TIK3RAuKXsy980zOgqTMtyqlzpQ8mZqhZ0iR2fNrOp2she43fkgQV4Qm3JKqGrW
iUtcIRIr4rCxhwdMv6wZFV87sF4ZCuvqYaZud7u9q30/l9rI0WCCT2hNvsFrSeqOsaGmhXg7jTi5
qISsQ0OpYH9x2pkR6GAlCcb7G6xxxErMenIQsu6/GfC719B3HCcuaaDvuWzmpLQu/xFXZ/SuKAus
s9qPfdmWmvHg0NweQcyUGv73p8Png6p8A58okBDGcZLfJmqQzjTHbWlX9CUK1+2h4dtBr1aiSiiP
2rlc1Z3944TIG50AFCD2T1tjyg7IfgG7g7Dksqi4d8bP9Ix0Sq5G/omxdEe+0w25V4HYui3RNXaH
4up+rx/BEozhtwKYUZqtwTndehhdc0ux+9lL9fOpvIKDCgqMBHIcklcEBmFyP4TNo8kZr8fNEVQ0
gpBrn1bk4vKeeGbccN81fJ7+Ap1pycs5nttjIx64nCU0qYbXgg6PcqPUblC1jMhb+72hxbvXOfby
HEo0sVM7MIoopv7o7F/7hEJjuxtAQ7ulXWb/OVsMX7rg+QsgJgQJ/9idi7L5uztULXCDdhWlRFUq
oCPy94wmNGknr1gE348py/YSZLppajd6AguPmpMO5LSqkTQEPHkoeCSXPTwbDuQjbisuadYLOpQG
lwn/L8ZywRWs0x25sdIMhU/8euMPDObnXBRadafWbd8Swhpr7uooWG9hVB5KytV0NfsUHsbiuxKq
M7oOtlTnnoPdbIee0Y4wMIue5dG+uloZzWuE0/dKijbjoIORJ6SKvgz0Xqgqsc8/NM/S2YtgHe4r
PmlmTchPLG/QZoPz/6zTXqpcVn2UPyQRX4w8msw5V7xqBcxnZKbYFjPKKMfY6pxPFQLCpF1ncEJF
T0Mw+4WYFaMM4gb1jDAd+p9ar9RiqsZU2asmP5kNthlqjEec5c5ftCTVMg/3sqRfjsKMU5Ux18fQ
92izwN3EzR7mDZpP7GNVEKZAezgZgLgAYugeJd7ZBvM+YjW1cjbBUEXcWWRzNaXImPiArd5rqIMb
64EmFRjcF1G75JI1UjWiSETpGBpfkmxRzgqElQZBihL5W4ekpmOG9AurhNXfgR+hXI0jtDPnDxJL
no7PVYfzvIF+hM3r9SE4gnQQetTTiF4CVFSZ9ZKVWs2ZmKvtACDUExU0umMU2igFks5XBo1a6Q3o
k9bSQXqqobpsIDzyAzRjSmL1bgtRiC0FKgTg/dPiIWoppPuP8jAb+Oa9/xLBFJkKVUml228ZGpig
MVygEFvRj/VWa0EPfuy8MiRS6tgrehbzo6s8+W0D9k6ERqt4JRtIVrfT1CcRLbYhuNWMzPEo5tV4
B8kMPqHklLYRYkQf5H892xfNN+T6JpFdbynOsSGdOUVcdQrGa+1dvnV861UkCfZmhxICkedAZPPR
ODolnfhmh6ARGb7KrGg9xq07KRW9g/8gayOwpiWoysGkaGoGMzWCRC6WeitRvI4G9JONbBCUUh6U
dPeoaZS9J4DF2VXS2dM4w7oFE3ziRKIk/YMoXm4jHKXEQsKyf/kxCi1QShKoZX5ftZE7ayEeD+Be
yKSSplqiZpvbq4DlZcvlN8ouFjT5qdtQFjZg1+YbuisKnTUO27K5qkjJ6LpIlwhyfgrqp7KfHPZF
ez9tyoM51svGj9RQ8i5xuJz8Qz+DqXfbx+eJmw1TNna0RzgPEKiMAQzegycrcseIbagkvw+rUbUB
290ob10cyVOIhW4bt7z7bDAb5zo5Hsqh7iysumtCwcWz2DO0NZxI25JFjLQ5m50/nqYuPmp7VRsD
4PeTFjOUUJII39DS0EK+AELTkhUb0ItiTkgguFBQfANQ3HFFc62RrmWcVNaysqbAb9I0lU2FGB9s
5drwHIknzz6Z/YCZRXguXLe7YFqp0/DEQM+MtCxaXV3RRsraYwETI7J/+F+KQv0GlBq19LqFO62a
Pjc4A5uW2vRhsxus+9di4GJvHxwZ7/zmpDXz5bBzcGQvFyU6laB7uzU7stSa1qXkkgOzLuC9NShZ
b0GeMX1GZ5zOxXTxvRuWC0/RjSZnnyFChkIaZ3s8JdPpa1N9cIEDeHXFIPfOsj3/qhseNVUBH7oA
/27T7IU261Klg9ohahLqe/k/fP0ZY0hUL4ibOPOFYKZ9duoeRT6ITzlX6HIa0Xlb1h/SIF+USeQx
XfJehV30Kk5iJDeAKkcc/SVQyLw1PtXyZl/Aab3jKyFE20e54y+tVpKntdBmSwTxq9hqoImqCf6S
5Fa1uzp3tFNxF0k52C/9Tsz75uqyu0yir9u5RYmgUEOIqF62fsyTbViqkpjvjZUTDMr1ktma0IJA
G9DHkjnchwFj/rDcSdkzkyeRtwzrX7nxVBSE/3R0DQzke9E75CWKAbeytiXFwz75b0pBf6jb97I8
UDK60xpCc5RUl5AP6+hh5e/YCEezcnvlFDbwhQfB+OSZRKiNhWXvQeL/1QLbkCxKwhRn0VsmD2AQ
fmq2fxIYsu4qiKbaPD/zd4NzW4aTubeyY23ZfoLIL1CN+INcfM1Lza2kDpqnE40RUVgbk/kujlne
E4MWGQ9ufAh0WpvjdaG/vzIPXjm4cjPtIKnBoblHPxQD0q5N9ycEKsXWJrDOg8s9QJqMO/JcKo6n
qEtIaEfPy4HLrYphMAsBE5k5G+h24boOEfmbzPT6ckpZMeK0IQ9p6nrVxunG9WUb2KUPfP2d533m
pO6ARJgCxguIXRiXZqy74XhZQ5dEx0fZ1NiUbCh0YiaKY4A6AfAc78z3Gpxa9GGNhGXmuX8TAIpX
kqQ77x99c7HiwHiDgyuMIb324hCmsHoCy32ZZLGyTrLVZjF95yFT5dlA4PqQA8jYGLVIkxBv9axv
voQjJMp+xIp7iABFjcRG/3R0P8URBu7I6omrNupb98URBBq5TlUAHpUllY8hqvzJ88o9B9L4Rchz
SDQqlVMU9a5n8/VK4cp+vNUm9g91fcWPnB5DiqmgWdEySKbTPnOZTqYhsqpfxAAEn43IULXeKtun
QZYB1UAXvokJR2n8k5Ox8vDsFx6PWWu80xg4aGgxJz0yQcqyFoFOZW6sBrR0cso9ScCgiwlQA9oF
3zjsZ9cPT2hg7odJfCreib6j0ec0FcV6KK5Iu0fwznq87eJ3F0D2mJG4nT6lM02KY2HoOKJ0fjOy
p1l0CA3GpGlvs8xNM5zRMb+VAHm16Mh7Qe3WF8nibq8Qr1Jp9FOzup2eyZ3AoDvbGpjZQSbsA/OR
2nvrIf/0uIariYAgFsTp/hrvPWCTNtBrgbPsTrzD7pXEDbbysdNRKk/spWyCEL/sOsBPJuhsvfEh
WZullm0S1haHgPxWFsU3fXX44tWXqEYp0UEWZDXWcGb0YFDQC4j5YmdDUJWayDP+TMNabVO2D6Mp
1JvrPww3x4BhPmAkNEuFN94i14jUXgpuzp0rNXg13AMCJNCP2wZEierPH60zKpD6iRCXGtp8SEf+
2vJ51Jqy8qbAADi0K5g2sHi+z14aFr0F3qsut3IZMgu7R34XgGQoAeBv+z4QOqWWY1HujaNXfwN2
TzjWVfPDY3FQpcE16LjtvSGvlnWS7gxF3u29E5rkVR3l2D/lj+IH40uhxMUTogYXzEj0kAiy4j4i
1jZTM5dK7LZbc123Q1AMIhR6yKuzRsNhSz/UOCeK7qAFx13ixNAzyPdig2ERHp3QG1W1u0fVApBS
OBHBGJLokk26aSMFXTfQmf21MgVJcg1PgrAQh5tQi4qdzlk7D1BAGckG73tI/2LmW+rNl3M0WfOD
NkNIzdGoII53hURVUujZs2UEH9AbB/F8fxVcmhsUNcQH6hcddN4lTsoRPjOn97lKKT9MpOnr4gix
FV86SOZjS1wnxl7SZ52EVUw0+aBaJEiz9Cn2ppw8FHeYhC+BioDoTiNO1AASNRyoSm3UUjsJBeZs
MuiStabMeAd+ZBo0N+scaXjSVBzs50z0deUfF335b3G2eIWAWHrH074kANKO4BH6UyD2vBKw2tS1
JVlR1XvfQbdlwlwNbue1BLfCPRzJliERsDkksBK6mdStq4B5wVvFm+4+7lFQGKGbJaWek0wG81mN
SDZSnx7bMK0k9Ol5fueMZ9o5vvPznbVVXRRs97zHpmeQsR2bEM8kG9ObbotPgdCZTTOZKX5w9Qjl
p52ns1S8hh03YtuT3hG2eYVU7HNT3k11VNKS3YBQeOpXjK6ZgPUpwC6J4j5KQqeT+oo+Vm4K2OTn
XaxM03q6hNYHRw3dxeFzVgzPnT3aXUaFj6Xrz8TP3TkMTX+I+39C+s+734kR1zZoF5nas8RWMM65
iZbDaD7YIhCLGDdqsFJSvzL1+lQretL8X2PHC5XFov/vq4AjJcbJVgcMy5obSGCcCk+C2Qgtok8c
7MK65dIL4rPpFgxJtkuGe/VzwOrZJc4rjsj0DTzFCHjqU9+EzzUmt3AARY36yzIYHJ1aZb8wbEGz
YmhgtpYdZV+dFEF7fxWMDYz215yzA0LU3RjDLHE7MVzNH3akBGWIKfsTP1+AUKxjEss9XU99XCqW
wNe+HE2E3SLY7BwzIYA75nLQyTmHn6bLBe2fFvnPau/tT0Xom9h4vmCcZNd8+5vCjtMHX6qicju8
q/DtYpQruroFkzremhKcJeQc+7U22dYm0IdMEP3ZBKXsIAyzWfYCfSGfcI0/rj9J6rR3e7pWijpH
TmwPNEpd/BRny27DYPSg8ZTEEjOXZFOuXlvf/Vo3hmlZhDjYGNWplZikfMKNHQtqMHJIMBp4G81Q
r7hLu2tAhpbSekiyYzAeT+YmTg0nn7N/ezfHk5KdPKvv6x/50TNPgNKRNDH1JknCjx/ANDdCiv/L
FQnBE120MF/59nEnXu284ppzJDio4hD25GFuPFBEc5WpjUFYqKY6Pyp9CDmQcT+QWTP0wdnrbts2
//QubuKbDbqJTJyv1da9fVdMTVfxJnEIrAzVB3Z+sZKQLPaV9M1lKKnp5Xp/UVtGi8BTIx4pUkJ4
5Y/Zbs7RxxHe3lAgzKseArEfYzUlf8qzWLqufERlqhL4XMuqvdEwcxeyQRbK8nosAqu6X3Hq4/Qi
biqA+GrVg6KGTL7+QUWBug9f+IvLvseJw1i8mV5QfGfyqAOj0CkzR+D1e5TFhZ2j/kdOuKgKzGhQ
Ku3PMQUAbt1KaChBg+bQ8NbcVtwu+v9UEuJyiIF3g+dD/poO4heneFBABeT5tLV/q9azkHvTiYt8
kIxbmXkDhrjwUIOaDqn5YMre4eA0iUBo/CHMmneuqmrjAQQgb0FnDOGJDcItpvYOYPiS2qodADTn
ueD0PWGjRIchWSqBIssaIVJXvK9zuL9AHYcHBMMQtkqfeQuuMnDkhOEoa2GN7LHnPNWaKg6Lutql
0/ivI1UYqVyNehwYDuMXbq/MH8U55PvMGEHDga5F+tnbRPt67MNs1eolc3RNzantCcK6j13zs3+7
JLoi8e0Z4SXPqxQ/USeR0UzJX+9lA4ne1MWCjhF0aKbk6Xq/EMIZCQhlFbFxrUtFIMIq1ZCzKSvJ
Sj/lLxWwh85LB3aev7xRhjJOVVpp+d9MIsB4jC8nERmM+dUwwM/uf4gy3GewOTcjFgYcvEVU/yea
Bp0i/HbNBr7YN8Ef15q7bewi3d7Pu9g+nQEQA3l2wYpHGEOX4rBtDDHxh8e3Sbq9QwGlVrJU9khv
1Ep048gRv5KoqHZuFmI2H88bUHvPA0SLvGObiykNLndc6YvCG/hfZIupiDmUakuBFHcHMuHxmu8s
uceFrPLmvugoQMc7eolTO0BvhCUsDQ6JgdGq0x6afCdoQ9meIIVMXeSVPWBDFwB8wuLSn9iY/JoM
W6ulqw03+NFS7eF8epglUjoA0+pBVvdcxlzX0dPov0D8MpxwLeuuj5F66INHHq0Mxdv3lUcrknVl
Oe2o5s/Y/nh3iVhP4rKbow793LzMDV6l+R4a84a4My2UsnjylL5Lx4WUgybK8DNYdkXtTN/c8Jvh
eiKm3H6NUXDbX1myrSLNWxBfe562/ByKlwTcrCvFNIK6pkZ6BMaFmXRi3rJrMFff1NeAODCejDRh
WRetv5z4c55fpolo6aR14+ZnfJakmPkO8DHi6KSO7D0G4ni2QiIsUZ8Id3SAOuObnmR3Yj63vE5l
OjwopRJu8lBwcZITWzmbPgjE+hZhUjnZKJSmBuW5+lyBYvSw7Qj4sQ3BNWa6UkaBeiw1wg/RLJhT
UwsLNTHI+FZe8pXWM7jCmzvNaKMqJlw3qsXG3bi4U3uJ0c1HCqBZh4mviA8kpbVQBbNCJy7e2AYz
yFt1REIFglz3q9OH6CdXaDzyMHhrmppxwJ9xQ4Bu3eRdR28Dc2z3qfgLMzw2pOXmTHXNG7ApQ0yJ
f9KGe3VQLoMbWuP7tfwfyrGUEAMcK/L17y89R8RZZe/2JykUA3Z7QiH6c9EBEDGedCF4kxwJm65q
hKUi8hTNW4JHvHO0Ab+gfgBUM+58dXsU59ArLTZuvS6wGoRFuGWC3LFf5fBBLdlPNCcInN9DVDiK
aElmVQ6fGYb7ZM+ftCxy+GLxselpXEI66YxH4N2z2lxl6Wlk9g0zxw7WSerwPlQR7a3g+xkeh8+G
zvsSshm5OBTfAELguyAyg40K0ZVVTjeShyzGdq8ML3GUghUTI8lVhaMs5Evg6HIzTJW7nx3yRVfK
lkSJ21ZCs/8ICAteW9rCRiMY8LeuNtVAn7p+dzzwtToHNuvwAF8BuIm9smGA/exRsweQnw0PPpri
CHPJ269Y6Qk5/P7/OZNwoMeNRherCUoYG9QeETRqxiXKQgAA4qE4auDwGxxmjW+zhxZJaeIXeI38
OQOAYCvtu+hKC0bREz23ip/IiR49caHVJUEteRjZFhv0ncJeoojb/UKxe3rNPrmG0ZPl4FfHC/DQ
0c8854SjfMxDYXIlzXvNcx8hNqed7Esx8oIXNVQ+ZCnJVlZWD76gz5cZDOEVcnlIBIivJ5SZ8DVF
aMzve0zcPoqhSOlMbvA5rlltuDqCKOz2mKq2HI+0kcfj3aix6YzlgGXDWAVK+2fqxK7yiy3tCAUD
5a1hA90IBA2PERH6VUjzxrXw3rSno3l5sUJ3voImSjq99PUGbUNDvbCl99l7GJjkEetTwyvdMWBJ
2UVRaDPXMzh0CwMbnGo3/8+OGhHEXPQzdCA2a/WyfyfByIgM2IosZzWYgiKj8b46sspRoJdMVOwZ
fj6O85luGcNBfMvd4bdVYSxchZVzeSAgSo35CkgHp10MFNjT4YLXMD5NB8WUGDtXucS0YG08Dgpg
fksVcmZ4jzTrrEmBmAyPTNnSBB/8APBJVXLzJerHIM2mbh5MBhOca+dHMAW3jEZDM646LLwdO2Fa
TouYAN/nWYHbUQ8vcHOHG/mw5K4kmtSIljVW4MJcjWRszb4fNzYDxMdqfDij9N2/zSebr6iTa1mi
3tGgA9a4t8kChvnhKU2aqRJ5SATJnwDMffgFtEbcFX6bvqNO01oWZN3S3xSq/KtfxKaTa4Yaa5ZE
7Bho6YFzDJmZ1K80Nxvc9RVNH1S4jb3uh1e7tJDtRfgOxo9U49W5TzQtURMPeoZq6z2EaeJU++LX
TfNtvY7QXd6EjwE0gdu8f25weOgOFKeAoil0D7G5vIKy+Ux97VYlXRgzSsedmbj2hsxdfO0pToph
YOx+jVMK5wtWb48X5ouKbXliwYAKDvvEqtEHO0uIx930cEG+5A/SiBR+2pTpTZyUW1RNneMEke/D
wGqDStEZSZH5tIBcGsvpktmzzsC5w3v8hLnbNtFbB4w+xYc5AQk7z0OTs4yZJ1rn1cGfvVv/8abU
J664VadtwHXmyyX/lp1WLfW4aKkg2mHXdowsToJrCjKpBNP73ujfYvubBnbXCu+F0Of753iw91Im
K56VcSLokqphs2sWSU1taaC4Bf/UOmXM9PG37WEO5+QT5cTV3MQkHO66hfN+klP4ETy1ffJ4DKq7
Q9BlaoXSEKGiVqrJ5/TkAtsJ4DbNpOP43WKQcCh4+c+pbfIIq4yK0/3gWvSpjNQ8r201CNiwRZI9
xLgjtxY+1LnuLGssvLuTii2ui4MUfW0A3MHl6GDKT/FSrvqyhzDjRR90BKOxFF1xq7xC+0I7O2jB
rWQUcBUAEBS4tXa4jRDhAPSIRVdxW+2MK3H6a9Rkw1u0n6a5u4jei/NavcBBtftp42yqzZaJuyGo
8f/O62W/y5iK8FTIJCdvEowfavAGypJV0Ki/B+VDBfpzheFgACKiLIirloAV8a9eQHBVCnTc7X6t
Gzf1Okk1KS8BRuqL7LBbHaAYAQDqqeOEqXKrQ8PHmqKy5lEDqKhAuytABz04kQ38a7hr18VekeID
oQSaEnAXQSK5mj7HroJqByTR3RxYUx0QRHwpgMj8KdP+DB5hHcwsnm/a7tftfMuSQOk7qeLjP7Ss
iyiyYx5S3CiBvAQ6cwlz/J1NKpF2kp1iRc2nqBSsAdXbYUvsOifNnj12P9aASUM7Q7anYW+61cHp
9kkHIiMLNDPdlvnxRXmNlhdgaQRiRmNLHJ2saLvRyf6gvVVsbdSOeHYxkCFAJMKfjMrukoGjdoIi
sII3Hpa2uFPE1UvVqNz8uzgOd7D+hyTfLfZlMhG6qsncQeRWtqDMnKK9k/hrvBz5Uooi6OLuN10h
4QYMOUreGWM7oMNayaJjQuXATbeb232PTxOzeIqPKZEGCQeq7G/vXxgKlyjJ5D3SFxJNHGavjmZ/
QSp1HhyoK9AQYHPgb588mbkDKkY+u+Qrb0WAubvP38SxjQZf2HwrxuRJNscEAySK0CP9LMt522Hr
L3QLpId6VZjKdu+7pvm7Y8P0JeKt/vIvDFeC7Dem6KuumGg+VY5a2amY7KrllkrVcLIZmqwz9+R/
YVaZbug+pNCOEP4GG9TBu7AK80L3PMtI1+HE7T73ERv2SJkXmMRJhP2g8WJG0rCmXibMrbVm6qW2
Vqj/KDsGFT6hsqY53gE6bisH/Q4K8dMBv3vq4jcKerVcod6xnnkW3/0cicgG/ZlnFP5dQ4pI9+VB
0kQBz5GaYDPQMGUlc5Tumr4x8QKBAZFbTGgRVmbj4KPYoHrjvAoBVlwCbfOrbGeeqKrwQhUqX4sJ
fTKElZU2EbabkHDUZyTqrVY6W8cZsjfWUIHq+bXbZwSo6pfavydghqOhnv35uQCsKXHocEzxzo0D
AGHuX0mrvCJcciH+Ifw3hs+rqwe7/QZFGeprtlAQE7P9/RT0JHRwjArckEWXsrqPyRip+GdEqbTO
R2VlUFaBBYyLPYVDQK7+Av+rB3wAb1dLKJnZ5L1xAQwLNCjfJXITRypgcFPM7SZOIlUlgo22KNHD
7a12b97WEXxFwbmWoRdlAoY7TNXWY1n5kCg+HR8wUc5oing/Mlzk9GH3C0WI9H+4YY9ka5mWN1zg
2o3nQG8/Epa1i35e45I7SzYa9dOT4Xjd+VG8ZGlkFTFRINFWzxcqFXMIHj48buws72OBWCoEebhY
BjwnMXMl8NjlVJfqdNmREvQZGcp9k/n4TNAd60UtRJ3bowIyNPfYdkwDlzdcFCK+cok9JuSJ4Cgo
DLpBhwL8zl5RJvv/OlZeESeAEQAB9RZdbo0KHtt7Ttupw9HxMRLOaYFpQ6gYolBuR/ChK/qA3n4X
kiG8PS0ro5/ILjUOFTE/EE59p3cBSPFT7Y/5WDEwqufk9IoFJUUTgLQdmpMyDpxAiC/yTETc1tSa
fLOxuD0RIY8SIA4RvNvkNbKk8AD6X7CUbMJRYmwicQ0zE9Jnt2C3UXxngpAgXa+KZYXnofiTL3GY
BScN/AIuPJKfvSQ50WhnGsSnSv2CkC4E+H54ZzrsmQBXwuRV5oNvXVXWO0LDZ30e5cv9ZQ+3BnjW
pxSquSwIS1y8PdCoS8LxYPaokonDDiy+F/UR4jEGwAZnNWDqwNa0OPn+/eCkVcNVBKb1q1kOeLAS
cobWbqmZCCCrETqV7FbeZKOeE5zjOP7teGGULZc0+7mxH4h6nLdPuE6C7Vg4R4rjwr953hbYrcsy
zENhIEu5gSIa1lXSXjMpqLZp719fr3AmuK1xGu6OB3s2MDkaZdwt3S2j83N/wl3rt7bi7Bh+kukQ
09+2alyV6llV0IBtQXmOsEuMNeSz+jCsmmqta/n/ciS3RUO3JCCx4ZLqrpuc583CEooz+yyhNqPM
tJy1Xv9rDQp2kmaNRCv72NipNJgKUEu5FZWGmibLcGRuvYBWyRiq2+JGy8LiKJ8t2tfE+P0QacWv
MCIk1QUjpszGdaUyIfTR6kGdz2dMOjKG/lukVjfsWJ6sUbJwCVoT8rXec8o9kNcFKoSatMFdn10X
0TtGNmw96W2+cJBZM+uYtU7o504kgchm48a9c/gLCQHApG9Yk2rfKcCCtey+1VllXl7D4yxNjVvy
u3iSnnMgeSLZ7ck6qC5nlsgWTk8y4FAFqzq14Yhq/wze0QO5lwaLHxL9S0IVxM4nx8LIUJdzJGM/
5qgh4uqqd0EreIWHU0SDQnS3XiT9pAO/KhiKKJMUWCWd/yrqyRJI5Qht3/FNrvYcn+HPMMOQhaSL
OXKanaFZkM/bzg1qjL4sMNkMppv1jC687WHSKFp9Hwjr3MXNnNercmulTPD41GXcxEDrkwQE+QD3
HfEeAcsNVzI80akvZWDnd8K1JcBuDPAGeSVcae9vWmaO/qbwG9dlJA9layp68pNtaNbbYKJ1P0No
hnJWQ8G6v8SOAanUJqJK+u2/NtbT43XNsMsNsDAlb1oc0D5lv6HJ+EUp0D5MgKYNeiHc1J/osflI
Gqi/xAF7FwRoHAnikChaafsM2h8WMOh1ozNJliHCAI/cZa4hqxlAa/FSYjt4wmipT43fj2/kI7lq
KLQQ9fVZ8c9wtEwO8G+JRqQf8tT+rb7QW1fqNAzjErEMCcnlThLvS8Si74GoDILAaTY1/x3ZT3Ze
GR0FB6hCouD+tne7OeE3+TNTEV/9E3YNkaCIs/iAS1oCYs2NwEEKRdBhMAhJDY9URPF/Bi/rnycv
67+tQMHpFllwqHfpQlQuAJKDkkjexU1Kswkt2NHnJcUA3cMP89YDkKcTwCAFDFHWOeFt2XBd2BNo
Nts7ypEqlPIaMm4KapZa2BZtiHneCsfKTm2JFvld5RjK2N2UPNF4gLJJArxiPJ1Fy9fo+eXif/Kx
dOC9GRoJsBSCxRbgCg1jLA1mRvM6qoodg6SBUWQtLEvG+HOnPPOCdhTsmC0YtJLM+tiZjKuvxBip
tp0M82cVYgLYNvmlzjoQ3v9wFoZHLyuMheDK4y3cvXYj0vkqaIbyqWSe5b2QO/qHB3GstFD/+0jD
oJPkGXjGUebVWm69Fl4binbq4y0aImCxfvAkJXOiC6GRHhl3cKUfZQH+6iom85b17upvPeqHMSSg
O4pPiI1VIXTy0eMNKeANBMM0rZUBwFQaUxNQvfZmqZxKs0RkcEoBUmi9B/1yiTF5dqoIsNr3p4Bz
shxRLulu7Z+roGw3Pv5vVWv3S+teyyQkuB1eKC04LNE4012CCxeh+qnA+WTJcX7iBRtjvrD4KLc2
XKns1VKKzwXsdlgTquVNkzvRPUZux1U26GQrRotqC1v7BVqTRansTtYs0PLpSxxEEAfHvKzIUlgy
KPwqjCGPc6kls6kwbq62TfB4XL7tMwv61zaQUi8e9okTttxQ1wNHZgqNWEloxT80Ojb63rHZjN+f
xzJECqM9TJhJKj4xLAPIPEnFm2pfU5EkSMiSiqWdA1+tegjffpAKepyBuHdLR1/P1soblGZZVjcH
w7CWrSDtPxUSHYfdLn/mO8OF0BGO66kCG1CwFU8jAg/SotrTp+mOWWhAOrnEBfa/UTQXGGkrXGo+
kh4a5We+zqnzldSrVugnipOUhpDswCNSxpveDQC/2prXvbeaeei2WgY8ImDByOKimuiXYagUn93P
dETn2TvLcm0DZrugv8KoM0zBDl522BgtlPu0pgt8fda6k8+6HKRkTuzNRU2gIe+V/hd7aFBNIxbj
NkuLAcebfApLXGOUXP9GijWY1iYUxJ1W4a7pkMNypV48idXJzn7NwI3HwIbM9MCL46Yu8K+zKVN+
+HU8yeYNDSjgQQb27X12NOz/xvvmD7rSQBysPjaG/CDV8SJGQPtD1QiyB29htmE7qzpDfBvP4bhT
ysfkLMZbURIF28kr2uV8OT9Xdr3MLBLK8FpF2e2A1Sw0b4aBrDn/7HGPErEW6maVkqU0CLZph8/A
T3lHUhkEjJwOt+kDQTt2FPvIewVBv1zINJcvItRKpzeK0DAnOJohS2ilS8jj4xHBqAdUyETDBXF1
AEtm05Ha2cfpTo15NqraFkb/I8zz74Ww1FYk/wkHBj4FPGNDXT/OBrmQ0bP4nx+Ff1KrS60yMHDn
dwHQ2VTuEAAAQ6z23UOLvp15ziz3tvw+xHPJJVPE95hNFbOsmB0J5wQphUw2dUPi/9fmND38qAMg
kKnW0MI1Pe8fzcaYAVLgwY7JMF4uXZ4CdpRP8trDTJdp3s+SY6qgak5KbBegRPSy3hwESzkzyvwJ
JxXmCok8BazkbHeyqzS8PYB5hdFBnwqe43a6dst/iIi9KU/CvWNYjM6pKAdVh21ueG71I7qW/tiW
XJwA4Hqk909jPwdysokeioH44JsaHf+FObhWrk3kxHT055djERqwwbOr3jHHLwA03jgbCJBbKRRO
oqCwGwR5xa9HGDYPqo8x7pOh5V4KrV89GqNE0Ytk/qoOIHgfxLY9wJi1Z6Dhwldx/DEx+QSvD1UI
D2BfgvfdHY4bI6HhUYm80d2Plt4GX4auJantWu5sBnMdQAf3qQg6abHDeG286dlLS9d7jPuNS05o
vyTX7/meozdskDHjHj/AOUyUfzpXUZ5IACnkEcKR+6g3LoRSKgmFTk8gFkMZqx+T6nZ0XiI+2gMa
wKIBWt/wK11F9vRsmMwySy1OJ5dASsM5qFZZI9dqlEOne3YTGQup5tsodWguPIPyuMlHtdnSawZ/
Xh2gZfTg8FzSHimBarbQvydABeYKvJr2oCS4rxwL7wZkMjsp96U6RqStePoTTk2CRcGWwdxntvIm
jvV8V1hhRTRCwOVSIBM+arD6t4d93pIEjF/hxSB1AgJWXrqWYr9/1gRlSS/KnA1ertnK2h7xaOsf
mLQLw/w1BMBm2FsNr0iMGGQY+HX8aohZK3mMepQpJZKg25fdqTY46FMwR853hbOG42QPhcBCF7/B
9vXh7kn62VPX5G02RVMgGxzf7hDiNOpEYDp6gkiZPcMpXwwm43nnJFPpyiWt7xhnkUdCtfyBJLoC
z/qF+8F57gc0QAExNnIRDiIMdxz5nsxd4KEkB+LwnH2Qkg0obcqLTSbaQyQ8Wn/N6EQrcuBmpssB
EkX7y7HV4xEY3psvT52Fdmbdq/61zqV9Q/TMCy+3r9hC7rMrhxLggvm/KIcu4F5aP2DLMzuYkIii
EEZ6pACOCM5d0lv5n0X/1oCuMzeVFkmmBKOA2bhknWc/qrzBNX51ZNv90HFT49qr15/qWMA8l83S
DYQEf7njlKMY2RdBbKa+seG7EanUMVFMVSXNzMqEopAH/J6MXXL/5mbsoIqs10vNUvHZzdYbZJ3f
CNCq7au1dcEnDMEXFtbL7ATwMPyHsXAZ7w1nZJq3MEX9B99vKB693X47dnbkU1KA130/1/0hE+si
FRP2DYHyipnO2ky4YXd07CJnM6UsZmzLfTrgxKz8GXjbJ22OANottc5DFktexjqMKd863wfgvjQT
dYjom9TKBZ6E4YbZu707H4jT39OMXLdiWcfvA7FxlYtvIkvGTOwqUSYBGj8a6KqldkgtuVOv0rRf
4k2JWbBKO3YlxkgUAHZG5Sosx/ta3FBTkc3Ye388BoDHSLMvX55miGhf75h3KdRzDSA5rGagDt7S
gWyF/46bWeJuRwjFggQpuOJR/9NfzeVRKVYeYNpRi1cMMM+cSLoqa/MbAO9rd9tqax/yzePcWuDs
vPIH4tgnx7YJTf5l+ziE3VlbiuwsPgqX1XEY1feiS53aqhIc5nehRRADFIzrpoAH2/TYVK2YNgVm
CI9cSUzvSgCF67ZqQASx7ZdCNQmb6cqTIvXpBsdtIjR2kiZGlP0eb4yzzCMMpE3C2y5JFQJFzfHY
riSlTt2KyoIX2pirkJkBpFIlIafmRPsPHVF2SORKUZRhC4Jf+mb5mey+VhSyUwbJpGipBtkwevwK
6TpkCfQDEIG+6eyvuxJGZjL+1P1gFNC0fPYKrxLoMrNK6Ch+2QwuuyUy6x4DJKjk7qB3hlJhX8p9
sH6+pa7TR7h7KVhOhiCPY/B22jr/DLYGE9j7OJlN3eDEHSU7fOfIvaec0Hw2TC5I/jzwgdAPjNpU
1zglyn+bwdItmngvWD8iOfRb8+XtYJk1MVE4pV4ZX8M68u9E0AsyhF9eyPtxXAER18o/ZRC3nZj5
rxaI2A+nyhTl8aJrV7RjJXPIRMJzEu0Ga4jhGH3u2jEl4kEaBs1vCiX9B3kZ0ZDEETfT24Prz5uA
dLEQADNkI4LdQQgAHN0VUm36/tGCEj+zQBxzE/3TTHBf5NUWq1JS0I4t3yyRGv6sbXSeuueNTo4a
eqpjlTPO4EpRI37pw/4oNyKfsqljy91/b1u3oCPT19KJwKPGSf9LbIJOHrciGcIOBCO4iIjHvs6f
WYUPj2gzzDVeYJv3FOBeYIARNaLxIOvu9Kh45pKT4luXUuzQz6whqvoo6aTAwCArno+KtLZyQmC2
b7w4/meh2tcNfZlcdBSElIA0F5bgox0EZqfhlas4EaoTF9BpCea7sRh+GzZEyBy/MhJhsiWF8ftq
x2JVMO5aYGYaIY9nK/+cmHkvZTQApyMQO14+GA4Hpk6wRhPUnjPdO31ux8nEO2Q5pDW/dgWYLFgw
KXbwhQLq8TUF2dN1Pzthr211W6dhzMSCdJwj7VbYCcBfD+/GUubeCqc0OnDUbv1MKB/gCGzTtm4A
J3VwvWa8MHM6bfd6ZATmUrSc0SMjMeSCKTNYXnW2oCqckOxMQ/q69emSpeq/8tNIa4ogapQl8ECY
YQUvORdLqJJ4X8tvU1MT7WT4mCWSTeoySl3f03Tq5NxQWN35yh/oLPJD29nlAZ62GKqSWBm/pA5p
Ai7muvPK3g04sEs9LradMiAmXSjmq1UBac9oAgsecF5As4zODh7DNyFCfE1W1jW0+VnQ6S2z5d4/
2BJijwGk1obKevAWmoNEYnvFbabUzU6E4Y8YUIhUtThQUoQLLQpJOZ/0q1jjxKBDeK7PqINSrOwd
0YtEMabba8CQdo9zIllES6VeD82xuj/TW4M6pdhR9b41QQxQclpucmRrpaZJr7Z3TLA1T8ozy7Tn
lpNTi7puvKA3HaZg6KtTxZGmSkEVGmft/eQHQe+86ZyCvXcDKvtqxqpgGD6BGsgbmtlLqpGzN+dx
gOeTgt9S+bEnKuMvpjznqr65+MKrYkDDw8D+ODWIZsLJM6HLrJ5oOlOQ4cu1Mfy5RnFsWbU1WN2J
y1Nk+6VN55hJbCmzHWL1+EDN7pnx0xP5aqZlIrs59igsMvSjHrWfvqqxJ9OmoBcWSUdUMAfTP2o1
TD3f6qX9saEhwmvIlQ31ezl6FxfxGLXNHXWStqmNJZsf10OJbIfGMR6Ibb32SuLcxGK6TPYXkCd9
/mUVFNmEciVJp11JT70jEX/YP/Sedsh87kBAa2I6y63LAwBtUA5dtLrnscZbgvPq8IISl8IZsvYx
WY37Lzt1cGK3sq3sY2LUTjeJdPN25biGeRTvSbiNEe0uCsxCHQR3oTlDAGchq1KX/sxmQThFRMna
jHBOmxNxcaWuicCfvN474fkMUlap38dNbCeW4VH0JTWRCFvQKmdEWbXqtsOEgVlsWh6ZiWgr0B5k
Sshc7okiu1yWL98vx51FMKri+k410FT2xpvowIPUQ3bJrCPi8YQSeE8bVE2EcwTe7jggH6CGXDf/
IgopbiRSzdZM+6WxV8AA8u19UyodJ46oMMkP1IKpUDek+PP1eaYMQoyid9o17vZAR1CrTQjpJGbK
qpSr0z0sgNU301EUD9Na3Khqxl//Ud1a2lmcSMmYLybxGoPYfy0AqSseq+bOqrkrR0fZL9xcondz
BPFD21aiVnYH/vP2iuHytKhAyIHcm81oKLkOdLTXdRZgXQIi1ZnANiHQdRdjtSAKsVaxv4r9QR89
N+kO/k/Y+QokQ7xJJ/ZgTGRuUjUZpBuNztVd0CNUw51QztnK5e4v1udGVmGgdCV3A2IqS7+n8mJe
SyXQdjz58U3ug9iF2pBQ+D9XJlFNWmQay1sxnQ1ew7ZhranwKCl/2Kg+2KCK/a5N4W1WqGyQxF8i
sfbLQmoCq6AKHebBjn8ThCNx8CDuhnXHFG3UrgIUREwf7FIX5N3VatCA2KBYDPRQvHKCwzDkaEZU
Aqj7ihCN45qk0ERKuTK3D2gAyJNo8FBDtNAmBXMf9Ni6wjrEsJ9OjSwLweizu3LqrSuB3g5ETOZs
q88U+t1ggBDfrjT2rk8Ii3Ec1tvmMeHERbxEw65HADIwwoYpHIYJZ0zJf9XEojn0JzAshDy+v+r/
kE/wHUo5tzBfvsxU/AhsNZiFR9UeQx2FEADVOq5jAD+Git+HKFJHyLcMsno0uwS5QT0xT8KPYOsn
z1sdy+pRECQSGq0LwcSHyH9OJzMASElVMnosDeHch21pPylzT9VGDKo2NmKMFA9kzJVHfwSzyJz0
amG7v04sKs/zojvaj2w6Pqh1EEw8+V2mAiLG+IbbWuLpKIxXp2hF4zemh8MQ+BRCwErIDipBF7eq
nRrGRaNViG/QJ5ANtqDugk664HLJs6amNGwPc7FVoMEbFDc0m5hygsw4h83EHCt+Wntme/N2dcfE
p66ckR+9fVmXfXwzP7bYDlyfOz+q/Kc1kAh7i8jji1xDe0NUU00DUP9H+JPnXmVO6y1TcdAeO2ae
QHukA7I3A1qA1utHdKxXzCIq2jTsejJsWcrYbbniF56j4RQWLNcdkv/2uLrigSmpKO9lmkSskSoL
bnIp2qyZ4zGooftHCMOwMSUckmUtVWbVQbx8YNT1XYPi3Zu9SbdCvUfILF/tm4NEVwZmFbdbNjX3
+wzGSX95t6xFdXk2rOpFnWmeO8dPxHL38lromrvxokOPNoPLqhZenIDLgIlTcAdg9xIhbWbBr/7U
QjEg6q8re/teQr7m3Y7H6GgWsRcu2MF5iwUQqS569/2wVEPbdxWEYzQvXDJB7g2zyh/SEWMeCal5
0Vr73MENel/lfBNS/ZX+OPC/wO7t2KSGwgor0OF/4SprYYTwn9fLjRtynGfyp9LTiZtiDl/KYCVm
QyppOICLqUaGE6guS3BkTLXfqbuWRYW3qHxyMR3U0tvtwgG8vHXtysVKZyJEAQL2enIZQSmca1X4
zr1J8gVfh0/DEomFArp+ZxBsetQEidIoDNYRqcUE9oQXNSJ22OylZZhFdXlg54CMUK6g4an34p0T
KQKyCy+dAGgc88huFutuceCLWQY+qxyiN4SjueL6d9+TExpperolWSCzNMGBLqE9IV93UOyyR0w8
eT5zdD+n4W7z4tpC7x3sjUp28FsAnV80eCKWertRFDQIe/OSFm3quCuDBmVzN/t8Pj1NXjOKmwQ6
cRYngaVWIQfOeB3S3hQLhDM949azO2vDLPGuzB26TrWgreHMfMoUmxX7rzXfZTwgkSS091DyMk8M
i8rNQEZDglKoFuHSs2/BUkNWi06VP3rmh/Ihh86iD8Sor8I5tEkthrbyczA4cYNbR9LCpjZ9ncTp
DY1stPFiEzmZwYB9sA3xSD6ptwlmnSMgw2dRAemZn1CyrmgJ1ivwtLlBYk+rflKgzI5snLp6iaIp
BLoGQKfHtJC+3vJPuA7x/KlJgaXGEinKiRWN3K38J7UVNyOCSNYEnBfpzAFS2KMPT3X3cHWViHro
UKC3s1Llw7NAr+onv1j/tdFFVj9k9RlHFmER7iJGxuXF+hRoK7Xbmi+v6f1G69QSCnMtYmy84koX
lPPg1dlF8OajP3Zo69ShF3OV38FJz+jbuPideAIj68QFbxiX//WtyEuTeg9mVIUoCYD3t4oO0CWB
6ID/kK6eX/VUsDazkx6WkdLeuRHrJNBuzbobkwEXgCJAZWeJkQ8PD/wO8Eg2Z3wJbKC0wxbj66hK
XP1a7iCNbowkPCuQ3P4TyqFSm+waI7Wc5BvaqWqmSJ+/zBF6cqFdBzMP4HPaGHa299FAg9aEKofm
Ken2bIahaSN1NMbe0EPX1kPDR73a/8E0EDV6cFqWvZpyd8RMM6Jnk5zf9CEe90qnf68kk0NOMYbj
qymK6hcEDyclxJbY+TXqTnBK0UsI2fiwe4zAo4m4GBAhWdhAZL9Q6Hs/VAIeUxhoeuW51CuMq1MF
+sMRFhkeprexqx++Ksxn2CGIt4/nL7Vxc7snFzk2XQwq0scAd+3KCFJIBs6LPzbUjVUpqXhRc2Q/
C/zsgxs8REJChEDqbQ7e7qHqvDf5M9WjYkJkd3bg1gtAfOpHOeQ4rw2dzxSGh97LGFpWgmShFBAV
v2VD5UhAg+CbzIbziyE+T1TheaiKzfeSo6WFF4ENdHEbLC4QQnlcDvzXk9atPyreVebx242WsD8J
86PiSaSkKJ3wTPEg52eKe6tSQHDgH7d6dzbcS9hNRlKo3XLHX3HsS+73OeRB06HU5CIIE2glfaSe
5sACVmTHuAWuPiD5oG9zawEgLn6zlHXoZJXzByNBUhuXjG3l59mjW6nw7LByZEd8hQmXHybEZ5fp
lRGUuApnjDodaOdpTAo8VlgM36sJqO7CF+OZTvTODyBXAaxZ0NtTlO8PsI7Ztcu5huTWazxb7JR9
SYCOgf5B82JB61SZY6BF2+YnaTRz7JSt+Oe6g3Lq+tB4vstmfBE5eiyAKCHJMtt6NmHgGV0lXZ82
AYmdWCIxtWxuPeazoo9THAntS3FJK7bcPiJtLWSfmjl4aQwgeX8aj4t68QaLLw7ooTG9TSLFoX9e
Mjb6QjuPeo4SFck2tVzW4QujQCTcIMjxRlvQOL148+XmVS1DRz3YWVoAU5w3bvQJDKaGaOUqY8y3
MSAWLbkelbX3F0TXQsJnyoMLsfkWswvmeEUiKHhoX+xxnTgrd/+xqsKV1LPdec34KmO1XqN2PhUZ
W+MvUE6L1azALFyMfv+QI37hFB37tbnxz2XB4yPEdzBLSbUPhjfgErU99Tg0YHw54NBu1eUhIauC
tYrbZTrs0WB332Bz7N0NroJhjZZdyfmKJDMdvweKuANJp0Bqa7DJ3HhfnrJQ32FHhIppk1hXftwv
QFsvbE3+PEzxbxeao6F9fFMx8EJnMLpIp9kaKN1/KMoWzBLSjMcbdtL3j8LRwO74SGpii+aqgHlS
TU+59G+esDcQLJgbo3t+QeGNGS1XTE64zSXiACH6xqY2LxiVX5IJWecxv70b6+p5cOH8rn0CerHU
LyX7b9gLWjVGXOktwXyoAb+i0BJxr8NeE07U3JUXd0qZVeTgM9BrFg79YTvCmweyKxzHRcZ8Kp5T
+WNJDCyP1e0LE3LZ5woCId9CsQ00Ts0WfzWWv1jcXcUhQmamjGom3f2Dl22hW/v5mJU2+kUOLXJM
wL3Y+/s74flK9/tnA5yXP6jCUbza6UXPTRNJgw9laYjNvfvFnsF0vl3pAMjYSMA6x9YaddcfehS4
2j0DXU9JMZW4ZdJHBqm76716kH4XD+42EaW7n5mRjZN6/NoPDcjq3kZA+vKgQHmrKzhW598SrQhN
dkOyg5TALUsGerP4WRHtcLLLZla4YBK0KZVPZqpDtCJzYdRZ3KYAFg17X1u4epKhFAxSsbjH4Q6U
Vk8j0pzzgrUdD17I8sfwR+yUeWMN6UTJ5AflaXgc05T5tgtBkHeBu2t6cXnmSj9ooU5Da+ED9Fwe
CkN/FbBcZKF4I6ga6jLVX2is6VoOyRH48aiqEyufSJozfVNoq24dSR4DKCpQVq+n5QqZEukei1zP
9ajzodDd7lrT96nMbXoAHYc1ftxcTkgEdRdNdSFu2DOBs5eGQrCyvmnphAOEqqcQhXDHe9VXtKiY
3mUvuzWVyvXTTdkML8+C6/3YhXpq1ZncPPqb+CjFWD2TgRNx0b7FZtH0cTVxKUTf3IHHkW1Kbb1g
5tzAUR2DLU7nQn/7UDxJ1o9SLb0typ/+RjCjPsu2y7FZkgGVxcOoEHGZcSuXTo79px3WYTZvIrOo
RPs/vfWRhI05J31cfozoGFlha0H/dHHx8mTIAr5vuhbuW0O/UCutRYCKLQAUUhttGSH69dYcvTZf
VweO5u9bxmc5c1mC6XSRyfif1oG+6CyH1eMehTyBW2vFnzUzVASxy6bYFUn1A1tudiWJD4u0H57P
XL6tQzWuRI47sEFyL8sX43T2+FQJ/jxeUy3KNI3S7pRF3WXWu/o2hEw066OpKx715GDvBRC5qX+s
HnVmgQfqcU15s/QyDkXSPHPPzIweu6X0JtQrtqs1ZlgSTVbwPvYkVz5C8Y/5dQrNiJrghy7r9bgu
xk5HVmx9upKgLTJBci6KkvBebbj5AHq9NaKJ0MkbRqvKSij7EJG59OfyfwYWkdow/saylerfx6W6
evcWNM76GRzd50aJmd+/vj7oUMFid1u9+vz4tGqfnvtLKissfOfMtEl4PEJ6xbXPtHNlkB6/BILC
4h9yNbj4nvnTZoaEnKQ2N/ZoSGQwe2gjkRhSHCI7A5Jg/xtFr3kiy7pZnJk3BXrn7Yn0zx9F6Thf
1YqiNxntgPlvHhB5vfsdU350fRP6G7Qj1wX8nFWLK5rPsxl+8PJJDXKy5A+WO1nEH/nPoxggBCl+
DN3qnETZvJOBGw4EtR5ziqIIYRrgnpq01h5E3jEc91XjvgN2zIZwg8L4ELNjnGF0ARcUrq5jcTf0
WIlisXunO93CccwnQMkJeb3CiefUpUhc3Uck1jzQOHGqxPK0ECAOu+ToWaAj3KiAuTZKG7A95Hcb
HPUBxsSAaMNUFkvIwRtkBpIkq4C4g4nzaGSt+wh5s39JOEp4gNQl1Py6hBPDRQuOwJWu4IV0hRSA
c61mRCdROn67lcMArYLHdGCwFOWN3YXmp0smVRwvNa03vbQFyBkBXodAWzGKFTw5TWcciwapEF5t
fyeatpDBerEWEKAoyF2zotCUQ97nR75En8SefC7dBs1lw6ew3ex/g+zofmlVZ37Dy/IAWWw6lv/5
MU+lpWmLcs3rgXR/W/J5Q8I3XLl8EL8JlmstbrHINeO1jweHjpShynLtQQSUcepixR3KfEKQ34Uc
FCu5BS9RprZwOaG4O5HodG5BsGnNJkZ/O+xEv9dHBvm34bL/zrHWtVW3HKaoJIftWYdCSnCta+T5
QJQOQH8+iFlK6V8HmQA/KQVHqoTZHhb/PwDL7ZaZ92jkvAKXKA6c69tyl3uFRXsNJeB6CfaEF7IN
IBOSDZFLjl1Ujs5AttRekM8iXtAa5UEVKCutdtEW2xKiwksxZgZbt7lItzJPrLybf5245I/7FjfD
Etqy4zmer4ffOx+wtdtQomDKVOY7yGKe6UJGQPvtsvsQomXsLUuwsuuDTeMaYSMreJaulBc9CYXf
hED/q9Se1uYuRoUgKH42ElopjPx3xDLiYDm2x15DgImE8AIAG0HXSP515u1OT0XBFmTRMFZBn5KA
XAAjV/H3hkhMXqzSSRkMuIFJjhqUwip8ejX8kVm/itTaBYriJPiL5Ohdlciyw0FVeIlcp2ClVnw0
DKw9x52Oz5Ub10evN5n/2cYoBxgYgcu6fU4IerG6fWfl3lof01MICyyOYvqpLQjNgn1rl5/cuN4o
6cyLASnlotm7Ou319WqOwuj7fL28Ck/UFQX0PBiPQFKww82tmNk7GsAJbqhvhwS5pXmTLp/p83zZ
ciEb3cKcglf/n5vYCjBTBGTfWvf/qviJRu940fciL6lpdOnWKJSkzQIJnLR7GvYp9biSNU0MOXOy
tq5hHkVwHsdGLxaGHLUDNB9YJtio/dzNKFw2Jb+nUr69tHxkfqFFf8MiBckyajyNNVl3LsxEWrHC
vTF9pssuGPdsmQgyHe81KwpF4oMLlvf8Dva7Be4q5zeJiCvoEZ8SETEiTBPh+aDie1rQhRIP5FGw
O4LgOvgc53p1XLg1Dx+BgNX+yG5jSKEyZTWIRWC0rZ4ed5pF4TRejMnZtQ+Zkc4A/guglqP/a750
jzwMzmI4d5lE5Ynlb0BQcrL1nJDL+r9rr75IN9oYL9kRstMnz/YwRFJHqNSS/fY8lHL83XszxVF5
okL0WcBgWpvdUl4ppunT4hwR2iECz65QJOFf6OYPHzdvwqPQ9z9aWOS/OQkvhSwiJ/y7IqRkae67
sXsn133EBc3SRCXq2+l2VqQoc/XWIoIlc3v0rF0wJXU4agYSZYwFTtexKZ0Iqhr+iugX+PThgD+I
VZI27AgKdxHHyGbFVel2nwZ77ln9BLyOVs4Kix755Q98BfG4/uv4ohCdMo7T/Euj80OXrXojz2kO
4QNB2BP+8QZh6YjFc/RHvSnFOF40CJzoVsTeZEjKTVSmAfCCzQjFtlAF73XHtkuhLvWPYqe9/zP1
j2FKNKXo/OyoQ6dJlzTJAMMBJEITdybhVW8yHDCUFAQQnsUwBTLXD0c1OC/C80f6lf++5gm5FKrW
CIrJjAUkPBjwdAYB1xID0DW/qYTmQb7vzCPSIgtUJZJpueGYCHEcTeGZ/3OzaUVW8HCGSvdULkir
B05PDkr3X2XyYTlwKYX5UlYKaWEiIeHy5eoMFAilbRtrW65SCG1M4ZGfJS1oyB20qxIgcRnF+znp
kzmOa4ehZPvnu99jhFUR40x5r9qu1hQAf1BcmUvGfUXd4zKAHxHb8FtUm91nG1NOcIAC6uvnThWw
l+TJqx/nWqQCIMIRPvxf8tc0h8ZvfdzKpH+QysOxuJYXOfVatKKuLvYyxUlO+8+MCZzVYBly9Htx
7n7Rwgu7AX6A/hQOqh3oF5c4crDwnq1YnuT4B8MkDEOu2P5IO7tlTCFiHTqy2aQyFBbnAClJRGnn
cXJr/tWZSLOY7KCHQzUrwMI5+gXdUn/vzYFH1maebBfcqhC1U/SRffJ2aWcZVROfqONLCIeqVOE6
aAT2wO7yck5gQKhcwqLg/AN53cF/LeXr/xJb+nhGI1flWPoGs67hVtI48eKPnjHNuSzQ/edXPHcw
WEG2gg4rUTaYnClnPYeU7YLxMED17DRNivl8g5K7GtHPMCEo77Yz7pr1PZVU6MIycCskGwGCOaHv
otk6EtiFxjoqYg6gSVpGcKH57af8ydJICzV701cvSvUQhW/4BQOejcJbEiOrfrKLGas/YSRTwJcz
m3f7mWePytag06L4UwN0wuz37p1sM3aXUTxQt1e28/LPrVyIo6yGV4hMVM2QK+hXb5tpA7cOFKMD
nAYG0gkMFICq1WABcMMY4VFp/8ui7SM4ZomM7HEn5PCdT9SpphYmdKupaGcogdJjdK566/ygFzd7
jDEiie8FgMDdhMC/F4Dv/9l5fz/nUrdVA+uP83JHOavfMhB96yuMCP1HpFXPiUsQTsGxyDDE7Qgw
kIUCraO4fk4sbxogI7L2m+JP6y8CImzFOul8Th4HlQDrPqD5Li6eg5K2G7Uhn6KGgb/hpapdxQgh
p945rriIVh7uAMAtB7rImyuZCLLk+q260zm5uPjJkLfpbIKyulegnweWohAyhpwZp8HpoBr2XtEf
0j9D+HmmUb1WL5/C90tv+/2Xf3TOl41zh8WvXqmSjzRNx65IR3RjBJnJl7iCmuLtSEcIwsitV7RQ
2R4FGnki5fxfla5f6vEjvGG29hLPpx5SVU53tZqf0SGWf2G7OCOFfL/Q4CnwqTC+PrladdigJ4AK
hkKwFg16ShWYOVQaxesAkaJKwRGnA/i15QPtYhnAdP+7imsl15QhsbjjKkV3ivFBuXds/M0bJwvR
TBjwhs3mCw90U31YKzoZ7WKNF9g8p5uZsXRSqEyxtilpzRVkqiqU9aW6RiXLvwGoxi1jdGYOoBtj
PRp3yY5dRCci/hutj0/6WPWsbHtDS3yLk/DZ8ZfAEXQQRR8ExF7cYweRIf5n6jr2p9m8mj33uuXt
GgdjQrl2ENqBVGL+y0yVnMUJnl6FN3LppVUJgkSiNLiIAoGTws32WzQ3yzr5dqzgb+SdHSweQNRj
FWfqP6z12FC90dLr+LROFDn08KfQRamawPwXDDX3x42cHVPf+Weass8pwyvmB8Nfz9CBZXzbYZbg
r/yFWBk9Ik9BksEG2Q/fd+ekOUjc/UzgzEs3jkv7q+AsMn18Dl7MmgYZ7DDf2Tsv0MPl9wXHUumH
UaCp4f9hCD49dyw/JUmKJn/nmH07cgNiDBh2TxtcujL7UspXzv1vp1TMxI4CGLfIS4BYPfsxpJ3w
aaBg132Rnha8nzXjz3zGsxKPZUvwTOWTKIRyBQF2xitw3py3uJkqjKYMjtawD6U3nY1OvkMbrt1J
rC7LtnvNVbC5LycQ5eNueOHCyXaTGKQL0xwDhRV9jZ9pvQlMakKM5FFxI0IyU3KWiJcDyxTTFQum
gl51yz2/ExMF4Ztxw8/wzRjpMg7WNmo5/bLSMVyL2RKPZGQ8tU+r4hKPyC5WmRikEFKV+nG3UMuB
q3oFaCq6abMgM60OUpOXKAFAdL5wF57iBzoWxR+U+xyccS3/K139X7LhWY+8dzqfvzqnbuPlPSIl
hGG5lFPSVho6ph7MtEocDVgs1Ep3wmnMV9asrjJbXdI/G5IYrFbXQP715HXtH98DzOzK5lHMpUuL
gdxQuFkXvyRmCxUYDKigMJW5SEl9dN8eK0G9pw2IEDpaEZUfM7L8ksRo28atUjEB1wlnqbxTJGL7
7Z7CIkKNDR3FredpCPJKXQV0nrDEFoBLgMWXWpCEhKtuFe7aWrvSnUCNB5UGIZlrVnfweHKvY3a9
VjBbjx+gWCfnfuUmmVdcryn02/h2lVNG98a5rGM0mPMU1dsdn0GErlo88amFie/EMrL8mreIe1nE
PmufpfUC+WnEb9hARSVXV+gNLZgTVKcouSewn11O6mSQD7OpqlM6GotlX4VvpdM6EzZyLmX6x3Uq
LVGy95c86Wyxeyi5lr47Utvemt2HN8Xyf1WIkToVPEOsolJtQN2ksBGNf33tYlu6nTxeXsFIexRv
ira8jzx6Kc9gZS7fNGHMidwzLJuMgUJ4d6CFqUxy/zM3ltexXCZzI7vklb4ghOesH421xBFtblLl
yVmk6QO+CRXwHAK5vqJyVmB1hI7QQ4sbC0DUny/4lDQArXQMlThShT5iP3L02bMmUQqQTRyJMnLk
OAEa/qg2ySZUjKPnImy7ezOAFozJ6GObLJp9Gl3ZT4Idi+xZaQUkXzkY/DlbbTrd24dq/kCxdKfT
OZRED+iGz0Kh8nvZrv4Ui0u8GJSuNkAp3fcojv9kJWik21+iQmFglrizifRoakcE9CfA4IX14rpG
pAXtmGyop0v8on9mEas7gg1yO10KFAonxbqInTPK6NRKl0fTH6LVutd5BhFQKjxcFx5bbmBKXKF8
TDfGCXKGadARpOZuy9ZY3lwj9KrkDwbJZzsHNDzd02bJ8bpwiGCOeL6znq2xzpl7fy13gh5TOoVa
N29IiYHj12I9YosJ5JPWu5DtrGDNh+MjctUL/jTlWTlvZ4ZQm5rqlz5saYIduvJI+rXqv8s4nZNf
V0V8viToXit+BJl6fQ6mASmbSOeBooGaVRGoAKgPYfDUOt0itKI57DE22ljpx4KGSHpqbeBDIJa6
AU1J9lRJlT3w7ZXa+MNUEBB+qmm9eegOIljrUZxUxqs4Ius52aznALk74kk6nlD3QSEIWbxqB9Cj
IShMAhRr/JgXkOpUWpxFgQdRDVNhV+o9PhfCWgr9+uWkpWvN19j4ecrqjn09NMegEHS+bqforRn5
1xnh05n7bt2f3l2RH58sf6ZSX9u4yfsZNtc0+w4q88HhkWh1b+2LRXrBYJ1cgtKKZbnyCrkUNvlR
6BifIM+en4N6ocr36wttaS2l/tdcH9r7KDhluxGvf15kzzbhpjvkkxVqAlzWbld7jsgRKrmJqZ02
gzqsUAtcfzlh2itA3iOVkXx8nvtlfFThdt8ecXf+pFx+bCAA8/y8pX+bikrG1MLKE6BCd+TLJ8lf
bQHh9ybPhIiKcq4VEq58BdVC3vu0Sc831pV+1wkh8w2X2qTRdyun1VNbF+LmFVBpTj7vMyudLymb
dLlpkB7tUrEiN6vpnWpu2lXM6EquRUyHLYa4h+Fmx9+TmBmOz68LtDcszM2dNNJ2z0H3VU7EJe3v
YDkIZJnPwbZ+cDxmljbfQPJ9Q/5F17oyDcC9EsaS70wEMrnTW5sbWx94M9NtMzOngGK0Yt25tgbW
sDBa7Posmn1DREI2m3bUGcwdotAF9jMQosfuJcytUl+lRaOBDHjqnYIJQzjO9njZl7I/1QKqWN0c
cB9rQJhXKVoiskYAklgi2oCwUjvSyDx4KX8VJ5e3Q8q84mgGp32KhR+rvWcflYWPAe33EaEzYBV5
QhtMrpNgHEjsaty7ZddAT5KsefkVxEasKVor8aTYGhLkuLyBp1h0CtBqzRn1WMDTgcEAo5FCnmRx
388KNshNC6JNqirpxK6j/U5Ym8d5/TD0F9P4HxOTdCQ5WXnUuZlAb2GUflDh+qHSLdE1kM09a2ql
/h1yR+gHVzmUiZiSOFQJbYPJTHk1MGkzFWZvFSGRZCQVtHzTLYMRApSaOvJC0cVs3X0cuUp9IBw/
BTZbhzDS17UcMjj2+zlXfkCy4JtCQnzfPRyONIoyb3jfjBVR2KoryBSgloGq673ky8ScK6jT/dlw
pCAm8IPwAK2p1YHibMBO5OnTLvidggvpFYACyWcq0ErgYcXBPpssM+JegSr56PLZlYVqUkHZx49Y
UVbwWbhadG5eafQPmN9c3xa17jyr0kjbSVXYEmsPwGGUDwKt386D3x7yZm+S0QuugYjdR+pfd0SX
kdbEcE7GbWTA8qZJ2xFypniv6n4JT5YcnzOW/o6UuFAUAfuYSQUrDKNPjrymo7WWPHv057GbJnef
n59ULflEQLmomLgqs4EVbQd4YGIBVGzZukhYvjt2khd18jai7Q+y09VlgzMInsd/+NzT17PEkw2m
nEZ7ENIJs38SDEbf7HZWAu2r1/1Gz2O/TcuUCoTUN3Y7+IySczMQe9EgxsQxDDl5qLkxxKw0TdpH
BfUQcBy8vDQZ9/1BaKkT7eDv+oaWCwE3foYfZ6Kl5z4FEdQeEzozSltcIsGI4v5NfiuBkE1hmwEd
hKdYctNKwOK3qqK2nreokRbTVhbl5AlVBVj67YEnCDrsZRFWhG/3PW9mWCqucXmDfj6YS1kC9I/a
m51zgkI223Mx0m/Q4XlqybHuOLw+oCphPZPM827VuihsFdBpQfDaRQcN3ebAEwQfUPrnmlFrQz9b
strmlcG730rb2x4rgOc6ua5qt9q6C1F7HUp/gcD5m2q68u/MxB0Y+3dkuzNU87UbSqTX7/d5zRGp
qODHAFvHjyGzwlbtRW49pJZzklG6nEIGx/Gz/AI0LcgOC54gGAxYCmxyyBpLLnIlLLPvF+1KDvvE
utAe+GPNPj5dNLy/a5nE6c78uAGQn2WEqQZLfrng7KPQE9sPhy/0d3BBY/I3iPqSzookErDsibcI
ho8ec7taPoWMddtxjB3EikADGGh1oINPPYbvfSN4KDWKJ6qE5OV2cDEXlO3scgq4sNDM6If41ghe
n+iUjiN+BDv5UEa5EEMLnxcytepVjztVccBnXfdkadFV8gLqWCPLAwGUwV+EspJEYTeJ/Auzflt5
hqbtRb/be9Y325IajmVTAvRjdvzbISXh85TEvGbjmOCkTo02XJp4l0EX2jtYRGloqHppUbl1hLU1
ivPXnob6S60rcf7JPSlJBXccw6qdRHpFfgXfWPxibYeLas0ELBU/rynHXhGKFRT0OUIMcgPmhSEx
PcXsf+JIfEH2aqtiPyNFumwojD573AWXOROFQNH14FX/GXDBnEDmq8b55Fv1uxxL9shdddk5Ghfr
+Lln01htdrimefZqqa+ZBLjBZL5DzSyvhqS/xEkoUDNDtIqbzQ+OCQ7BLEg20gSWqCE142p5LjTK
JEAoFHxu1t3Dj3zvWZ+bvDYAFHj4UCsy0oFXH1YL/FownIy0mZW/E70gNtJc2LixRhvHNFoElFr1
GIc0S/DuX8OyPtBdRmEhv/KDsSgxhJ7FkdzTv5BxB3Wnumg5e5MT8XhMl8ahKdkSE9TZtTrmw3pR
L0/xKVzfo7ZAauIR5dUyp3GCOUztFA7l0Ivohum7ZujWAZ6bci32dL5hFi5Q6qPzk/EmkRgiMANF
FjNizVA2iHwsy5PdVc0L04CuWBeS7aBp4wt9epMqAywxgO0kEHzmDCMdQM9e3ymW4qBB2gXgX2q9
HocyKn301WKG92tkA2a4hd5S3ZdCNHIs3BfSQUWjxVw/wzNWyFMijHMZdFy8WjNp4pjpLZUoAl39
238Ow74OokTgaCIRt8/F6A3HSBWSX3PbLBREFslYC55OqOTdvsnooZTLaCpOoTN0Gc3/kh2g3kiF
SZoQODlN24jGvaz5OuX5bxqN7j0oVbij0D9Fcz7rruIBEV36bColxtx1SPzMtzcZFvswMwk2CS22
4tw9EKG9WMgayKpVacN/XS+MC7O8BtYBNR58an0EPsmiBZJOGWEeBZ8t2PByAwrAjee1ilZxFuen
QdiCAoeRUpM+4hjfGzBTeghpVzirDb20XsQxoP6D1YVsYoVHsLW921jx1OOPRm+KFEixW8lMQZr8
LRPR/vjMBRl3i7gpvswjAa1A/1oKLgrmuWE57MVllvBKXTEToSqilKGyHGkAt624Oy7WaL47GkgP
LrDvCUmCHZZ7sKX/8fcFl5+c0g1CR1vipCqr+dR3X79RK7Ib8Tjn8Kbyq7RD38XIOOX2fZ0H4flm
8sK51/lwhJqzg4YGt7kahYv7JDzXfOqB6J3ZPciNZ9jehyfeMDYxAK2iqC68IH7OrrA8d8QV8D8B
DuLuWMXSgTYuOv8M3YVzCqfMj8AG0vsMvh5YpEtVHSv3BBCy6oBniNH66cVgekTjR+McDbBBAl4R
qOBU+dn6H4zB3X/PPcGKqbME3u24bcTirabwqIhJRC2TPIxkEbNoR78zm+tSlVIEOXzpsYlBOkq2
vzGKr4yTqJYUdIwrV0iNd8Shv6Eow07SwUgxaQqGus3HjEGvv9CnZfLiCLt6Jrg81R9jQihZk/2D
Tj0PbTNJQ5pcs1g9Q76K7qpK4LKPc4k0NhwnDW/m7TPz8swP9o14+YOCoVrV0af03RRDskHs+wUo
OUr2ICOoj5lvrBiwp0Pmlf6Vsb/Kf4Q3aO1d93FNOWNzFlRblqonq/i/BVpj1UjzdKaYjYB/6/2X
YXon/YexW/jlMJ2K5PKyjHyJSPqDtn7GseluUU8kUqOoqUJ+GdGMJXerMhvJUhuQwlM/jkYGixO8
asJBzjk+/73z44X7wLM65Ndg18LcRy6l38yG8EIhZVFoyRJtqdSKI+pzekE4uU93M7gF9AH7vTf0
IYC/UtYnMyHsohJ33YZM0kw9e6HRDZxtVeH1hjoYZSbXG8YUM6T0LfgEvEgrqKW4XNCFMz5pxEq6
rGqbdt79sMZnM9IVrftjqUVi/D9bQGeIVJJ53ty97IucxVzuhignup9KkX5+ODUNpaNftRFNG1/P
k9wdXif7DmKH1B1Qc6+5BT6zk1PyP0PQHlqt7b+DBtZHZR7nLtV7adxSHbFcbjvHSa5UXyFVToyE
ndJmGM90NrALSy0rQPEN1FyBDWYOQhFYEOLohgfQVMrvkpevPhmT8dU1gDtns4h9IZqPHJtpX9sd
Q0ybnWud/EgyGFyPFLL04N69htV7YudvWBSJVcfzDg3+jTfXWla3zYB8+bchvd7yAfUeg6KJVrDe
lOFjkmmJ/uOPpcuT76rpVB/YPeFvLaWnWoW+55bjcJ7nRcH8B3tE0+14pJuK/LQXfsRAgIpzaWCF
4I52eD9JB8w8vpfM45A8JtJjnglGerv5vpYMTkgWAv2y2dP5tThlwKrdrIo5+3Q9D3gqiSVcG27E
FEHtRFYXmoE0dNubAM9rB/+Ynt4iny7CxfxK53cNTbDGxauY8fKUtfVl7bZTXZrREmAkAYoSQx6O
uYph4NMdVIVWmnAMvKoP7EhTKkcaltPpSa/tVwPeDTFWyZYx2AQA10yzVfs6X7xRLuxbcu8Cb/Zm
Ui4VaQMFNHotIJs29HMdUCcZRIRLTn83Nw+fPYZjxELIAVrShUIYEl6khjeDCyo0yfrAarn3oHbc
d9tIEfCXGSOVVf0aYv87O11z/+THiJYCIN0kiylO6ZJDAKyBGkhmcqOk29Kssfy1THHIqICp3Csg
t6BeWlR2vumSFqy4iO/KWAVtUIRxsy9vZdemj7nTs+46fc9mG3I1hh4mlq2/hIOebjGmRh2Z7VKs
wJIP/XNH6uVhqUIz9aT0/JI2BkXHdjSID8Imy42ewb7/Dyi6X+MxyGCDc1buoGqy1tYV1to6ut0+
ET+hunGfEWbCCWUPyawc+wN7qP48E5+rP8BWwIvPJve7JZWv0rTY2S8MEBagvTggX/H1yeoxqXEf
93nj1ZjjyhY76rbs+c00sJPy6mmLVGHOmLsR/byomod1k0f7klrYk1t5e5oES51drz+HGy3/SCaY
k+uZuYQOvJUKQUUgpk/JWb3b+/IuiMn/WuhrW1AkM1GUxzI3BobC2l8MZMrNWnCK7n37QSAlV7V2
pm00zc2EMmv4VNWOLaOLCRm1EGWei5yLt2GDb8lGA+Y8W65Syx3ebAtxtHKtfjLlBaWze0N95soj
u3YFoJVNmaASXZzpHqdZsg80Q8V6KEHuh7DuNFTj5Y5A+S6aHs8zqh15e7O3VfmnRXpQlAS/zumr
fVx6/9C5Bcgdkki8XW7qoim9DjKRgvPQkfwl9ZnSGfpj1bT/jX2Y8h8huf42u+A1EK4feRvTmokO
IB6qRQATFmauNuS7VfJw5WzAT2oDsa+zuJvPipHf1vYuV7xAcs+h2yiKSaKRXBkJ1NgcQs006fHN
TKdWB9pwcTuc6NuDNnrDYtgfyfHIDFPHkwxK0PFD7DPmnf49sp+jzORpHYvgMPO9I24bjD9JtWMn
4ZZIWA6F4pK6jufHDyg5nL/401zx8LquObK/kZXjjmMwgumRQoHpX6zpQgXISdWTEELCVWjz/Zwc
7HQUtLReCGpGjanRwGZ4Vfqd2cAuNEYrq2jIRNsPqnIrYqLFTkQEzbQPjfiYk7gk8nHnsaDJfLN2
SyOYSndVO5cZlKNwJFC6lZvwCflh835TbVleTsw27VB5IbSlAae8fdeeZ/KI97jMSuxq4O5VbPJ9
nnOxm64fNHmpPJVY8zywgdFOcvzcc0igjpoq0dzFnpcHz3DGM/9AF1EqajqluliYTY1IXohW3c8k
hZMR0/exUcntFDpqI7zMcRsE+T7BbjKPetiaCmnbFSlPtnpyB1ajv3vhfvwCoH8VK0rDuQK0SdJG
mTY3nl/JJZhNKm9N7gUE4Y15qUXIYkVstKYT2iTSDCSZN7GaHRk4TON3Zca5GnV9+kQAfG42EOR7
xDgNxB36JQZDBxKfmALTwX5t2c9/igFlNnqYrT2CgxwMjeLPagKzH0t9CvQERd7wwfU75+iy6HPX
PHro7KEhUle6qvqE7YiWKPzOxcUgUe6vpUp54HAH3/aWUylS1xKfOhWgzzvzR0wIVO1CJ2mgcey4
w7tUOhbGIALJ1JimSr4T5zlTXHOLI376orot87cPswAz8K6hV2Ay86N/aEJ8y2r63N1wOGfgq5M3
f4UZk02XTL/WQnKKjHOE+qCy+O6OMufbBZbYhYmcFM2nolxgUqrY4sdU/ngRADhOSMQM18no3hKC
o4SGeejPOn6pEzCQwjmI1rZPcBrC+DZUs51RaNKsM+P5jKyC/w4beU8rlNj0oh2L9i9IbQcXd4Dl
+uOIQq1JJd5yXdcIqTa2XEeMc+07Gn2J1Pu8E9vBdtfnHdWfc7eCvGnla5UkiJiWMMMQLhHpMKvp
OUxdo1/biysMw688tayGjfJhYoVPUuEkfdpjOSLCIOCaq3dzOfLS4y+1jhL5+wlbVGm5b3a9zu9v
CSTLKxcTofwspk9zXbpiQYH5aDUX8JF0YVoDOKSWCo7Mm2jjY4RP4jCUtsHu0SqzqAJf1ps86rOB
qCSTN5WNJEuTH+82GAewjKgA01VT9jUScc139qHYdwfQx6GcEHlweu04+chEl42sBwfjVnNWGxBh
wAZEXQVNYK54BPFkXWEX5eqDVVVlTegvwg8UwX+CZN6c4byMABx8mmo8bRA8OfqE4XYfAts7U+OJ
1/zPBzhh6KNAx6mebrpbI4Z3BUgt9YvvUu39mU+hCtSWv3ZN6a30I+0P8hGwk08z5gyOKdGCoK8t
gp5gWobL+t00N14kDaJlqDOLOM3L8CcSMX7d7FsrkOSoH2BcphBUh+H2chdGl7aVOexbTmURb2Qn
GQBr6fruBQbYQk1RmcRsEBYgzx5Iu3/LwyQj63YSo1bRzDCVO/UbbFKpM/Ji4ootDCPIo4HTsa88
jxTtl8iYlFdqBU9fPBdV5oVgJ+VcqmfUl4Q6ptk/mv/8rfr2uWHy/AZBzham1RxIrhkDyP7l3f/s
fRz6YmDGS3mu+dlMjltlpMzMcoOy/MxtxzkqiXXBbUhDirs87L/oRrzdaFuvo/RQGcNwMXS9Bi/u
e+X4A8l212rZKx0dVtUvoFpjOiP79p54o/q7FJ4kdTUHvZrzwT0Z3sQsJR6DiMnGcwy9D6dUVlSs
FESB7TOuBGQdVeUb0cLRj+tFkKCTcQTC5Kwsw41OnrUqM4rBTozWtxNvwrFlLfp/iFu9hyxl3Qdj
dmUw3GTEOJmaFHN+45zua7ql4SMqrk4Qw3HpOrgEMeG6o7PKjxBaROZjgVyC6Fv4nEFZ9cUJ0ir5
wktos76idg2PL3gZ6Ff7u22KbMqoelXSQKI371ZktJhBc6ITNwi8Kp7jjDGk8qsHk7mR1SMplyPo
hHtn4zoS1X3PZJZqbAy3AVThRGQLjK2mEMO/VMn2GrCONg1H0NX0lQy+jS1M4vdKSpbU6etH0Vsx
sVaw7g1J/goVDV/X/xt6+clyOnpCvizoUFxdkmt7PIOMmAEChkQsQKQ0VrKtxwJB2AOJhs3BmjfG
1GUI9edKknNv+dJatm5Ph6S0C+zmmsjpXIvkimwZgMbMzDYwYVa5SZhiEbmf52ghPO/isPHIevqs
wxszumPbLPbzF3A6VHT+Re23lSDo10wavlXqu36Vo/iD9KTh9KspGr+HNjgEtU8eAf89vDGd+XlT
mr7bHByh0X7M2RArnDuWnqFhy6ldLA/+S/dr8/3DMLl+K+78iJW/W+zcrPE7e1xmK9vZayRrz56C
0TjUg/N0t2xnZNNrRTDji2p9xSBRzqlOgz6DR89vUjKEBiKxtJK5XayJU0b2XrXeZJYqQvZ3JR82
H5BWk9QVBYnvd2TsfPr2QJySEfo3BDPZy3IFg+gzcWihAXVFJ3R2DCJGn1+n0Zq2Pot/b1R+FOSL
1EfKP4SgG+WiEXhU5uC35GmvKY+p+mkTuKPdLLmAqgrzDtkAxm5W1XNmKM2H+TRrBF0BTFso2SM+
EhV9DfhMVzYYcmCyt1bBWJrBxRWLW/bbKOYySYW7P6SHC9DbkC7piyGSvp927OyLYW75qKt8nO+h
UmeMNX6B44KTvt5ams+noTdgnmZKDC2oRNrABJ8eeCiD0Jqh9HGLFxeWl9wtf9qGEW3frsA2rGg7
vk+2118gtxoJYkh7l4qlbLkle+KU71Et8Ch0m6iOdrhTG07jaaOIyfAW6XlUrobZNz56ppiwsKra
jDrKJepXSxKeyl0LDss6NA0SkE4f49qHTlPy36WGJqiPi/nmJzuTkl89AaFdfPuUKyyC9Y6mOPaO
gTfOwgd4p0iTPr5drXzEsn028hUgMQHQN0i+uBPj2EMlfeuLv/+E0AuAndJWzc9nBbK0v28IbPzI
HM+zLFywReZVlGET/b0oeVXzvu6eL0kpAWpAuQH0Doeho5Q0nZgXidwBZeH4ps0rUc1tsk2cworl
I1cS6VFKnfEeIWK1NWktS5VZZU62ljzCD7Sep4yvwbRe/Uro/jb7tvQlSC+/8qG+AQJ6W+nHJvWv
g5fz7InAGek0B9NniTNeTc23CUwVoQeMr9GfVKBtUD3420zJysy/gOM3bZJ53BBRakSZCqi2jI8a
yVmSkZr20cdyy8xU8IbRi98fcs+GJzlKiLWEZ2jHkTULz0j7jRIHhi77qmUX+d9uErFbL9EMyf6e
usS8WB07XEE1oiAlSWyfIKeZBgEfVe7H4ObP6Qftl6mkkAXZPiPvGNvwXYhvVJcHRjRa8hlEESfG
QxUB6yBcdTBJZ6yvSGG288d6JFfG51aFUDv/LrgQNoMiaa2sHdMKqoZhWC1PnO5tDma4IaJ7jltz
XHt+w4Wf093iR8BZfOz5rbKeXqHuwPS/ujFhtQdMzmRPNqZQNknjnXQNHO7qJqqrONd2ndzafi10
+rJgFiBIM3x5paMtMyBzv3qRtYTq61llGJRIyx7M9PvaP07lEEjkerSQQlETql9HS8SdP3acR/Kz
QqQ9X7TzXMAv7AIMRAv4cLZVRfG+GbTKJhV/djCBzrkf7BrTX1UvsCgAiDI5/2FayIpl5N/mW8Ak
KN3a5Ov4WevgM2hl9eUGE2jmFWrc4w1xOEHqUEip60FpRQqf4KOA8Fs+fX4DzfptHA7OlfpfJ0SV
oyTh9RDd7LKwOt2Mc9TWHgpi0rg6wgBO5d1v6UyRZr+MBJ+r2h43SJjUdeGU55sAYVItOLMvPO/7
1tnYgBdbZEEQZIilcac8dDbnCJMdb4Y8UTzzO4tXPcTDBwvJI/La/tnct4ZxdRFFlBvv5j3CD2IU
17i0yVCe+VEqEyV+0U2cswV+vRaGYqclv3A4aieiRobxcO4ZS+kP3XayAOep6vkyK/mVg+BtLq0i
FqP0ZmcaqsyXb57GbVQEkvbXBfR5TnSB6ItCroX7JWEt0yEyugMAQpi0PAMx9w3jmOLRdZ3gepyl
9YZVeMQ4KEk/mI9LRncyojlAfYT0gStBW4PHUXkociRjCAzGARWoboFDuJ6BTdVYsNDZy71bZeCp
sNKXWOjc8+CTv4G7OTLE4wwMAp9pUQXyedE2dvPYvqGeEDPGJ1h/IiJ3OEqdvY+EuBJaUSslbQO+
i3CM3i9Zqy28SR4EvgP8TN0ylWiXTJ4cUvNDryrEZga0UyJ7tqwvML/HMLrJyOgLYQ0RPItdd5R/
FZay9DfiCS+m3PCdDawbmWabiYx3l7/yRg2tfhBtxMPjToNM8uBT43RIHxAEx1FKkHqvyD4W5nzK
K7NR55+sGHffi2LNhn+6U3rtaPlccflOyM07ew2Ep0WiwxVQj/aoHP0z6u+nUx+ozQvnUeCHgIrE
+AsK7T3wrDJcyrcO8oQq6iXJCXCrh9ufuPyf3d0urjTJj1coYo+d9+ltB57RoPC+tahymAjBENb8
A6OoLFh266WtAv43jwb7bLXU36E0q3XuW+79WrmdFLw3WZED7E8Vl34jKVCdVdgH+PnW6DA9t5p6
Dlp5qMXdM9BcHKn5ObzqleLOM2JX15UN9cqKC9IXND4+Wh+gFs5ARYfv2eWJC8weuqgwYK8yDJCq
UEtny2bpXY+shZtyUncKcqWMVn50hvFI30MhjUQnFFkTiv/P6jRFv788EDszau2Q83Ww0d9WO/PB
UPRbIhRZLqbcC5X3AclzCJ8N1Z9c6GNPxqlsfyDnfhnq/nruS2UBTTGhy07H7sUcQhgtqvkc9VxI
3cpO8YbSA9e8wplUzmV6w5kV/NviMgOwsFPk6vyYnC0xPdrFl2yNXsIDX+/76INOnoUaC1PTKwWe
ReUqx0DlP3RpFwzMJGNYcKO9SckzBTMpQ+SgRYuL0j7cVEZIpA0w737XICaSkcLdeiZy8N80twTo
oMb+Sw8cPyJnJVB3Lo6ivQ3jo605JIaamqp3tESmbG+BH/YbX7LQLf4h2LChHjBNLJU4pQPuIhzt
CJAxTuTbbZWArx1biW5+SdOYtRXfP7vHDVAAquQGyXdj+U3yLgu2aFcvcbkActawywlkFkY0s0WD
Z1PDEkrSrgN/7Y51p4oY+bSbRuI/Sluk/3dv+egkW2Gp1MrONciKAj3Pi32WMq38Bk3kg8vSsSF+
H+shm12V3W1V12cEIIFpaOzS7uon2ieH2gpTbvIFsMHep3T6xIzbU0jV/PK/lRsi3pQzUhdPEKjd
tkHvErLqX1OvXGe4EJKRrYg4YKZRGKg5Tr5fzTrsP3jpAHtHBmXMmULDW7mM9Yp0z1nu9o8nRRNh
YuRG2/0sVcUM3GD+ILnluyursobbDuV4kaklQ7/WhV+PE1V8ZjSIO9ym8Xo8CW6Mtck/hRfBXLED
N/mUHjmUil3A6vqAHMcIXyUweBa0u0Ld2oYJV977BxJvAnjp6eyKkcdYNYxdFRrlzWT/zbwZQ/JT
4GmTK3GxEvxyJYHBCRbyb+TfioijjptZqYBto/bEGohca3rOEPm5kIQfGV5xB5F+ZetdV8oHMI6P
Y22bRMfdOGqBwtaLUwU11+5ZgMyBlsvgknX7+iMzWI7xH3bqgy3tB0COML8y5icKJOkueVSDAV5K
aByO0kRBVj2BUFkYSiyCGIk3qrIgSkqlIfFsgRDqYTGTI4+r7Ca9mJ6nJRDrlDDlQZG9vNgIJOah
gCctvOA/Jynfc+OjoUpxqKUDH6yAgi+eIAb5R8cbWsL65jdFdsagQWbeNx3D30Io3U/mTeYTE/Xr
qJx80V52k68NY8t2xlovBUIK3I7AI5njSibyv8gj7+qrmBsVLorzkA9teLwGD2ISZnojJ46YMM2d
dTDhYbotuTQXmBqLVjftLcr6rhWcbPmMFLHRvaH1qxP53fsN+x7HN2Zew4+UCWaSfo/y/6xSTklF
6N38u/7Y0c3vliKKkhmalC4po2VmgY6HYYZEzdSm6OoMauoxe60OmV+7Sde9QiyxPD3M2U7F2Fx8
6CvqE3EdX437yn2+qXFNcQi5S6/FJeCg7oYAD8J1rGxS7pwYfSeIoMovfXu+QyOy+SbK8xvVIHmM
LCZeCsRk0LXRKUBwUHQETrgbh6qaWf7hkT4TVn/P3ymw8Kxi4ga1XbuV7XegjR5ZOs+kHFbFOA4E
CnjOSmMujbfFoFrBNgKmusE7c+O2nIsh2sKFHCZt00eo0qZ9vkwz9VL1hPtjhJWIyp+8HKk9yaDK
PLeLA7MtAm55+710cIZRJoppXL2SL279oJNfPtdAW3cGgdMQJEZVEZ9mGPSyOz9nxhmPcbxk1hq1
jPzsUWAWvqetHsB72PA1L9r4tuR5WFDF0onl7E1RJN8gGNctqb6U/q70EvWL+mfKQxz4zSwlLTQa
9P5jIW0AGDou5cfLpwK/5gRc/7TDYA5o7fV2/qYwx82628VXzifGcaXHSRxWTFBO6bomQz5V2VCA
WAXtqvW/iS5wg1iob+XAHavl3N3EdhJLd5JyMiTIGSZt5UgirhnBVMvFh78o3A61s1sQl/5gjor2
M4FR3y4ZumzSj/U+e7Ii6fTWp9O3/qFnDD3zYms1eRbzdXWsYC0SKWjk9V86U6Y/+6A/BaQm1OIE
W2OPqLyjsf4fiRJ/3oiqQQ/qJm3IElk4Y5phlB9nhTSSe+jhB3vvweLZRjH+T0gsJsJXyX7v4ZX1
SWJ2Yy5LpZOHTZOcM3s7PvJbqfuypNJr842+qigow46iMkBOVB+VR3eWdUagDvH6wSDcAW3U1ruU
YNm3Ih7wA64I3nSMm06K+JtcEPybCsSesnHC8skPhRW6oZVLGCmgOUNgfJht+3wbDwC6r78qcnGk
TXUxmkVOaAPSs0VfXYKjNUW4I5NJfRijce0XISdTjTS6FWlZ+aniYUrIoVATqbwnPNWQiFAi/J53
BzaW0Jcq5UeqzAQeMC56l69SNbnIzheruC65dxx6eFRhUwkSmBuVIxlo/tz95k6gnfOgnqNy6WTh
IGsdIJ0yc4Wm3RDQHqoae0gYZheKP2sEZ21+LGUrFB2nSYWWKSKMTGamx091+Kyqnzdn/eftdOdK
/yBx0iWQFxW6A9lT6EruWuzL013D3coA7oKCJVV/WTqqts5eU4/jt9HffrT+pc71idm41+mMnBfi
qr5ZyhtzXTZr6tyre3FF19W81+l7AkKEFPNsANxDaDFHoKHSZwBWOvnXB3aZECzFPtPmiwVxLods
W25BnqEbjqKZ1duKAdRQLJwxD7g/9LjYolHcx5pSN6/3sanUWy74LccAeW2OaMFg8VvvLZ+eZb8w
An7vYd6pcZgMh4obv+eE8H4bD2Zh0sl6Y6Z0a+a9hMnEJ1qHxpiHwcMAHGVnRECDbcTyH0+kDKt7
mOUs0JKeAsZgnmkuMhw+Z97x6OOxthV5xyIhWAC5ZuKTAW0HKxMI/KnVHZe1MeewmRLGWFjZNODZ
ghNMkmVcZ+13txtJwHqkQF0gV9cNlacUK0HUUo+Yqgy0uYYIN8vwD9N+ERUrhRfpAjmYUFQHAHHl
OwIkpRAsIh0BSkAUnAFpQLtEDHpEYgrL2W2kw6B6bu1oVJ1MpPpJ2iXaVIi0rZYrim+VbePIKo7d
97X7WlQK/d445F6TBH/UCFhINxlKng+Syw/D0Vb91FMIt2WTKcFVU+dBKKdzmgy+JKrf48lPI/TP
OFsyJx9XnXQWI8dzDAE0fxe3Rck++HldOZKWgisOwCNVGDkS349AdPSbL+Z8aPDLwRiZ/c6JPTfD
DOYSkU5CKREd/qSOXTtI1PUGYUNzhEYwqT1+YHnQLCLO5oG8zSBVXnkb77EB7VWQrvt02s5hys1c
p/xhklQ3tzYOqWMT+wdMCF4WWQMEC1p7U87pWVhvDhY00RmyzPtIpozGeu4bma7l+faQ9pY/BGz5
zEkVqruczMIntXNR1p+PdA+Ti0eeDx+Ig0GyqcFjz4wJ/LoTuQ3pKNKNOEPelh5FO8ZKLcvKv4Mb
uaAkDW4//daJOtZ07zkzL6WaEbhPIU2SMKLahtgmfsCJxQEICpCA/Jdw2DkXbZAogkdi82nodGAU
BJzO4asP6n7vs1Svc613dWagYzt/toLVStpMArp3CuYxh2kEnYOW05dGTCNiNog2I5yShdxdcoK6
WbVIQGt8wNp1SY7Z2X3UN2oFImC62e6i4tnRpxh1UOS0yoXzgXcr9YfrtnukNQZyWWT+9ml/Dm83
It0Qpsk/ZxDdwrVQOJNQsS1Om2kPg9zi244T9dBebS47aKaP0G4dsBjIM6sMj0n0ejPrRf8TzAe2
Bo68FoxdLKth0V2MbHNZKRYJcNoUj2ZwyDYAaIRTNuBlXrwDdUGVdolo2qXo0B27hsz1uvu/jjWR
v2XHCSqCHDmF414sj2WdiXDcoAC24rJGgLzbzhXz3BvucLizYrvmrVjJMFWt1HgDjJTunPnj1udS
R8fKJZ+lstwFXs1e9lBsZ+xe6HEcECvdyyAWpHzfjcbxBFBqVO4CxbckOl6Puit50Mc0ULXgoJoZ
U77jpWYL+ihdyJOh1nvD3KnoclNGEbTJyHeMkgIu/mjHa8k5b2W+M18Jloku9niihdi/X4mWsP4W
/GoyiRC7fNm/KaGdB42RbR6J8BBx9mw0uRxq2/DxcUEmtGspqyTxe4Ka9Fa9wMrBuxV+sxAGjiiR
44kf6tRBdzMmCaEVYI1p7ohUWEuUJPovJTCfrXoL7kK+YzCt55eUwkSNdUULCwDEn5ehySL+rhXH
sHAAsWbrJQKG51KWblGUO/40h2sZHCgL92MqQ8Jqbu8qM8ErWzZs5ZpQOgH+GoZBEdoQ+CiOTbq9
Q3gWmVjp81orZ3ctvD9gFyZrnIwBroW26bRdEx8u4YYpZ56ccrArr6DQvOIy1exe8Cht/N57Ws+N
J/Fl3Mx9LAfKdTjY4CHMsDa91+xadWivlJ9E1qf/7H10yXGqcdc4LIL1wEBh2/IpDKNuhuk+Ix+7
us68dKbXV+B+VHEDGH0ITuH8pvTFakFHboR9SqNtRU0RRQU/JWlFlQ7eDefDvnuo9nTL1I3eKLJr
IOrI3yP0iJOC+zlrYzPbCGle8nU00/y0APPSBdbNBZNU5bytNiRRGweaY6QqcXcfMGTHGVYyXzVt
JLhNctYCfNJImcqQBpiokbD9JiG0fPUF0vVpzEc5+ouDCO7pcf21hXW700iKflb6Gn4lEPckvxzI
+2h+hmgN4yc/SkUVWPhgAAuTjYAoCCLvWoiTiIdGrRFDhfMuzcuKxjbirbSJsORiB8pb4zlaRWlb
mqUvLWmPghhnZIO2w3FJm473EWoPQuDtWHtp1Ip4pmmNJcGo+oOIq+oiaHQGVS8c6pSq0bfmLPmr
Ie6GLLz9bVb036cQa/nMsv9xxg0d8QxkYvMy2KPuIOeWVXIqyW6trIVbDkyl7wpPumiavfLkQLCN
spaGwmYf5G9CWkf0xNyyHyDAkCtKk2JsBJNDs8qz6l+uF3htoqSqm1cGS9Z0dRmKL6YEl6MXAZT+
+QZTh4jIrcWi0+nGAsaOdTTbAAxiV2PpN3eQ3acysaMtHU4vtl9EXRHpcDKsFDpF3f6Z7Uxp6Ivu
pGA55oMlXm970HdI4fx/uTWJgBhRMio6NCzu/BaUTtWmaZzg04MC0Ja7+AjTWt/BFnInso0/q5nA
a9VR8v7U/BAlL/CVTB6uIBlhVnPfTHCPwXM/ivIzGmf35FZlvff1wuV8HJ/rG11HfJRyAp5wKGwh
/ETdzEgJ1bqk6iIg5/oXMtcC1Zg3aDaLD7I+8jpx1OpKl74MC9KsPJwZju3PLVBwJg6ysRF7s8uH
RGLrRjbnKrhOvZnE/MthT4zOsJfoxdkiNqgWLQrsWt3qD54XT8fIU+gn4XkuWDKKv3XECyd/WE62
xWzbu1THV7+bxG+ZrbXFyHVvLwzhYVFo4pWFKfwQhiHx0OmktxdgU7RAeVx4ow8v9WI9np7Q2oHK
j4R8VDFuJIp5zjuOrX8X5KVJ5RELneJqWtRosxDOqGfO+1GLSKTcoCwiLJWGzvH1E66eBPAEe1VV
V+jKAromn3lQWPmeAhdKr/aCnx7jQP79++/ViN6lturN3kzsI1ptSZvC6TFMnb2BJqEjj95lTu8l
N77Us1Otc3JLV9EuqnSovAydJ3nGLXlqu8BYuOT8d7DxPlTC+HyTTUCtRVvSJEFzEZe5efC4gIMp
IDn7faVxh/QYaD6TdvvYlbu2i5Rn64AVsU9YGVziXHuwLhEof29lL07CGhz5l10XEMGrpm9+Y92H
e16XbFOJE5ZMN3RG45qKYwsXAPhFKH4sX0nNWGYDW1tCB2FPg41ilCG7wJO2XNTg1h/LVbFjzAW/
jsJvkeIwLAtyxk9j6/Sp/IeUs+9EXm/+6gd8Xr+E9tL/uF56Bb2IWmROborDXrWpAvHteOYF3iOI
OIKiSsFyk3/ugdgrraHyHtwjzijnLsUKZz49Wt0iRq9qXd0eozUrAzcgSPhuUWrqpeZGwa7MQJ+a
39V2X3CB6hUpfyFffP3nhMssBZ56ofE3fgtYuc0//ImGCZPHuW7bmgTrPQ8npY6edxUc2hZJbVvt
tM/U0zxZnEjycQctTAzDHR7W3bbg+PFZyBwSt1JAF8vvGHvnGSKQpT6VGqK0TQL27IjJk1hXyEh8
jjciH59DwGUlOBYFvK18ELbvHE64lD9LWL8W2VmUE4My3UigGfB0ZZo3Yi5AxNc1PLEQZZvmdvza
azSkAimScmDY1zuYu+9AtNUffR6mGHWtXT5DsXM9UoEqQ58Lt2aGC5yVBpr0tX/tnOvIXqWoxL15
25HmrWDZXdBjZbI+vwI3FdFy4OL4hibwQOLn1Om7sDTXHCz0iZVVK/UsUtE2UV8vUrh9qPGFPaCh
24Ty0MCbQ1Aw2yQC/oiUf8QUz2n0lesQhkknsLdZP/Tc9dTVQ+k4NwcWo9qgwdESq+ata0lLQBdo
RzJ3e+ioOcOfJjfzOdv1gVCMq6csP0YpI7RpAPuS9XW0kvykwKPHCzPJCjEuQa3eE6cqZ181Qngv
Pe70e6sg0UsY5TL909ZTbyfLZaiRKoeAbEC/N3RjYPoXRW2bMsS6/mRMahy30S3rB315GVry+HWK
I5W2RZnHXHP4lNxaVbdlkijWsRtFR3MZ8Gb0xumY3E9/loNRjzZlUCnbXgY+PxtwxW7S761A7e3Y
Gkh4A1RA6lsHOopl9bP5qfr/FQnYkJDV+dSx3ZXL/z7VIWJCsao95lpL9htjVDsza5AEFjPyaZOf
eSv7FlVnLe1lVFsmVY80JO18j0HS71IhlLfflWb6TQ8vLGribHbkVgA9ueJZE4YUsURaGU3koSIz
IKlkZaVy58IAjLjfuIMI/zrbYblm8+SUNuPMISbSL80ydmRCz/rXoS0WCM8RBsEK0Mh8cdZK0hk/
QRAFHbsI/aRYNzbKixpY640vB6/nFVh1Qyc1C7cb8y0ycNhlEkV9Qcd9iKE/QeEozs348ehWDi9r
K22lVm/0Wf8qOLt77P+b2qieVJhHpZDu4obZLjj0lk/eMbw8zmCa3115gC0kpfogInOlhsyWuCjR
trGkzlnXzooF7I7/dPI95j5T6Cj/mNc1l12O298m9zRS+kjKgMThVhfblRxJRexb65+cacUdudY1
sXpoGZQY1vbspEeVQx/sfxnuVJ1ECwJLyp0Vi0lgTUsTmuVJxNb8m3u8cirkUL4Y/Rmx8UHDC2/4
lHJO5egRy72f1g2Z9rYRYhZ+v8BAmp0uxLTMYXaY8JmS0dqI8pqc7FmL7SOZHB7jQXNEsxDZgly6
d+VHAGne8zDR+c5Y5/jSCrBgqZp9exWOAxux+M90LumIzI33k+ynki5ii594s1c1nS6zf1XKXpJC
/VhjeAxN7w4IMkO8JXjkY/UjRj18dX3YgbUnKMvNPXhZfMWsQK9VnTPw+6UR4/nbUz7dpTw9tevd
rkpCdsPWSfYrW5iHP+jHiPH440rOiZyS8MCJLXA24FAKEJ8++xDM2QcNWPM9ioi3bMEoGmL15UCQ
x3BebgaFQF1yeDiZN93sE72rKT3qnV1B+xolGUnQbCq3SqZKR1SK9NM/BXrcJFvDTwAmiHhp5HYk
rcmP7lppvlWdPSuZpyM+RTP0gSL1/0lxk5gZu8WxGXUg2kxQz+veswbymxeUg6ZzLw+LJgzl6otE
/8d3v8ttBLTzHhIVr5iWQHMYzAg5Ow+1/PjAiLHR0IsQ0fs+Y17dMt08FwiGGXE7iSibIylFslQg
jBofwujqMV2AYQ52+KjMJ9Ls2eNUgJMvODDAtd5Yz12kkqTiPx3qO+ubsXap/f1xv+0y7w0E7mwv
vYWPsPdzAaZvZQ0Np4uv4EKeZprmPJBE6E4gibV0Ea5YiGnQqelh5ZGq0DdaGxoqiWuuOQUPaYiy
kKLMwgNOVAaw7ST+w9X9bwu/YnDLSkNW6g4jafo6O6m8DioW0RvLOBjTQyxMj/zXf3UOzj74pSsH
E8fDgftZTTRkT3C/vNJcI8dz6ysrsnYWa+8D5MSP6Yg8meWcSTTEky+Sgg+OdW3gVmPVM372+3wJ
gfFk2o1cREuBGG31cE/wZS4LjMkEvNBpG0VUuJdYZBVNBqYPkZv8hrX3XjinavMjccq+SkdjT1dE
D1xvJ5TlVr0RphmsOgE5+TO64JJ/WtXR+FSQqNUeWDnEREBzci4h+plgIZr3MinQb8D3ImMBH76n
WivNIKPROMj0PvLvRMEaBWiZK8irRdccBYUOT1QgMQyH9H2CdL9S9aCmmV6oDgZURE39cadTTGkw
ugi5xm95+zY5bQdpv8DLlBqMT6SQSzVlB1zm2L9bYpEHGvWUhK0c1/WF5RTvD0nTclrmA4daEU/v
/wRNpF8tSy6wHhI0aByoh4qmCartRryewCpV6saIyVqWs9mGl4NdZ4v6kOY0K/da/7Bz3Z6GgfYV
MR695eLQLI4zAxWsQwhhfJpo6JR8u5FpDqNq6cXv6H/B9kY2fhe0EFC0YUa8QQacITySAuqEujqm
R3968ntNAxwBW4/XkWspfVeLLArcYSxa/rupMbMjMuxdZeGhAUqcrcjq/9KeJhbRsQVRWQJFB+2l
riJv7oB+GgVJ3kA5x5fux2vlJ5oYkMUynvBb+C2iCnjXEsDIdeFM/OE19VNevhMaz1Vol0jbYKkW
J/oFfVmEq+OI6FFTzopRdj2UCngIa0qbwCj8poCiognNGbephEDIbAfRVce6YcHuNTkfxdt40hH/
2kn8CqaB2NCiopKppV039nMPK8m9vKpdaOSjjTeUSpvAKcPpOKLMbmbbWm9z42VcwkxkzJUykt32
AXLl2A8QcaZHuVJqhQ2VOw4l/CcvK3Y+2vhi6H1W2wuY0bj+a/URHxZCu/xJDS/TK0s9ZbjEInN1
Uhuun00+rwDvtDrJMI+F6nVsQch7dXNJw9D52MuVauLwlm3XXvJgs6VqRJrrQSJYDg/zVjooHVS9
/VXoKremJKqV/TTdMQCkMuR4h9Iww+WkEfg0RjJhNjjNCFqoQK40ETnLaKBPJKDw66v5SF/Lq/t3
WxrUFBNvYTN4XkfVI/nLb/Cs5/IRGfKPrWvvPvjZHw6+gHV2nghnrhhNK1DWScPEIidFSPNKEpa5
yyMDwqAxboAPOPQYAg+7HolddY8MzjJfXb/YOknhRZl3C6DCAFhvQM+JMNRHhNXVeVvFWOgY1Jhz
xOsnP1lwdFW8vpI/2AMhGtr5KtAd+myOSOjCLu1Rs5oHHhg6dxtXYBNoZMqyRqMhU2yp9x2+7ZnY
RLyt7scWma5IiZWhWx0H9/LoxKkB56e9WyKGu0qtNLYvYxaxcd/hdN2lzR1ULEFyVzqqCJxfPRry
h0qQM5rrp8DYP2IqRQMktUBSRvr8zwFPR83wGME+qjswRFp1qRzAFc7d6OT/Uij2Zm/8fdrO4f7d
o9S8yDZ9V3oLg+4bjzYzc1ElpezVQMDcwrcpo8mlKchB5mAtWj845PKYIlmqj1uLNQAnOklqJTSG
zpMUUWo4QYFu2fdhigs7VsB6HXFqkd+8AhPrbuTTkmDYeXf9PYQqVKa2PSNIpYjpUr/InekkjcH9
XYF6ZLBzoJpmAz0oIA9uEC+rii8WBC9cDYk1Lx2JoerWM0V+RATsZRdyHVM7qmKiEyypdQyVthqt
nz7XFBlFi56iIqjg/qI4iIqwiI3KpkgqvdeWHAnUGdxECFX/Zchdup16Av6KWCcMBrnn9lbR0he/
Uj9drij2lfAHUPI8TMOLAB8npzx/KxmuskfJ+1vJGDqc0fvee4BAerXm4nnBySL0mVMeQPqBEKNb
XwI33oyg6eqFwZzGvC0ShRVkS1TxZ/Z7zi6USP5f/QftPg+F72+7koJgp9BAFLiCCt3pkc+kZV1g
iJz5EEKLwwzWHMRV/Zis4Vq4jrtVzX/mHJllHLwvtJYhcYJPE/0QWoqn4xKytAAmaTlXcdekP6sI
kddpTby2Z+6QvgLY4GIA4QV3vCecUSzq9/H4MqKZ5df/ec7IJ7t3CkoJZVTCKeetmtfW/J4UEUr+
Wp1c8TpNhUvKhfLUcNwgqepMmMsZhhfaNYTlgm0rYy3ZGkHg0zd0C+npptnVqOw5HEyXj5ehmj63
973IYcvyLUgR8l7p2fzQfT/3Osa8udLRCq/ruQxY97JtC5DPfBsBxTnEDXl+epaCfP04S1C0xiMZ
H1zHjv1lDbAymdoMQ1XtEbvTfozq6aCkA5KZXnFs7KsWq8gtAaEqWtcgOzmRR7BGi66UpN7+CjJF
i560LC3BTrAVKrkovvHRodzwW2hV01EAGXtPRiy6XLpueLT60Cd5lbRLxOsB55iLBahxS/LD8hAX
Vh7z+u4Oy/j4aoOcO0ALkfuQtNyL1xCs/Zhoof0pMsukxyC8CTN8Ove7qh0VeS3gf9mu3dRxO2Vn
vzVpW2ru5p4pv0BmEq4/qP12mRslZrTL8MPqHclu/93aJh1Xqundpuoee/Y9SUYyF+v6rd4Ez9GX
ECeMJ8MLLWqfoy3own1nDEL/iWUNQ93/PwF7O3m63IX6JKZ43wDnMLOY84kR8MsEA87jhA4gQBBg
2AI1ENI5RIo/GhRrBoi1MyaD5hyF+ki286/pPaIp2NSaWKzSRfRTIlwDU3nuZi9SDVUQ+LfzmPbT
v/QPz29cNZk/vJTzLvS3T4GwfNAJ42Ge9tI+TObiV6yab8EHlQh6JTkY5jMmXfx3Mv2zYpmtTmKA
6EumCRJ/XleEtCbPfmNrEbsNqI527RayHUb9Z0UF3IbfFzApAI1g3yAp4iQle2iRZb/pbTCvPxJf
v/RupoUTqX1K53C/mlBKNxTXV1P4DOlWO4H5dDo+WqYj0N+439IE3yQU0Q7hTIqsyU02876DluvR
MQ257ASfyfujtjsbAi3iyvQMLsvXKZ9ZTDfCC1cisFwz5qMvly5phetcVbj7mIXLmMrGE7661tuG
4jW0+g8htU4fzcd5EWnK0Ej2T8tU7hPagHoXEsvVWl4UBmSeFhinYb9zu81aQSOImDKTDH+KLBwz
H1BV0CfBhBxw3jVeA2AlnBa4Jd4Mtc4xuZ8gAJLzQFbOrB43k8C7OnB3lc7oUwi947kBO8SqXrFZ
taeHid9lpjL4upNkv63bVxOdEYdyxExDPOXYwEBTNI+NphfdSwuKxY2+0TsDw0jHvvQfnwLkxniQ
bZkJHeTUGABZcaZtqjEK9rfxWA4XsWy2CbPeBk1aXdBEZTi4Sy0EOCGIBO4DTVLyWy0rU3P0qa2+
2EdivzHh9HTIsWJ6FSJZLOt5CQCXzMTtCw7myILIkvoMeHkF6PdpuoVmCGZcQ9uTw4UTXXWEm3y4
SL/52HBNcszIp2N1G9tq7KinlwK06BhHrBKrtn9ruj5OniBsIxxXHtDaUWrHtrqq0JGyIom7sWwe
gPVSKQP2Xlv9hV53PObsjJQqmAl4xM16f4YlBp/LnC047H+CUnOAxfsfWACWYKheyQpgNvFvBQrI
KFm7zM1gFSh2QElvXFEPhL2kMUfAIgo65GOAw0mtyaTAydWclU+HcAy9eBaEzCXMjEYUQTb/EmgL
y4dZc8aIbv3U7Kfac/Y5qVuoAvmEjnJrSSA/9ntZsXfgtbu9yjOzsY+fQoEqx4sfkLasyJ7Fa27t
6UmL9LDcHFH5YGF/0YFN+tQt8STzOdIMzzGsXatMzPVz2Be8AjRq0DY2q/8MMoEsvbVKRRUD8VwM
viB+PIuW2CqJ5IfjxAh5px/+v4p0urZ54ehxekDWxSuADscGx/mem5gilJe5SIrj1UAGQR4b8NDZ
yhoFxOjdoTwOPaVnrdMwHpWn3K/0tqUrj+3K+gDRIOEXr4kuFpTx7oaptyNS5gxyCrB/GLnmop9/
WsW/pOMdJt/k4FsqTAdgId+5Mes4BpYD0Tf4PGcPd6qq6Sx/ZuAz0tGj9C4ZH/FuUzGG8pfEbmLl
3dYC1TZFJiUFkKEfly2g8qpNSjzn7y/gB4PyfGHJ3jB/eYBK4e4PIpepimDe8aW22LVBz+BRpZGW
3kgGsjRA3fKw5lfQBGNNhuE7c7O2BcSwLui7dhK2BTkxaIcM5DiWnd+NIGM34g3NVc1qjKp3fzw9
zy5XehbopKfpPA2M94m8P1bQXvcTurm4NjLUeWORVXkuX9isZsCBceL/Xka8wUO48/pEuUj+9zME
hX1DiRO68yAUDs/ucg9x7VdCx2+HsAtM2GXSTmrYAE5pEIphoN8qKLxDWcRRlDYJXmPy6df+QOrs
VIYrcVa/wBe/OEwpTfqf1JwyhTtUPnoBeILQr9ZilwteuQeohJXJb+6Jz+9lj6XPLdj7P4wwXUhW
nGLBII5L4s+Yfsg4k/bcZlpj9A98CQaDTq86dig68ApYlMOVDzb2OwglzNOM8gTeEXwruCAM9Axp
o/bb32/J9NWoH8rudbDZk+4t52YzcQqzEpcUyxOBm3wmBbKZyv15Tc030phBhw5vuX9xELWbjqSO
ov8Zm+x35QjeZZB7+zVo9MHopOnIApDVmHYnmngsl9T51Cp6Uup5Dh93cLpQp3m3yaJn+Zxjk9dT
VAYE4ph74dv6VK6WUJPB37PFLPVlPe/56NNZ/P951zziV7q/0rczoAJO0QhZoxS2xZgw3ciUxgg7
4zRFpAR6SR3Od8XtTvamroy0fYmEBf9yo4HgnYqKhP5tVyiXGGlPs/7gZBCZKzPCCdH+yI017mIQ
ZRi9frHT3Z+F8SNT14grdX4g+J3XbVdKPO+MKvLTJogUlLAH1Za0i7lqUyTH85/uLxNHU0UIhqdJ
McR5OSaCFSXdYSSAlKBEQaNFVmcVm2EmvkJEoVZFNSz301uJ8U4ITjxwfMBPOLLXbgqdn7Cy4X6N
zvVAYQmYjZiz2q/g6pR79i9oiOxwz7sBsXooO4+QjGNx3uNsCQmWt8cq5f3z/yKdWISbNMULywM7
CYCyVL5zJbuYa5tZ847pDkNG3JYxHOXGPK9Gqp+nZlS7CC1J+6D8wqpfY/YXLz0q8J2uXDQHYmgn
2ANCdWe3nJluLoadeiKAMlZk6R+UtZjajM7wAhtLXdRACWEkNc8CUUA5bYiIutkDX9QAFHQKpory
12kgAL0xnKOp2KMGb3N7cybVEikA8dhS7SpKEjgFF8cF5CJMf3mNLUVVXp8cd32Ffuymr/JCIOQK
SHIp/OnMj2XQHKrmI4MIvZngB6iJKqaRuuDOmoZ/jVZfVZAGMbdb+Fzp9xFe3ys1gCiWt+APHtAA
HwpbLHX8Pqlmyhjh/pXjuNVtf+qnQ1UpI+T+FsxSoY1GRDdbvqLKerzADqTey6Husz88BgQwshij
SN/ntPNuoSMU0dV7dYEaJoLhZ37AmiBXkDqcnwJEVxuf339WuyfauCSNISyNHbzVsReU/BkkKJgu
fCBWl04pSg9IpaCQSwlazNeUCgK3LEOeUkGGWabszHSOtyPqtbFnxs1yMg+qWHZoz0DSShJDZmQG
XtZrmVjno5f5ZA4wInDEoIAfQzzV+o6CAdM5/XaefVSFqPjCqn0c2yEK8Fi4V7RoyF0nYDC/OQCV
DOZLsLjOPFRfJG9qQcv8XaInziI96oA9hJUTovEEcm9/EnG5iGrwF6MzH2IsyNth+8pUFbHqmUZV
grvKpp0+uQrpZ44eaQwy1auSzZwyXSWqUOvViSvEQA46ykiwY4oUKul5ylCn7k2NwDbWH2+nwCAD
Rymwav6JOown2VangJfWQQLo/8GPL86H4GumeMhBiAMr3Mmm+s8UI8iqKnSWQsHA/E8MAU11XWXt
XHtnbPjyPGwCtd1PXB8EI+bkixBUqM6/mwMj0t0TfNbALJK/zEkacy0pidLT66W7TeHjNZ5A3j1e
drJur6uw+DYUuAeM/ekk9VbZFRF9yAnamj1w/1xVcHPcJnGYkG5dPx4N6jHaX/jqE9skOyu8xRqJ
CYoVnAqyInxNlcwOpjDWI3FoZpj5JIfBjxiaikMrzlW60SQ/sKMonNcodTYq/jfy+NVIYRqFMZO0
giLBnNOXPBSDkfu3SRVSUGWtOoHOB2R5hE0F7JHvy3zG8wT3A12L30cI11vJDtYwAFNR0+NGmZoR
5EYQWp42QPpc8QfFPsftr9gclmaeGx4/89PVAUraIyb5u1oI2dw+kCNzlIqn14dCgO/2029VSm/U
nw1WXqx6kUY/6cDYP4OcsiztIT72HWshoJKsVZva/nM5YV/pNX4jFGSfWhplv/goPElutLE7Maxd
qS6vlgRS+PgC3YEDbYWOPKt6XiTD5QSW5/RgTVV7qlZezuIbH0Ss6cmO8twLUOMQqmcLNl2F6gHk
KpuLCpp5qelbzNJQ2xniQznUmHQymn+qNoVgP242R3S2L8vh/7mDVkGMRrd2YYSW2MTuNYG6tE0V
Q/31PgU44+eVKsZekL/fgXU083IE5dcsWeHDifH77fkVv1y4h+QbB7OFnW6Ge0ZV19tPJWgy9FGy
bjfp0LhvEwh0kP/SoZ4srn6a0fAgNlDG/wfUWcZBBBwO2D3TOYVVPUzTFcTDwHrYpbkTswifE6ZY
9Liu8mjLhxXR9dzVDMg5pgNvED29ewIC2jqkOQ4KPto3eaNJ6Kb4pqxoQj1SG/PHmgw2yCWK6mtx
WmThxqcfnMm7/+M7JK57JO7WMKlcDNaulgkOGhEr1LH2V9UuG4TOr7LHBHsThhqnRMwQfflzza75
+r8dLIS3DAysUqAjVOothoz9AjmoXodw2H4+SIeEjGTAw7rDh9pNzYPULFLiRQNni12NBEFQ6gbX
dhTMgrWXRH8H+O9YuyuWMcmB9YISXPWJo6kOnYnKH/vuiL8Z/oMNYzGOpOqX09lPsSU1lhDzNbWp
06Xh9L8LREqLYOaxtYNwwaR4nqhkscblLvBTMOB/ltNld2F2PIuIrgZb9rsufBPwjfQ+wtLNc+AV
e3IvLv5ffroTBY9kyNwSz4IPKTQ4C/ORTZy/EjF/byOZNv1g9jsmfEBxFMxd9voXdYa1kjikpl6o
jhbf4CSF9xaAqk0jsuYQli86MR+OeIFGzn9r2zvMYU60I62eDOYPxeXTgAVGA4apGISLIeTbuX5F
qYX/9U8hw+TXTaNT9BQ5f+88nQrj+lk/jlWqnPNTJljKzeWKXu8+eKm8D4kJhr/3LojKTvgF0VFN
3pX+WJ2Yhz1QtfVGbsbSsx7UvE6Tz1T6VLJuOoIWzVkla1gO2zZk2vzMjFrjQiV+J40p4C5X3mgR
n4VyETy7MAmHdgejZxTvBgb0DQ8hz1PtuysuTKZbr7Ubx9XI+GbMM7LckghmYkr8Rosf8i+A1PAg
Kq5cbAr8rODK66qL2P3tHGApByk2obO5d+vd96YSqwLakX/9RmZT6QlJ2xoR/vLbG7lLCpOY277Z
npyovzsd6W6UdvTLSvFuZZbvC7sSeqdUTietA/gIV7FK5Y9JxFcTrPPFbOFIkLLqT0g5I+0Yw5kX
6puLBryt3bsju2I3/mHcP/y4KWyDiWti9BDoaR9+AW4zmZ7ELnAOkrGpy3CJHxkrSDrgzk8Whu5k
X+g+QpYg9KPv+wPNjFOT/GMmHNUPSf8iCQKk60Jin+788W4xh0Cw62tVvfyUOuYXa9+sPXchSB6T
MJMOw48eP9x2/XmqjxyISEZO25wuWxgcIigurkNa+013iP39Ar+MQ1mz+Ppas6olyp7FltsnRVRt
3YUNB3Svmn+YeMCvrzmbti/lgVi5yAoqlbdhsjbG5FAaDW+xtVVbNTQwTbjD6R5ibYV1uvaMRcUd
d3fx0S8BZfvTD8tDmipbvwYmVriMUr+x8QLMZCysDGoJ4etGJ/Y6TSFZZXUKa//vC0jPaXkEbSsA
VBYc8tOOyPBmRQIFJJfv41N0clbD1QH5GTSxX6eGz/srKpFyIFisPwkFKqDEwCadtF/rC9RknkZz
aDma6CsVHv1IjWgyryru8q4XSPipO4gjmyOF4Zg9GzjdQy9y0AuCTKYippTKBk1j2rmBMsrDwtqY
tQFDi8Yf07yx35Y/lqn/1yzKbrzA1f69gZcT4hlY2yUujx4YHzA+arQrGFJ7e0GuuRrwbB80OtVR
i1pseV8b6BmDVKqx2DDR6yn+adaaEQkd2lck5YPtHko8H6lBQ4bli0tyt/iUudCRBG6zo2VX51zH
9z4U2gB30kitg8awaUtz0WGgiQRmpgwbGnVo5rlAyqbLIYU/QKz1/BRKEcKpzUaS/fnrc4hXu4+u
rJfoOoEXmMzfWp7nNy2Dgbx3I2eSlp4YhCF9LhATDprTp2jYE+wETNlam1uKSi2+ErBGDW1JQHvG
lAwYU+rUVhp106ziSnRDjPttU+fJVPq+LU+iWoietMBuMCiTBYEw2Fg7CEJINqFcvbzb1llfj30p
SreERU7M8pt/tb6nv+W5LTfZUCR0ONojDMpxNV/mLtl8f3qpBEk47jmUvXIaYZOBt7iP41ttpwPT
se3udogt+z/edQxIIlLsdX2xbPZ7o2rvnM9Dvqdkk/NC5Pplha9kyG6v109585fTEKNgWx64NRQ1
YRuFSJKw1lvlns/Ex2xlpYGrbHamTasG7dnzE1VEBS31CLMCvvZLa/l+iSBLrIPNEy0bTUdD0BPs
jARVL0K/NHI2mrjX00rJNXEbCu8GZz0CplCl2NA1fct/9nViMMw9RnD2QQOt5x0xWPftsi3YnYXy
ptdMffW400rrht/1wMUvAABDxBeqiwPMC4JNXPkDnhqZIU5DcacqCRVWJM6T0j8Uso0GeGlboLDL
NEERA4ivWvho8lo5gM7IyTrNm6NGB0FzqISjtuAEwh+wpzta4IvAx8mgdVEM8osCDjs0k4VFuFr+
xerxXK50Su/DRr+CBDcF2RWUmjf+zJnAL/dAtGAO3mcnmyoGXfPNimFNF2by4muQK5VvoRD3UXQ1
Gz/pGXUf5dWu4djq22DW95UIvgA15TcROi94NtbjJYgL+/XC07CxZDeaH8eSOUxYnw/K3speJFOq
MK62rJ7mq+kFT+1sMjXmu2VCPVVAsKWJ2XgigQ/AETMqML7shHqitBAOSNfE6J49fy5CB9bWM6jt
U6mayzVRo4IgowaTNvqOr9ESZNRXAo23PtubOuh6Fo1Ak3pjf6bDW7ctBR2uXws1UWOb0D+XyeNa
ny15h1jLuJmB1cxSVJuK9SSCPpTEQ/YZiDcPJW4v8b32biVe7CG8Bq0fLhMFHjRYDQAWrCXxGu/W
B+cffCBTPcguns2zbuhgq6epDkQt+c9PeJItp3lvCEw5mvYMcEn5FAmZ4MSlLwAiytZMkJHfBoTi
VxsSC+OsO6FuGAFNmi3vk8eHy3HlXzujPgTEWuLcGwgQyV55OpJFqymMJPAR1qAzvNqK4lMI+kRI
KtNdf7wRkE2aRscgaqjwQUiDFA/EMQ5wuuOrnH1gnqXNh1AxZV9nloI4b+BXMI1vkxaaf8c6oGd0
cShQa18yIIKaVEcNxTq0ZXT57ujVeoiq50wwjvutNXA/l4sa4TI4D+SxkfqQiNJ5S6Xs7TjNtSM1
YKNevP1OOeyO4hq/LP5WLPvXVjjXiG9NpuSZRXvU1vCYwmv+rDCxhICJXB5IacWBi71E4j/reJkv
onJbAFLOhwjB9NEkeT0/TPIzZF8/+9BpBHF4sTlcQrK7OU6xlgM8Ehf/M99vYpwdUiDiwWon6toH
nlzuBtPeIvQ3K6ySh7KWxt/Y3nD24uj2sm9GM3rP2DjUPxCjvQJQIBJgP8j7JeJEzLCr9S47OFb6
W1EMw8Eznq8M6zSbt+iWi0Rnr3uTfWXna1mCDRGgdTBIrGnfcYQCfMKM0jTeqjvLtgrgVppOAd64
TFV9U3bfR7gEzATbEEahcedGNIfehkoqHb+FgzHJnt5Dli1Sb+3p1oOX/eBtnr9gQjovKG+rAf0Y
zIeCLN9iCcl435Td1NTSBqTC3hYopd6c4dkpoC4fBsQi05IxKvnlqmdpO8wSC18WAslpy2QLubBh
ningrqfjrV/B4Wj/g87NDjstg2bZVYHOyohfj1/HcFMbTRF2geRfqnIJHUHQ5nu2SW8YFYKY9ML6
CpTQpDKR4Ba471cUmFyI5aMndkjUaJh6bsA2YgCXIMbfGmUDKisOO9sRJcT4nDT8X1eb7DA5JKWG
E9V0z9kNZESsXY2Du2VZh6+fSYAxw/AVQl0gSL4ASdxjaPTfHnHnCr/jute6SRPucxREe7teqjQW
3LjmYPoyulgijXR7DND2RAlZC5GxYJ5EZHQLqgOzvRIawKjc7OkaSS8sZts1hEWbSWhwP/WvwuoH
vAvXDKr5jO0jZkc8pU1uuL6+hMvF9owkULuLVDG580ztwNFncGPHblZT/2hckcdQbt/1cZrt9QcC
oW+g7cfTTlSkgOGxC9dYGUp3X56Pv1FpuDmORoOx9y2Mnwpkup7hSl1OFskMCKJliVQmcVTBd9go
wro5XJ5ZIfOu24tq8JJa24Vk1ysRExCWqDMi6RXjo4feHdUznEZT3nWjFLeJEHEtRstfWDLu83Ss
ugbn2cbAi6w0JhYsHlTB2mdT4dfmpAGUJtje1FNbqaCgp5PCD6+wZlgyNGr5r39jAztZpoPG6E80
Bw07aU/Co4e3sw7yL4Cidj635966zue4SyQnIB4exVCOtr6RfYnkz8jSLPtbJmGFT1NFyogA1hx2
asOfxpd3j7bACP92pNE4LZS49rp4zdwNWbDJK1PIs5JO8Tf02JU9ewQ2zfXA8oBl9BA2ZjUq2mNT
PFHPReh97wgslJ8n5bfIBd8A2rOe3nUSGSwEjn9imEIx7tZv96wpAu/FPP4CvdE9338lxrg/+oXv
NKAIsJXGYreS7d8Bqo64AecEZ5VNU3KHheXH3b5vETclzLt4gpEO8CdOOyo1waXTXbhRanmKedkB
cMqVnZG3V9cD65pQrB6QwiyIKT93VbVJFe7AsVDU9bmgjbVUQP3oxc8AHnTDBZAM+rGUKdeCeP3O
a+ivDsQ6AtNDFd1h8EESVVaJ3E31EQ9DlL9n/dwskl6Pg1BSl+mPzztQhs1b28qTzWUfJSEI5QCp
g649pZ+lnbwpXej9amDorZRjLr+p8F50DJRPo0DouAS2gwUDKmeZPgqDNab5DXM5RyFFe4GKgBaZ
FTCxWu0lvMTZZrGkGHzIUbuIrsVylcAuoNDe8jNj6L7UqcH0gzvwo5azjoJ7r/vmYrpWNCeZXEof
vON6kYDT/SdO4lIME7ObDx6drhSk9e3sm5HKlQ7xSj9YR9Had7M3EVhIbEuDnA7li6pHqv2FbWju
guGpmHdm618nmFME3xwzr8k9w4iUPmlkYZkqWSLYV9g/LRSv0MfdcbxqZ0LAN2vgZLV6IDE8g+Wh
FoFOezmj2uUKEkSvJCdo+A0oH531e6Z/tWi8gIH8nfc84atpw7rRqGWkiuIVxM8yIJMgyN6QWTUC
wF4Dkx4wJXvgW6dR+8cYLU13y/mPQo8btmZr2FR26tJJC97waG+25trBEyeV4qF+u+zRXubE8TP9
QlxkeBnpAXhV5B39HnWNW1dfzjzNTkOhz2hfsqsQx7LG10TyRD++PbbS32wntcXTPLUf4iOaZyow
tw//BJge4oH60dE14Z2J0p5PvxFp7C322VpAv8HjpeYh5R5yR/bJFSVspSuXJCDHG6nIXqEi2GEc
2/8NVTcVYEvijwLcFP7H4Vx5IXSNPSXqq5EXcWhNiEfyF3o9GgXhUZSR8p8d1FXtYeJSNz1hAvgK
VWHZlokV9YtvqUWTYc6Ab1y0+iZDwkfm5rOVoQ1eMVUhgN53cdRzRPAfsZkvPbQmgZr86JSCta3k
mGqHtclhw5xoLXm11QUnlP7B4sfjTbFPk36nQTd9wotjCZKwMwFl/cy3sYt7tyjbXvDZdhBCMaQX
PpbJ3LvBs2uKde1uUZDtB+IaPboXQLMZhdjOo5+99vSVzYiCDOSYOJMPBhdqJMfCfgrwV4jxuUa3
OrBe9lcThcKJxeMF+5rjGjt+V7OkQq5JFHL7UdLZewvk15BmxZR6g1BCYNd+FQNjUiyjh6EYEGGQ
yexdG3GXDrI/LPyLjMdkuq2222TEteKbAcQ+up4e1tkSY8h12jHbs2POibCxLqS2hHgR/1W+P0Qr
AiUjVQYmJ1oGjI9YxJqgR3sdiLjxjyJvYikFlTMgh8bXe+Ro2B1onI8o6vRGYgUykPbTdlXRo+SB
d2QnRyBvHGJpFSomrk3SHZrCqP8wlqeQtEQ4ZpsL5vliUIAiloBseILItqOakMaJ3BsiduKDPBdB
JXndHWNKdq70s88MahIL7+3ZeMldlxkV3W6pAcxBSwMuQ7nOCNyE/R3JAh0MMSv/Uf2nKcmCl0Oj
AAsLGmh6pUdw+RXgJTcPXnSgKMIV/FxF2Be7NdneqzNCjMH8cCqddbQ3kf7onJtacOFosAcVBpS4
E0juXgYJHeglIVFqY2uvCtPdyAGJK+FISK9b4E7ZWJP2PLHSiq/pL6yxwKQfmSOc8eN6IF/TmR0J
fpVyfKOAXvHbEziR5j8xsfOwPBR1OiJ+fWQugkvLQ23K/ZX4VnPRTtpVxcHVdNcxKoXC4bTWHrcS
jD0vZwG4qZHCjcEwQRt0AQYNrCAV57bL0IPvYksDhYMAa3CgZHAFO4xiFaXxxXKRQDmA1bMm4fXy
gwPmGMRgRDseWjnWPOL6p5fev1rQ5kdhnuOGC/qsDRhbR+AbzFtXQR1q1tpuK2t67aYI8feOl+tv
2MI4seHlQO7j5kMy5GbdarqCcVOXK9jDxL4qQvBRahjpZWytJWoht+v6fE1tYXw7cuLOuOCkVzWy
FykdFiI3vBsxBoQmAP9qQGNE/TM/vVsjfc4qYdzRKm1YPlJ9yNkIdFEmj+AQaA62lZIkFsUfQ+/N
A7eLgvSV2zRxbEyJF5behjD+LBuWcidW8k4+eOToDHCDcqs5Rlb8BsuS0gAXiRzw7iy6obYnWxU1
0i7vFnWO4YjAiY3NoLOUQHMJsOliNV4uIUK7MdQNRGLrrpkQyMWrfv6fcJSF0WSGeCmks4InZeKW
ST+zeea1MOASh+Npghk5yZ6Jql3C9EZ4i5YMrHJNFCsnu+TpLF3yaUaJizS9KPm7u+Q5LM/YExUI
Ai4U98itu9dUrqYCCpx4u1fHiUjFEYgjIfmK9dglyKUbC3zLzY3mvRK0Thx880JhGMfDk8tT495l
8VjyiDHM8xhmOgq1vgUmYbysw4C2lDta7EJVBXlL9xiej5sFSNFN5g2F4O3edEViNWoJ2Y6Zsgpp
0eRZpK8kKxsZiPGdmtszuoR3c3RSp+AV/TTe7AE1ddilQ43qLiPOXV1gQErYCXc7nC7vh8Z5Z2oK
Z+1/iAdhApNjau50y4FlYYYKNGY1aC38f3NzYobfJ+5rKa88FPWx+uQBA11fC1XnJjwSKId48sOb
qXXNMTbVixJTc1P4B6lufqpwm3dTTb+BC8wt+QQaWq1pYFzf0c+ekh+gtB+9M4tYEE06IdHJ1v7w
TU1ciCfsULchWVldn06PEWuInVo77/bDGrGSBEB6YJPdtgaJpwBd7GxgybIgmFBIh5Wr8dJL+rjO
ljxoUii99bi9zT63/WOmPI0YpsdCACrsZ9JfU4C0vDwg5+FjEUFF25TYNBJbe755ViJ4rU0IXZbK
fLXB7DDes9A4KL6aVZfo8S+gkzZu0cM9IKE4r/QpFzrP44e/Jc60E/RdJGA/FE/DIbgQMSNoUFuC
BjL8OHoDUnqlzp5cjNeqHsFc1gu7QQvAKWLTPXp+ZQHmSfpr1gdfHzh2SYi0NpFIW9kqguoW1Gmi
d7llmpPBdvX3oaA2/JFVNnl9dzr22a3JlIbw8yKjLpsXjXfX4Vpc10RvMuGCgCjMVeXAGN6QsLC2
FmMwbUGDD5pYBuIZWO75gfbKXGWKJ3CHscI98+BMSZUiBSqcwgKBuHbZXJ+pvcb7sPg+HqjqMrKt
TkGxJT8WJkM4zbMhqXgQH2U83ohkgpFPdyT45DK5ghONsJibYM8LN2XcsszNdI4QyWMzdTFbBRHN
onfZWw4jONG1IjE3x5/VvLvLR3nhhZP1XZso9M95JF0UWRq6vT2xFWWp5+NRKT/p/3kofJXTp2jO
n+Jrj0nJYCktwOi569e8hx0vfgW/osMp7yDROqfHGa/fcfRX5wBJIgpmhDVOLyguuUS+pxBZPZmh
TitywuDviG2eXpyopZiBDEZ6R3pduqEY950qorIwjmsMVlkgDPKnrmtcH5bv9L8GzTWkMny4Hpy5
melJzG1ZMADe4faSQYVJfCMv7+i7oajkDG+vkbKX8npqxJ/Vyhf4BxPG66cbftfBHXVtme12Tk6i
XgWBfjEjGum+k80hlLgCWjJTgthBxmc2npM/lt0XhgYCAP+ScuDMW1OQ7ttiAlxHB0zSBGFyB2x/
SuTyXucmXhCpo1WsyY88c9RcUv1XCaJHAIPvXnJVl25Dyjfiqs/Nw+pY1sYQCeFc8uRB6rocGPhA
LeqECdpmgDgaQJLTuZXqL925slg3xUX36y/yCWMDWptkXxZqa/7Y+gG2fn9EzvWCDWvEm70tLtns
UNs/FAQkjNBEyEVAAG27o2EH3L34Ov+as1diSNbUvHqpi7BG1aoQ3AZRBvmetZUf+KAmP63URiKx
KQLZnmOYYoUD+27EWJg/u6lXArrW9QnKVVali6cyGaAxdV8uLDTpIyiJcbUtrtLMYrei2C4bhOqI
RvGZysTM+CzD+09QzQlOaefJ92177ON01/ZI3k1inL+ILX6dUKt+IfBcS7P/j6CR1cTvoaEGjJIb
VQakPPW7yL6O0vOxrxjWN69Onjl3xvfxREqT23ssxMExVi8S683nLhRSLxcrsBQMbUAxWK0jpHna
89WB4XvX1ObZC8aMBWnhZ09S1Wrvc5IsQVSV+My3pxyYgQtbxO9+BmzJ69TQWdrpgANHS7XCDRpq
n8d5SEFmjJnz24Jnj9AsgS1Cu8KVFFF3lfOk+LSwhMfbQpDwXU76qtfsHJ6TI7em1or9HJ4CQMj6
u10TxGrZNLVPwtpEpmPmSMoSTQ+dro18c90PKVufFMRn5OGCjFojKmIPptPN1rcF5Su+c9qe2yoP
uIpQCwtrE8pMqWwLapMMeXrCx8tOiZNoMPlHcRFqEV9+LaQ7PlywxReCjshF6p5CdmhT2WUyBz8Y
kzZIvYltI8vEkP1dIwg1mDAi4++2pp5gwGX96skYFZmuUlRTSqP6jSoy7PW1Rynyy6u78YLX1DBA
t1sO52iFfKP7on2jK4yW7sHqrhy9+S24xiaFC20oziDy204KE7PkmQM2qFFmLhLAHDPQaI7SsmYA
Tdd+g0/AV69ut+yrT4lVgTBZiAvi0rRmciq/H/96dzO1aS/JfqsEVY/mFqD+gCR74fKUt+S41Ov7
n8Sgkf0Cl/mkk0PokUg0ijzGQk1fvFbU/pRFDLuzmn7CQhyJivXDS+yA/MeIY9FjlBFM0VJ27qWo
ZugagqRFpL7xOp+lfKRN6Waq0LlkEwDaF8cyrYDuX1UR2r+xDiI4DvSVtF2VJCwgNxtVSj/gewys
O/gFDrHbJNXNY6a2RgtSNi/kq7Fug+55nKKfdrE1qFec/CisYWaPPFiY6nMQTYINteg9zPNhUII2
JTBOdazABSUJJoglx/DHYlYXKFjZW7eKhy+qD/ZG5+NiPvGx00iyLQyDyZaluOG636DOJgQeXWJf
2mQGtFGJSdZpT5jPyEOX9wiiT2Clenadm8abjP1M10zSRRGJkbFQF22exKqLFV9yuMdzpqXxfRKk
yujDeGblWc4tk6PbVWUNt4PZrPnv75sbZSibeFjSXXerb47gHVcBvvTyHHIhr3zDo/ujdGEvaIN+
9B1q6HAhVZ7DmCClxpCS0SpC4UgcFTmNx05TMzakdKAXMKHSLmzJaf8NR0btEcN8CKZAVdPCOs/L
DcCDwm6nlJUMV1IYqnoaYZBbn6ijigLCr54n9BOHunC3GaZmoeHnb5gJk1H0QrokrLCWr+w9P+2M
t4uX9bhRZthBtd46HP+zTeL5KQGk7s/1vuZILv2fAbF4Dehg5K/dNCKQDNYNM7qWanX2YsDIj0NK
XpUGRDC0FSpHVBG/cp+aYY6BJGy0oklOPe4g2wmDOsOmeOeW35ysG/KJWC8JsNR65t0kshW8r3w4
n+WGmsarDpYsD1cDSUWvO9HkbUL25JFuDCDdORPChatWrpxdIIcgCF6eT6hJfZFapzBbvf+4K4Ut
z9yn/++GdFpGN+PT2LdZIutVhSrrzyR6RF5R0XPrHyEV90Kc+2R/KE5e+xSHIyKuzOJfquGheKV7
ghD8QeY0sGzmMQqKi2I4hwQj4obmvpcOxG5NsMz+HSHWwkyFmkUyUtYPy6QCQfV1b+Anmt+OZBTS
6148tHsGkGrWDRDwjfoKM+VDxLI5UpmmCxPJYcgcpl6uaAZT1J02EbKNE5KDJz5gS0ciZT4fOK2K
KetXFbYSg9OyuTV3Vi1aDRja7XOx7QdlAfrxi82hJrwQKqq4S3CjIEJm+wXxHR+9k0YtYfb1W87k
MhcNvGK8THXfx7g91nmWnJFKpFx7R8MS54/YP8EWDww+xMjmVXQWRnDHhIwKY+wwMga+90vmyzEN
pIKck6K6jkqddrn1H+RzGcfFmyh8cwQ6iDv34nOiKPuwOicSFD8NRLsuIxjS/xjZ55l/XeB/XF/f
z6IKs6FM1nPa1YcpH/R8jSPBEMJeU8gEQ+j+u8W96qGyLQmRG/ShPVMmeM91Isn8rMGE/lbut6/7
o8t375oVMrsCfIxQriKBSR7Z0PscI1TP5GU6vPKRz3SwE6l7eH0NcYxZHi0QAApNAjN04O3RToJ6
aaQ9eRE2UqIzLTGYOnKwMnZ09MdjRZkGcuxuCVm6s5Q4tnjMfycI696C+M3gAHIuUDmLxvCzFn9h
xMCQiWOODxER9ixDAf+G5uFbc3gDgVXsLsuIwqJonnTZtfHSvxZRU0MhJCPaCSMWWg9fWhvxiY16
SYVxjAtSdcy5cvgBbQMwqyIoDwt/PnX16Au+ql8i3/09M30LBiWZrzZrGpwGcfg8xLmKWKtHK3K6
GKO15V2PmD5iWyEYEuU6FM8vng4LoGhGmgoERM8H3SH++qIzFpcC+K/Uky7kZBhcQDLCFY4ryyci
rmJiutqrn3WUcYT8bbm2OrbZSrV/sygWkFOYdXpQIvThOvLRDLFObHdDdZpfiOL97TjQ0fRkAYoi
Km9TY/J5VgG2b8LNSyU6k1mvck+K09fdVVKJXE5RqmJRAKJ5HuH7Jo3j9yfy8PdYAxSzHxe9L5JJ
IphG92vVrY/PDeSAnI6r8MwGOdMDshlmtmTYBoDwfbjOqvLCuBKZji5BqMP6Lmv4vCCTHyo5VUtv
hwGK8qQvB25oM9unMeWzukoXGBjp7L3jjlexoEyxHYysjTbU3pppNTMp3KRwkHR6go9U4uWtQRe4
PuPt7y0ExvvDBe2YqpPtROqU+eEukEiLXj9FaiDL7zIR+4YQH89YxfjE2WfdW12bDBoQQHEQYXq0
rfrjRG3+jUq+IOpnmSP4v6ECP962wH+vRf2Kwj0tOR/AQz6aKIOUhdgZwymilgAfyps/Uja9CPXT
OcQVQarTdo02NuXW9Z3GfmS6+S1jNIn32rav9w9VQoOQy+JmrNBfhnxdX3CarBupDMYPQwzhTFHY
iVqk8+XqE9dnFKAbIHlSbEf3bneQGBjnINXWw66fQYGfZZrUAayDtQ1h8np5irdVS7N6dqaK7jiU
3q9yV180SdEGR9se6dT/xvn2xGy9TTdtmPqkDgRDs4tUV2hxe/Nq9Qd6snjFwpxmKrxepSIRo6Fp
HBVqGsCuiCvpMggGSiivq2ULmIhMXAIDH3S1ZvJARBvtBOTAhkb/UgjT6yp1jZ6VTXI9K8pJH0ka
tPjAmwB1SKE5aUvgBOh8eSRnxUD0ZJsRTBihRXFTRiL+Vr7HQpUJX6pHG2oscHyYhEhhCk/ACj6R
IBeIU/3Za6iXugN1OHILQm4gUEmyl0Ew/RrdMwvKx5nOvpqEJ01flAVRTxiNSml8DGRYMc/y3Ejn
5lW3rQ4hMVSIWVY5UrKXF/VsiiBQlKSLa4KMKiMawfta3++aFR/3L7ixQjEnSuJxzpDcEi+Stspv
FTQC2OXvs/+eHdmhnzZ7EBaiOhdxQOeuRyrRkX+gm+3Jod0psW2bzeZbaM+Jx24j9Lz7BJQhGf/7
XPs9Wa+L3JLtky/rn/H6PsZwO40jahlIH0UATUN819PJ4kGj57rEIlSQmichAuSVqhcTAHFeZ5m5
SXcS2yV68C/rCJSsB0Jd8JyjMicf/YvG+r7xuEX2xR4nmuahBReIBsLcSxPFlKSBi1ZOOyfOChSr
iojsuCYfKSYnLynqq+716vrnQDpPs/YsXdyo59van1A1GkqN3pdoZlnDM695rA9+dIxFybQm35KB
UayhrgrwT8SeDYdT9hNcOildzrxrOVXCBieSIRtgsKPpjeDghYIBjikQU2+mCGK6A+8oXeFvxh0y
Rf6qLAYWi7tzZflFABWIG8MZjQUHDUgV8LWDphh+on10gyPy3UF3H4Hqr15CQ2x3OVDEFNDG0U5Y
y+o9LYfRpmOuzxTvZuVlofLcnse3G2ImujHqGMN452RoYcP1mu7dIQxJhAXtHzFIo4hp5IVMH0DK
outYjgMtFy3KZ0lyNJUjz3mLylV/nTywMleqH24P5dAC/AKtRy5oBwDB7lSVhf2eUEmf/2oRV0CK
DyGG62hqr8jN4VNKsy0WmCv3He3ET+IelvZFh7NluZCk+fOK7jzRlKYXD/YiOvQwSjLdhjRLg24o
ZQklsj+KYtfPFHbOL3aVaVaUbnw7MTx454HR1Ep651vAAmJCZD4ehZ8yr2u3UxCI2K6mXuTtSHvC
P6AFnfEDplQ2jpE5+fTE2EEWnV/cIaGPPo5TJx6VHz66covMZo9Qs2bJeW1TE0zmwRXiqTeX7Eos
boPBk3qjzxktVapMY7TODkmowXKEwBPt7fAzSI92XoizNXuuQ9F3AhJPkwxjZ8oQlv+BPD953A6+
luoboGXZ4T4oX5NIh1e+zsSxJJjr0lohFM9373uuwHLaLE8vX8ea/8IMmYeG+CCRovEhvGFbQSYK
qCdVcrFFAkBdCb20ceCBVzjXVrXiVEOIV6wPRzk6UN13Fvl0Zsr+usOXQmhvgGEDLItXbREHktD6
k/H7F9lhUZIpoO+YUCA3+/VJgfRTMawOmEhAQQNkZaKaYT3Qvz9LUaFfpKfUfS+oB4A7RXd82/Mt
Z1T+0gIDGmSmL/fasrWi2sM91TWoUmfCM2o3H6HL+DthmUt/N2P6fCo1l0J7C6v9hgmIGgsnKz/e
Wudrp8xzQNqf7CshJSS7tyRVIoVYHplb3TtRjjJ1RCF47qlrmyt6k6uc9kpPtCAOy3flK2/iw0A+
RjKSnOodHvEO11OPAaUYSEicyhUXxHcF2+JFpSMcoA5wxChdjSKvpMUPCUeKmCSz66fwl6cJiX9s
zzWmz625FEXjiaTEHD+iezoHvVVpX6gLA2praE2hHh0MreNwRt0enmbyNS7l2MP+fFKXAhqHjDw4
kc/JgMLyROkZOakmj8s7vlfE7pzgtsLrCVpGmZjWMT/cR+ByNwhkX0yKVfRvWM8kTbPr5Er5pe4u
oaPoVH/TxiZNr+hdOPbcBH4UosObVUvboBLtylZgibCMUcgYKNeCRFYnMk/QbUKOOG5dbda6T5NK
Yi3gbGMMm1ktj8rkjtVC5T1IU7umIDrfVm1dbyhDtCFkpIxhEe6v77aP4HI508tZbNqHbv4wY5Eq
2Plbm3zgStCniBVQxxODNJkLWycJ/vMxu9vfhtTu/Co2OAT7hlZLLCpcqhFJCDXPCyl/uKVAI5EA
oR8JdhjwFgRSsIDpG7fgSsPcOTw4DAKzbZ0X2M3MRbsdxg2rCTN/2jOAmBmAMiasc8eqrutodphO
oT+xRIGzwaU0RTHEzqAIbCouitZYMlbyUKUO0DAFCewUwuUQL92KCJoBLML//+rJQNTryFBmPtog
KfNiqnxfU4VdRrtkSIKAYgUiAfTCSEC7lhkPqShkbiZmnUnTmUIG/z2p3D0nPLTqn7FB+P7Gjpq+
1O3IGtn+RFkmVs3bxtd8Q96t/pc/T+zsh6sh8OnyrDhQ0sgtDu9L2gaV6fLYizIWjYLwhme6hqPU
JjxnnbOYQU+rBvKiJHS0FTyfIulDkiPAlpsc8XAvsRVbOucdxtOnFhKW3lrp2K3sgdNy8vVhyjDE
Yhwtj7muREa/u6TsvJ05ZdKQROzvQSoyqQW8usvosAYPS9nEGJ9KV9jIWt5CtOnTd+7p08DV+CJ7
9EuCDxxvxFYIFQ88Uks4ZLf+l+MOa/6D4YR7VnLoMviINVqmoaTYjlfFY9WyvrUKKwsPkEYm87BE
1b9Z78vqsCSVtmnEYv84Edw483jyDD3fe37v2DItQffaWvv2A0wxx2CQEr4xGMQia788PjOwTZtC
kk9M763z2k32bHLK1Na5rZ+0aeMWAYvaDkETN1NS4ly/Sf1dkxZmgIBEk7JpNbgaOhUsIjutL34H
7NE2B/2yhaz5pKLfsZGIA1dtRq5VCqp8LT8cE4Ygvng2Pmulz/7O+TWslw7vPJUMn5zwDAl71kXl
So/nVgoF4nmx/gzq5lgW6ltkM5pkVSeJEpJYvME6WBa0CMGm9ha7Jum+qKuAzRMah/VIj9unkLJW
y+ZSIhfoSUGiXvNKM3fWQQYDNOr9RHZMDtA221jJP1NMyQ9eex/DXJibo1ZqLNyW995QhFNMXoW7
R+INwZwLLd77QKBdSypMzDXK1gwrC0zTkH+LwbV/YLbYG/FB6XyM0iC6MYz0dk+vFjwhoZBbQKtY
xueExgqZgIWW2VSB19fFbHaAScN79mpYFNMKMEESuvsmhpmgwMqXP/uUI1V5JxU35PLCC+Ezuw9C
crWvSbUg/KBdu/mjZQ6AeTH4aknIwtKD4fFu42OV4aJBbN/gNNNXSGkQN8nw23XeCzlxCIyLXgr1
fn+F3nZqK7eEENr7MwQ27q1PYUIf2R9u0ZosdxW00d4eb5RuDVGVlChu/vKftHA4XX2FpKw9ATFa
8f03RzgghEjlFc6furOtjlJHhlnxRkrvomXXwsIEJKmGuGSN+r8Ji+yUEN3UZUD5iSLMvyn2vYI6
dmgSZ7mlQcpQ2/N0yp435TYkFNVOZAZ3PPZyAVc9QFwr1fp36sPsavpC9t6StavXuNTxkhDOn+Eo
vq8OxxttKECIJ2n+AakLxsFY1BZh+Xg32zHPljFaBtrmQ+rTofkujUUrEl7kX7XmzzY08m5T8PN4
/a+O8X7oIotK8xeIR5xc9P3UCOc9H4dwuLGCrNVDQMdnqwMvu86uHhZ7Q7TClvgH56CfYmhSywRm
9aQCl6DVC+Ft7eOLEqZUXNhR4E5dUkzfOnRl4K3ExYddeXI2Ty6g03a/swSkHOrAndCn1mIcCNfq
OsHWbF0G2pkxH7EiT6J1ZQZwj+NS70edQQxRlBxpenbUrAQTPKZuvNPBrNpRkvmloKWguvRz/a7P
WxMJhU0OzdXVdpkso10GU9tVVaMXzrgA8o/uaONXA650lpLJEaATVnZC1UdSWvUKpOaLyQshdw+s
9UUHyqvITiT14qUtBxL8kbvhfnd5UxJrCO/z2sLWEo07zGORldA55/9C3lIV/NpAHl9+eFiM56Bq
zS7rU6VI506V11qatEZvZWvupUcUxNsx+TwRlH4Y37+8/mRMGYJ0ane2XiKG3wDTtCu5/uFVRt0I
Umzi9IpWotNGOXUtm/Y0mPpwv3VnZX10tplhenVRsKZw0iRSVXqkBGLp5CPxA685Y4qvyVDrrlLs
6TZVY73Y6NUooS41rUMd68a5Cb+kT1NbQyFKMlvxhFX14k9WT8oNETbdOQUZ1FezorJbIPMlIT9/
6tdFIS0UHPa+ArpPBIAUDjNpuSeJoUqsfniXdYPUwDwHIbHrx2v8cKN11McqBP+6mccaSDH9fFxS
BoMJGm+vV9wSSolD+opHYBGA1eOiAdPeCb8fXl74BF3A9/OQwWIKd7DNltDUf5iowEEtGpmmicyN
aPfkQUXYDX0MpOzfa0/vRQGJRISojTI5vqE/u++Z1RNY2Gl/I0+kKQJiPu/3xGv9jDQyVKQ3vLNb
5YxjL3CJkJ38trlzYGcWI8TdGe3Hm9mFnkEpBk41bJZpFet6eMHVvJukv2xpVlsQvW4a4KvT2Luu
eNvNjcRGNftzDUh5Dxp4S3KDN5R9g7isvyMKcNZAca6MZAeQTmj+qo/gmaCSY+1c0nyn98T5V/z7
9UzdYUXauUXoeuec9ndGAbyp6SIPGonLqPotk1yDKk7yMCGqlSzB16iXaC2CoUSiuMUk6Ct2TkHa
ItlrofmRPQfQW8zE4vQuiSTdr1yZ6xm9Mrubk7hC+R8SEiIdSZPJoamdQ115RImGomF8DBmTFEN8
k5hnnMniXVcgpFMQz+6KLt0J2ovNwMCW3OIohDyOpzedZ6EJFJX66qDB/NHLAZMNNGj5Kyp6t+BR
MkD0OBVW4/iFfYMWxwyxXNX++iwHXvbxULlJNC2O0h7WsGAQIwLHaG43pG4jR11bkuVZMIbQmBt4
uh3I5HKQqGKrOGYLrS+3OVIblIgMfgMPXfJsE0esh/VFVt5jtgxEzA7eUBmFv7+I/BQdU6DCRY9o
SN9BNiyciqPc4JKyb8BazNmS9WxAIyucKTpcfaUf5R5Xd62zyMaNt1SMKHP4cWjCOuwZQqWaJHKf
MSjlb58vgpLy5uuUpGPXGSkZXiaAlAKjvHH0KY2BvGMg8ZW1UqEE0rKRvWIbxhdPBzAP1bBeSfTW
C1B6YkkHLMRYFrRBWE9QM27pWzqWd1fZp4WVilDDCP7clk+I2ffL4Fq5OdDnv6Nomo+Xb3M9bWx9
JblPf2lRH2OPFrtzadD92XPJqgk62s3dLwFO8Ym/T+XhF1Sl0kA/pzz7oLzYa23n46l3OlQtteKA
UwAq1n3c/XrYyxAuDf6WgkIXnfv3BwcwBajz7C9NeMtxmFEAeWQlR+e7ebr0Nt7SccxvAWqRPab3
GRFgQVCiygTHcfYn9GvDV74RhjCqf0pNWnDcK0HXpaz+aj+U5SkyrUqEc7uDZqiip1Z3ziE2XR65
W7qfwYOyAmRKworWo935HOA9rB3HeO/UMlK0xiOY49debevHRW3aJNwnG+CRqhr+IgWnpJvVDAlw
mBNTyo3MlAVXU7WDEcC/0q1YZWTMbhcyYXgWd7qGUMMsER5pJeylVbn09Q1GIjlWaDkEf6ep6qqG
co4H0GLHv+DnIEdU6tZuyUJq482e+kuj7c5RW8G6GSF/q/FU2Y8UDdk3cAj6Zo7OX9FJ+UvOmwes
s1Fx/RNUnsTikbSreX+Wom3t+6MtVKNZ79Pf9Q9ejh8i3qRPbpQWbjsCojK934K9lDLZjCdvXui2
Txg3CJkP+f6hAL+iLIf3tc/Jf444C5gWbie6xhgyCP5Ph7KmH+j1m53Y+shKei91G95n0zCfiueW
z7FDX61fLidQM4zgbvmH95w6LuHvaIIly4tbfOjYNhnRKJ6Y1R9V0esDh+SQJPNw3g6W9B4RiNlg
gqt2Ij65VbyOlIvk8/IOVrzBA2Udf25HHGG1B57bBWYlpXDS8DKjA434eDIQ4Zoex6Apur44Mvps
BAH4o0xfhLBFBikyZwukgtmR3Xfg5eHFoBtmtPoIadNtrQeXeP3yweFjpzzukke4uP1K0nxGAhNn
4UOrxsDLZKLocjE19Axep1fJQK0/635c5Fu4805di9kiaDQgXbeEKjYXfyON4V653k6odq+4l0kq
TSeq0yE1iKSNSXgWHjGEGICCPs/OShXsnLlaMcI+gqT0p+oyhJj/Z3C79L2VHyrZDaepjL911fGu
H8rdsqoZTJ3pIOLGdyGiPxBcPSIrZvX9TDuOzFMbBIts7AiIsAU2eG6pkcBYWWcmFrllEByvGbVC
zjfOuD/oZ14WSNVO5EHjUuB7IdrA7mZ9zq7VionYyikyST4kpkf6pQ3lfTBgzLq5ArURt9aDX4mg
LrNlCSxhjyeX0qPa2s3fwvoTWkCpihgpoBsphGhNr5k8mqmz2Xc2wHEMuQG5jOeQKLXrSNv+amw0
KGIDD+CuZM93p+2KMDdSyHfd1ruHU00fq2iYNzNk8Dusxg9DwL+cRzTMooSd5BtC9i6gBvBYFdzD
xoLGiOSccRqNQD7C8AFSzvMIESEYs5npNrKDQGq5Qg4esX01pkD8dnmTEwtMDn1kMdzmz07Tlp4e
BFW6xIrEfbSrFudQN+lJQZlRF/3w99PdixAQQssFnjUKXWsEloIMwYgXupufiZEvL1KgNQJHCeCn
WP4X/Ft76EpYxNdSoz6Kxj6zGzCqP8q6QSHL0AUBCP+YKndD1r7T2PKN/Sj8pf8xgvn3IReJQMhM
dI5Xak2fQPR8VblYGj/hOIePGw7QCfHMvTC476qos69NLVFT3SPddo2BNFQt7sdrHHnRYcXIHOO0
tcnC3q0l+7C2VUn490rIB17NRS8bjPlU1/wg+A5411q2A0IunTCmZvhVnYMY/X+KwqWWjtTwVihD
7LEqW5RZ9ygMVbx4ralNgMQ3/Y+V3UMjVZ57waqmFU3YEPbAOu1GNDJJyteEg37VjcUct0LJ/2vM
Le4a0FlRvuuzcvyFRg0zF6ezR117wTmOCQot6RvIp8uTAF1p/3r1OVzUQyHe418qDoWbDrPHpj+6
mbJW3UTvxdu7WV7MZvrTp6XTXBdi0Si+fMHX5T/e93tOqEny9Bzbd5fygo8aNloE9K2HWoxtMKto
eGYHPao7cp35OkphvsEFgTI+UbvpZbH0DwJvpt9W2kWrepFyZyjdOC3MwM2Q5aN7cKOhvKPhd2W1
KXVJqjgO0PZrCOwsuQW0GZG6kKWSKMysGht22xvHBaVBD/hul6nv33zaS9vmtZtz2Pgqugr+evh2
USzcIDrgpVOYT/v338IeLpbe2fEJ4EKVFu4GKfa/o00AfCYoCEv5y09XydUQF5N23SlBsZf5g+Vv
L2JP21LWPHDAm7evMIuYoSGo6NT1IB51c9Ezc0Ifdfaqmd7gC6Rc+SK+bj4NDD4pcDLfIFI1VcYZ
RuyfK72XMUb+hhZH9Dftim1p5x6DMzhqzjeRzVRxo5fsNG9tdOoXsxk4RcjWl9p/Iqe1q7Q8Mamx
Wo5pFRCkGMo4erFYwQc6eulvfwV3D23NJcbuRmtguPo4yDIN74lYiLmoMb3pLMNWqxZqgv45Nb3E
RgRfLsOdXOfFW8EbF6U/RfRNlam2bx7kUxKm8pQ04Z/nWEjdSFQ7dO9cBLYk2oXCHJfiMEIj3dcq
rLECfI783S/R1Gp7tisPfkooahglNP6h4cDYdc3iZJ5Xrj5ePdjfcrCCj8OKzpAvdlSdrBMXQ5yR
IbFckJw+zzkgmC3PboCaGD2Ht6waA+ejIYVBQK2YR74S8Ey+xPk8cNR0YMd8ApUk8RUpE1zoet6E
3sv8BqAdLCIbsZt0ChIh2LfbPn+DT2DlGja5ULCOzynYjOETevgcG+4/n3+ftlKhs6feY5UobyW1
Zd7M1NBK1sNbi+xXDv8CMJt6yG3RIOraHJU3JeRt9zKaZP2rZm7FCU/c4RZxOsG0QgjlNCZ6u5Pn
iYX3Z9v09Us1YMeXbd0j6eK3c4xpTdFys0wezf1hX4xbNgFYsYtTkZfzj4rvsHwnTmckgMLXDkZL
aM0osQ719AV0rixFl5UmEK4rSDsgSMTTCx2YF5D+zj3q/C87eEKjJBILAJKChmU/rH1ctVbFigNV
1iCBt5QHdTVscdv14SYOIPessZA/bjvavrpUZiRgNgqyBymcSpFxiSYdbUVmRzcrA01Lr1JphPFv
MBxN5cz7kbQDG703rTuH3jQ1gB2oKTTnssc9W677YatqQckZI+SKNTclUyysCa4T36wlqQ08ineH
tU+8gE5V2SHFLFyorNLsUyBbnTKQjSQwCJBAfMB2CdZjC5vuoeTfleQ8nU6t91BIGX50mfrm+WVO
SvwqcwdY4KM2EnF07la+IWMqHEutCOqmOI90KXd6P0k6HoZ1SsmWXY/zRh33K0xPqoGX4f/rPDJD
dlV7vkXSr1gHJZ4LbHiEgwUOo6Hw/LKPqy7gfnopBxL8qorYjRsnh4PUpueAwJlsBoh/IQBejHae
NsORhK8sx2GDWXtRHY8qQOscOTDXREYRcHJkLRUZeXfgY/fGsEVyPa1TKAH5rw1v4LdSRHPKp+I9
APL65JPqwszChkXk1z+HH7kprEdnpMI8AOjGkDW+47e/B+W13ozhzXx332vmp0Z8KO3chHbIYsSz
p/IhPay0RWW472kC1st/vOEY3HxLdJtUAueetH2FFwxLVDLRfEVkkB90jrpoA19af53GIjETvni6
gG/F5yuNx8174MzMyqcVmUk9jgqwrm3i+RKQ4xHzjEgl/fzsUZS27mKVOm1R685hlBI3rH5XrP1C
Is+aO6iEANfUmyJb9FS0VWNYhVtWPtLwt2YhU3B4gYlb7ZxPkvE6xbb9H150I/7GLmcvjg70TJkN
et0wNh3J/Wo5RBXzNhbDzabTpmiGhJQoKFGRAEQLGrWtH6QZAGUD2vl54EvX//LNTxyRFZCIm08p
OaDrwlkhdN0a6vJmGd2GSCey67eugAfyGjpU+lxi4sgk5g2Sr9KJJ45wdxHuq3N7/V6QnnReCiMM
FaJIEeA3t0h+z8aSpSLtVtJOogMj0BJRjgk2pfjr74IgG1GMc/eq4Rcovb3Z74W/M9xCe5apP/ae
uj0v6a64oPMRQrxlQhNafN0Sk9U+jXQwDVzxr9mG4yK+nJjrYHCAMkMa3L+jXEr6kz8TE3IoDapT
ERCwoUNTUs1VdLmX1yT7XzT4xD/r20FsBOhtbz73AAOewJMbosWTW62pIChTRdpYJ8QWUQAO3rYf
hPZ/DEIYdP1kV+cR+Fxq8C9I50BdMXtoNvNnOh+XWB/Wh6vZz1OnafG2ZOgFzNsuz7Gib25B3dAK
dNWYiI86V1yHBR4oaDJwCoJw0btytaToZXWBDb5iSwvEM2KjOHjJENF6OUh2Jr847FhPhDPjJg4T
BOKpMVP/v+TqNjVxzRBtqUVJClYn/O7zWvoRipZGlFgtV6fvqABcwNvtdE5jt6RKKnmnml1DvFdh
dddhNwCJK20NWXHv7CG2pPruZmmuGsOnB1fqE2YMFPII0B7+56yK6UrmiFLVyoc4QSVjWOUXaLMh
sOPJy5NoilLElljScRYR4T+pIQCOfmag1kjXdxj1cLKrHQZ8ZDDav8LfylxrICmGGAru+oII2ZmO
L8mRF4YZFArcFvg8VbmK1LtwHBOeCnzkWAQIVhIgFUyLmEwRqt+cpfNEg7TkI3Es3Ty1pUd16oGi
6RJwN16GwwwCGra7q0DQLx1hR+dReCTCGy2tok5JAgzxz6vL1c5OoVOR/oYZ0s2VBcR0V7+TwBB9
0ReUSYKS+eJOVXfYt0hIx2AKREZg9D+4pGyaMqYkaa0C/JkT07DILBXZ7BnldJHX9qZ3uMDk+ZpJ
HXt9Ie3udA188grc9vbzAM7l+g/K8NgAEkXL9XA7g9ANzuUFf/8X3Ap46YGCivRS24jfwocDZer9
OfYIWf2Dopseu+ZYToBQ+fU6TSwLMfJrJFeAPzKHED4kHSi3brevQVanYX7VX1u99q9/Nf1g8rrF
/9krz4bKs9cNtj522+POQ4TkrslGZcargU9D9Tnk3YDBOeqijv33y1XBUZXFtUNfpLDhU1bh0pSu
sQ89ZmQza0uwH8Yb4DCKlD3XRkpdBL25HuNCEanjsbPy+DYmybZ4GFknAkMbsx93mmCqgm4O3Abo
EZ3M5m74Y+dBrDBvh5tTYOlObrEVUhxvpjKjv+tkLYc7e+HFEY9pMvZU2xSc+Ya7i8e6iS9wqTdu
Ijzj9Nhqm5D1pBfkVROSK46yqJ5f2XkYmGbflVhEs6AEgCVreF896iKdmiiUUWIbCqCQNQ5ZDmg4
hstJR1iNXkBFYQ0Le6eUm20ZXZrj3R4zhgESvHRT22hDu9P33nfRijN/8dWYyUIRSPDqG9jAIsdH
MP29pvfxGguCQaazLf2sEhayUaviEgk6Ha2SlLNFnLT+cF8jo0mHHialbdjf2javj26AeM9xsyWX
JF8/Tm/OhO9O7u35bnAZ4FZb9bVWokmZ9w1SSIufRCbqRQB7c9JDE0QsXuczYxcz2/YcXTYuuAXt
IAzaqIhqol4RicTGTMM+hcFte86kX1STug5mO7ZMTuew7U1TLx779eoH7YH1pJ6EKoRW0Wdyisej
Lluzzqo4c6kw3reDXu5DdsDM8Ku0wGFfHWDYacEkERiCFm0jHA4Dd5rzWAz27TvqBuJxuWUVZPoj
SIYFRIdfWEoqs3lgKC78JWkXPPPhKLPTNSJlA0VC5VlgYvggBZukUPJd2UDZY+/utkmpRNZW02pK
mnHT2BSPqtyQPUNLttEN2T8Qg6WgDhWKBuLTfgFMuUFKnnikdNtWys2SdkyVWsOsttplsxjuLBWJ
OWr/vdobbaYNF6L7ltU4f1k1yBzpf3JcUbkSr2T2ae3Zw2fhUSSDJfE71eab/aV1cbGITCIzlAdf
d+zLXWEVfQaI2M2U+AbV6aqyk4JFiZN5qIiIyqqLNty8GwLRZ9apRPxNI20YrmNYAl7TArj3/R4u
bOGBHFCrtpGMZYQtQiUyeux2V7yhZ6XH/S3EPJtVXHOTa0ZdRFO8PXZoyHvuVlj2+cftw83oNkdc
wDkueHV5PqTjuA8nEyGf3iJ/duy/rxFJ0l3kkcX7uHXs1bNN2lVa32RQewuai3h2THVtdpE0dKYe
Ronp+WQSnmeuC8c8SV4u2q4Sx9i/FRQbRRWQBI1MGsILhiOyPHXWR1A4IWk67+44sd5LvOUtVK/k
PHJdpslMR3mAwWEVzMV+UgPztE0vX2Iiaz8Vufs6zfe499gLD86vunI2cliLyZ1FLd0IIn0xidnI
2dOpKZMQJn0N6DH0HlO2koWIurC2cGi0rvuY12oNTmUh/uHgDjchYsZugpnHv0qdpAfm2RlLIEdP
/IHiRlwiZUdEY2qOd8vCljWlSpIwb6i1pl0ttd/L4jWQP+LV0Jc9i0Bl1YsUoYIahg4/hd4ubFVA
43HcyQpv+hCzxn0ZAEGvSw5qXKL1BfOegzx/DGWn9zVXWhf1aVzDjKWWtHzgUlmB19D7az2dsAEQ
DCoqqSs7F1ebAI/OwIqRmZyY86Ymph759DAizZcWhniWeSPiXkArVkUcZNAbypNbEzZc/NUQVIXE
m4zAdJV11hQoemHcj52u9+zkT8nKMLwDZqvQHTi1fxZSR3j4+c6Zvvgraab2gg/V/EgrZP6X+cDb
gvv8JbIzwu06ZmZuHQUI28jb/1w/x7yZvFmisjIbMtMJvRsE82mycCpK8QNB1l+RRup8DeL6x+QZ
QLWYwQQaCY/7eAdDvXraWpXJVrqyIJO0NMKhImyA5vsGUB9ACRQ8CV1EQhEl4RbjFC+hW51zmebh
MSVe2+F0GLuaInvKun+PFccFHkxEJ/+ClLKPbG/uQXJFhrPj0A22TfT4HGuP16GeN+TcbU1S6BsE
lT3v/NZg6z2xzcNQ/lNTUS/kMyrxywrlmdR/VneyWbv5gQ7/y9EBcDcb7hT6HnERLtEWET1PSOny
L/RyChuqTMRNeRSUX+KV7iQxdVBp9+o2wgZ3dWblPlfnMaWff87T/0pOtdXyQPBr36e0g4cANAET
y4MN//cPPsynqHl+3Uif4xO2urX+E1TQvOiWoT45Z9R040xf5zFtJNqPevWz1hnK5GroNRk3+a/n
6pqGV1KzBOOpEgEjHVJmNu8IzaPalHifYiX14dndkRD+GDnvgemV9DlSpM0l9zlui1AvIKffLeNp
xpAzw66fiOUchmdLNpcx+LA6D+GquHAvR8g2tTkmxbDC4NTtaU2we9joc63A+ETj71BuujcfRCwn
ZVHOcfXeyWhIfeKQtFtkf+m39TNWISxpYRYZEed4jRISXGW7JUN7x1o/o/ILiJsYlmL/Bsc/ja8E
hToaI+8EqAbcCE8G4/wXCB/mVlbkVPC4ehqHIY8sL8SR4NyzCKcMH8f3FNh2Umyr4aMBt6Y/JmtV
VVTKRluwTQCLu/uqlw473SA9UTKboROrvtEm8+wv3VbB3Y2Knn460gGI3POQt68OhsJ0F1xeTvoz
v0r8SJyHQKSV9ivfeDvqr9JkpZpV9Adnv9e0C8hoNN9U1iQnlAbTFExJleEf5DP+IWT4JwowdOyf
xedTbH3FCPhNxgJbWshTb4hDgykXKG/ctbjpjLDhQf/thpj3iqAnqDQqwx0HWlSkCF5aWlimGq/6
UJEp7amHuummurJL5rcupWgBN8EEBBl1laM2S78su4sAXTtZ9d+GhE0zVab1kKlUvm9tOauP282q
NJSCQWrKwCWtxdbQGZvfwT7/1y2qkybKOoAHp7sj8JYldS/wK7xeZR8mgmXPgYpL01PMa86J88pg
DCi8QVqWxYjfJR2VLl/gE8v0lAtZpDQDlLhyCeBoK+2fKDfPLNGeMmQ05XMO4CP9YndkTg85Gnzv
cBl2yrngffYMgLNHLuPSlEvPy9Kdr9eSRr1ZZFvbmslbsvV5OZBEPK4CLUmZKIV4JoBpABXlh3b/
GKxihPCRSiKV3n/jjs0n2ofHehP3M18e4/YoiDTWble6gAUJRhx/EzkwUZcG0TuohGGYAxAb7W9S
PeSUA/wPIz/6hysvAsBxI3H+FKsDqQHj3UUXD0Q+DM1x8nlaklBBccDNikCLogrE9ZVyH+qt/8xy
O5+gOM7NSTwsKFouDPT/ciKiiRoBruYnH0I4cexYOjmJS7MqT3/AlVOhkg31v1gVdjD9QCYpSkoo
hShgJwb8XqdrNx2MpvLqB2hTrgEhvGqEhfDpqP+fm2x8S3cCgiYRTI0jGEQpjJaK2VukIHjA6bKK
M8wd2jZSkfE3WNcKTghdP7oxYPZN4AhHjetGFKtN5Xs9djg75Nq0W3HEFvOfro/3o3Xne5J1RQru
JwhhdCgrDsHK/C4BoOljMnmRS2YQsyj3DHT7XW4LbwHZSkg1ILyykNPZogiJVrVdLFmRtHJQXFlu
VkLRGRER/tSL/dgiQfbKS2v252iO70xuxAUefYVBnGAsyGw1frjM4Ii7AKUz8UWmIlpV1BEIeI6I
Mu+KvXZqXOkSSUmSwvNUEPZ6wt00kg/HiIy/DLcFfSLR7S2tmgrqU9jaV6KXwhJNJj/MP0iTYrZ/
6nhh0uw4D5LA9WSdnII1Wf4KRRUjiTFVthJ65/CVM2OMWi5c69NMFuP0uE2opm13qGnIH3QWobLo
76wK6JVkQdTLKZDNjsGqjCgqDGK1spu0wwkQO5x3lhfaG0Qg3ph96E27q9CNpy3tGUDiR4AVF0DP
8VTnRFJuGmhl7zYAdEBCThvAazQDJ8QulhkIpIZmjqA78T4S1hVZgCZCUwNbY7V/e8REn3aaukba
I16Kbnm1EBSQBbmZsUDtRDVAPs03eDBgAMzRAeTxqjkdNNFBMtT4zDIa/imUPhLR6yssfYH2B046
GXbdjo4jbk7M6mXQIwpIAaLTBxdJHVazW+v8tSckQCew3n5XhD1QHox/2ux/jrEVCM91LEiby88P
7/2VxfFIlstI/9Nz4ddJ3r9JPdObOYENdccnufDJhYPRMrzHZIKgjrATLCN52AsVT0WO5OupSWOO
3wzVjumqPHXTUY1dms9MEJEzcxNUuYrxG6A1gl6Rb+Gyxtnf4CVAWUGmZwQlUJByf/G9JNWDtf44
cwatFQv8l5uimYUCpqHcqO/NIgDSVxtPjVNcy9KSuPm8xZYYNGsfwGUQfqu7bAeRqM9DjdYT5VjO
Mo/nJsYxZ4UDd/TXlWd06kFX7UjttiLtLiZPuf3XlZsep3h5/wr3IQshxMUUPVCmA7FsewDjnzl7
3LVAggj/RDUnzGgmRvdbLISgSHxKeRDUWxuLbr6V+oz9SEGssmfOHJT5H2IoQuTs8kq9rBc4jpo8
r6FdRJwGfV3v2NKOB3Gw0DfxTdeZpsM8C55RjQD0sRyERScBzXNJKlc4waocLndMJN+7K5SNZ8Tl
HnG3UlMfO7cD9/bDZytCwDBcxZsMZlY1dgHem+2SVKRGruioPwk066yqqMZlaNqswS2BBoJGGk1j
+NizLNtNA2Pezq3eOXtUmppIscjFTD/g7oGQPc7VUJ6bLZoopmKSVTqtP92SLyu3kEf/VH6m/TYu
h1EbidRExqyBislRzEmMo+tNiEYawuWnBBscEgTo0MtOtHWd3PauYuQjx14XsxQC82Wfeu2k5vO2
Mj7sBroCMNhgEOsEIZy4/E3nJA+mBbHESwKJwh0x6Nx3vJMr+olzVYZ87EwExYkaRddQ2VqPPxNE
us21jUUItUIbz1CDAjSca9Qyl9ioIP3gmWH0PuvPR5G/Ny1eA2dnujj0cDgcMRnmZ7eAu/WeAF34
QsYdvJI2iHeA/jOVZTD1srnX0utVdd/bQE31v43QQ/9e/xlxJyyfVgGcSOkxIYUeXXK1UkE//EHt
uqLjwEPjAjP6sclQsGYwRf9Agrsv+a/RHH1OvzJvomBE4W0WduTosKaCjRu99Lzd7dMvMShlB2W9
lpy6TEtmKTiExNbxTWe53zt0LViWgY/Vvnnx/acQ1tqvM99LgaWaXQPTv6OblcT81RGaIygHrH+Q
d23ewr4o7FL/jEyCTJ4/dpDkB0oO8bHH6EItWyuV5u7b5Sh/wDOk+6+uJjqxk4bAfl1TUFzQjzCB
MnEFw8wCYBC/lfTQ9A6qi04prDkTFcVSxQVrmCdSKMjQUC4TfzTb9NZRIjTkWGHSYlxLf6b6jNCx
SYYbQ1XEQBtmKbEeXXT7h89KgY3t9zCUPG7FdyulgGjDaEThZiE9tYU4f7+ULojA7q9P5QKpNgUp
1L3Q+/8dzBGg/LTE14kMThIjcpCI6ZFZivljjYKT7JJGtTnshBcLb7rFuSxKyzVXyClYDBzGm38g
w9XtEq7boMTsR4UmmMF0G/pUUlk0efaYDriJnk4Xvw/fMcQV+Tci1xbv/fsOoe+hV8xGJ7j5uU3/
wwOTw9ANmtNcIhDcXxrqjef6h3op/Smbxto2kzHWSJIVS8nK0jh9PM3W0W29bYBDxRGh37Qv7Ra8
wzYyeLpg2wGM2gpbjeCi8cr6irhOB5jC8PiluOVzxc6BfWS1qDzqYt0zcdtnT7KX2I95uG0SsrM2
cPbh94cVwkvTAjzUT1B6b50D+RQQ7ExjUUSoVGBwgntwoT8zChQQ07+S8Kel/gA8HLLBK3gpezrC
bx3hYBmopN5i3sIzv8W+kXjHGlVAzvQGd9cdObh9AKULuVuyD+G5n61eVdYK6G4FKFQxPhL3nKP+
Wa3jfZGuT0ehzSEsrmscaeA+E9pV92JfVO+kNMI7o3aQ2RdRkK+HZML5RdFMUAtkk8WRwQhujonx
UqRtlgeFbNwb5Db8cxjhSgJT/2m4/SVkTLXzzBP9WfedPaoOwkE9tRt9A7ZDXByi3m95aM72YYdv
AGQicxj466g7gmFsC6FBGGv5mFh3VGCyIJLev9TYXgyf1NWyuZkkNEnFCgdWTTnKIEz0hSaMTeUd
kxycHQpqareRmnMo8NBxZyjmhEg19NtPDckUFlYWnw2+biPNrBiFAHsbVa4BxYaLNPBrKuqtHIsI
C/hhe0aJE8EzLBHlPr/eehGPmm9Nv66+xIR0l9+24/Q4EkeH5GorNjaUM4EAQAQXs9MwDgu1U/7S
Ycg/UDkk31vcbU6Ghw3mIJWiFsuiFe7L6qVS6NJzacni4nKvwnxDe9qjIXgsMTKkmbVbyCHRfE9o
xRQxpn9tR7Yoi5AVvtEgQmDx9GXGaGlPXVs3ntKR/Zg+m9OTeMaltKc41nivOhZ1Dje42Zylt2PK
oafZjEUnCPKzF/J9WzTI6FZCZW0/OZcQBnU4TObedCEeyZNdthpqUM2sKjZfSGZrdVEs0QN3VwrT
Hj8CVpNnxo2MCsRG6n3cwKveJfliI5sRBOF2OK4O/k8elt3IE7X28LtvnOcr2gfrvypL4ffmQxeb
Bp9kHMIAiogVOOjIhHIFHXm9n6fBs2cM/O52DlsuVJO+u3JhOgi8lOKVjHRakMw+A4xfKl2pcsDb
p4/fuCw8+95mtesGaEhqVFwoEDl9zXo3PUyaRwhBet5dkdzyoh8CvObLY/3zTYRMBrq0+6BMIfIJ
MhYB/PHCfCWMm8HGYyydD0m/j/SzMBKINHUsvxPHELmUzvL9rCSgh2MiGMiWjlv5AYWpcih57aQQ
00mSCZIrmnTz4HCClw9SRAUfUq7fVKFwW/OxUVhBKknhDys0x5CS5xBkfsaBJRKYQUWlR3rXMOWX
BpcRRZqlinGZtDQ5sl4QAoSVv4HoPbi/dMtEGQXMM1aHvBFhihI4VZ7av/8nkJTstMce/koxvcE8
bY6RkPDqmfOWVetoKWz2YEkFXxDTcVqldPDovg6pB1eKR9YF3va0O5p+7A91K52F9AI74/RKlyDC
SsIolLHJNCPslm7d0aiGjB3bNbRGHQK3FSwCB3dE8yfVfYN5b6H89oY2EP8aFYHftd08WiUueVBm
FPNg+W6M3TK3n/+GPEAwLJV10yJBY1jti08UoPz/4X5YMYxb/GU9duumdFi1C1TEzXuxUvLtGRPz
fFhnH+joqPSMKGyKK77B0TLL3SVp2DV8nbStzWIe8FKDS+eGN4U0Ul8r77Pfh7fFNdSF/H/uy6pH
IKC6ltzQZi/PbiRaoqDiGEzvkVoK9nYvzUWy+0px0HE/lKKrUVTn5E+VczQw3JwWa4gebkEwPsHj
PiA34eI4+m5PfGD/6lX2yKXch8lZTVxXNMObw/4GcWh757Pr0UckyVNdmTeYRIyb3ruolEFJSvmS
oM1n1PW6qEDqtYTxIDXpfFsd/vONTcyZHtEU5e6Y8eo76STJL6f2qNMye9nWmbtG/hlARd3x9U/3
11SCHql5vYmYhk3e0OUYujIOoIQp/WLYyGXKFl0pVkbOlHsShCck9hWW8BSZ93CAbL+drAqNpeqK
07Nl3F2cu5YS+WfcNPKwsF6dNoV693qZV3Qp6lB4Ozh2vWtfBBtKGnP2DxyrHgDEo4wHaGcqI8I1
sSYAlr7a02A7xJWFA+LOx/Amimj8H1Kd4gWZ71B7EeYYKcOTXw4I8M4cHfn5C1e9UOSbIY/hl1CB
9voDYw3irpFH4HVFaHG8NFeqfQSjn9fACgFigB72JhS0orvQC9mDTQHMXUvjxddxHVKbu5kuWf1w
ZTCeMo6CUewD2d0jCWcsGrXQox4qP1iITkp0dRavfJ9vIuFCUsGI6kshpFaSdDWnW/S1mLf9eboC
6Z02nNR0/7EPaEJ2/JpBCZ2/M7Q8g5OI4we2k9rM6edWWuvy65ZToihukgCFCKJS97ZSeXWH03aF
WgimhTx59xcP0TsA+T2hYhiDE5BzQtMyOlZVJtVidCFkDJX9JkHkm2yMEeaIlwY0L0yTk9P8lAUe
qcZzf46j2ssYBNPlz3+3+LegcyaZMX/BafmAji8zbPcRBXTUQbMM6hPvh79oWPc4fkYTxzBWzfrX
33gRYuqkdOFh7n3cORSXNJ9yLw4pTKtstbXwVsg0lXnAtZKBdSl0kj3MASgjSwUXh9Hx75xfQtiv
dHxk7ZHisHgiN6Fkh/yRazrv4lsWFoapUL3fHNlj/pFLDBcT3NPLkLzpo7kfo0BdrC7Tx3UtrzOJ
z8A5dcOdyroPYFWaI6kjZjDeYEDIsvbFMlSrx78oQYIrcJ2oK6ArJ72aftztLZV+NF/v+TZNGADq
xjpi3VRlHb96qdCxtoo/LxK1vFVngY93W4Xw79XSwSlYSqqTHCWhW8mggv1IuCXYXzLdDQ1MKl6s
rD6n+znuPZi9mQGOPrc4VDYckd5z6zW2k8wKYJp0LE5HhZOsqNepeYLEhfni3sIKQ5cwIDYMjezc
DBHvA+akpZ1r76jYmEW44k6jRiPdV3++F3EcvEgtFtUn2AxdpPNwIv38jQadRhDmmrVbzK8vA/j9
6OszyXEbC7cQ/1AaP92nRUNUygZZ0kVlCdx70SbFCZTw/TNKDZP4gVtlilzROGdkvkGmUqHcPLdz
/0QoEY2cSiTo/g1gmNakONsvMLaXTE4S2k21TAth5iWMZPbtfn8Rl0ZTe1RbR+cG3jivhguFSmiC
bt68oox8z56S/yYQsunF2FGL8a8HwqROTlsQKS8YZV6LNvNnosGJamtn/g+gKC4mmI5EpQIKxNzy
OLQpOLvCm75ERI4MfgPmN6CyuMgygGqAJexx2aNYDaH4MW2KiwWJhw0D1qKsVbBx73lTrhX6ig43
PA+AkctuY4MupmrASZK82GUmORAICUvrQ2l4AWPWglFtDzWosgs8ZQh0dO+DdsGvfzyZmzUOAiFm
n1btqW6lTwA+EoH7ODT+EmC6X6dLJ5X2TBK6Maf/h8Z6Ba6FPjY5+7/TnGEax7W2RXOCxKNoAIN2
oGBkck2el+NAgOh9w+fgYmJ5o4cRMvxSpNgPNk8pS3wVm9dfjB7CDipDqybfzP2JDYfIkrxwmG7y
SqMyPlxt3VvvPJDP8ms/wvwWSy7z/avQNZnhlNpP6eZnvchA/eed1hYrwy+N9l38bFieE3I0F8s6
gJSE41l2TNMrO7Y4AYKiiD+rx+FyJph4sIQR/iGZSAYrKS6abPscjdZVK//+tltFPbT6ci+dNVHj
VP9pPC/26bpwjtfAjvysWxoYqx/XsJzWfXK9/roz5ReCThckzFtsZ6WjMwVkPch/0drILM0Kg/47
5XqIhskfZhBo1oXwgtZ2JAG8ojhLY22/njH8yIinpo2Xt1ys3cBS9NdsMBifhjQC8OLW0NEKUzmC
+W/CMdozGecLdi5exkUmrfrOBgKZrmK8g/7iyBSnv2Qox4XAZVGHL0RyRGdLs/j26TIUZIYQoH+v
D5IHqDwk5FwWaEVJVs+NvZGS+2jwzVzEKThReAfZmLKwOu51DAzm7+d7yzeEv//neb7loEWxbXhD
1Yi1JbVRS3RNLF0ja+M+0l4/6C4ft72NMPCP8H54j6a79DljuM/MuEaN1plsV80rtPkt5tU/p/dx
cvYHfQGFb0X7vHBsHHYPRnjM2BX7kCEPLaZkVd7simFESKT6ASyCqDV2qKiw0xjE/wzAJ/V6NaFB
c+zijcb55vyo+tQ66CvvjQ9g256A4qmgN5hWxjN8HnLrr50Zdc/rgRo0SkwMMPKUKFYRgH+tI8Eb
Shx1Xuvq1Mr/XUjes2eVyvCSwQ+K7jtTgAqBcSRWhuykyadhsJHV30TPMvqr7U2QO8Z7wGoB59ld
SvTAB7lwY34F8neZcKzry72T7WooF3RZxg6u8UoqPYqW0QQABReXKUfgMTHyxD8LlxFGQKguMQ7/
2d7xY0J3yxBXbUwar9LcEOFWVFuXzzNmBAgF0V8+f1M3Nq2Ft2BSP6cPYrd/hXqXZf/nzEsxPPdN
MClkC0sSDKQqUeIMq2oW+jQk9EoUfsKW1jHrLSPQlU65MezX4IsAb1NRMJkm3Xc5S5O8zwhXyEXV
pvaGWQUplzQtZCM+CgT0UV8dVtDGOGACys20NTA8CJ8LRZro/EsxW5X4t2KnXaackKpzuKGhx71A
qjPIRuAH7cWab1tE++W/aPWCKHtELWp/f4dmbqeEcR2NYva3MV39A/Tkcjrr3qAEgEgjkYtjTxzn
0XghUxc+cz0R+731Op0/SvnFkmU6wXzFKaFu0/KKPIsIK8k3gxkuYXP8dovHYg56fCo/RmkDJQlg
RoWs0ABZ7t/fGewQ7UrfB1+bOL8YZqa9ObY34o3gwzoWvJ4MN3WWvVJwW3LiHrl+UXWuJAtPzgcH
Go+AQ8ygDjtsZBEKt90DRudhXM47vv9jNhxbQ0GZDyGiD3UcUmXWyWABySNDYBvVpOIq4wPaCdj/
/32UUpuHmCFLHSp4fSTRT9GsR4zASfnKnvfhokhVBeo9x6O8qfYD2IoSNx8hdyA5jcnoiknEWGax
qH1M8tZstq64Q7B7S7lG0L/GB9xqcU3Nr0kXO2GcJOx0LM/UCXlRW1ju8MNGg2pYuiwJJn4ZI2hD
IFVnuzF0OvR2Izk7raoo/YmTp1NQMzTz1tg4zF06gsxJDnMprylXOPpQXxUw4tMLKlztzZkFm0up
OdGpXtxMrxzlQy98m4z9oShiw2VoctIcByt8OsYZ9yTPFImmV8rE+0bn/TF81f/pZgEOXAYrEUGM
0tPr6ICgHOGx1QelaeKcoQrjgGdE0ZyC7GPeU5a0Pa2wZHqIlmNF+C7S776lrRsR7f5Ku8tIo+9s
sLxYzgZrRnjpM0YqItoy1dV6gp2RXz8ZJmTVNec3ufllLpg/zOuc4ek1h35IYAPxOKAVE08mgFGD
vNiWUqPyE4OOZVO+qbniVB5n6uJphVt6JN566uboOOUx7RjpwTq9XY00WFXbz998q0U51lGhsifA
Tw5UHYKqmNdSHBuqrUTvPysc0qQA7gNuSuKiU8A+/z7bHzRqUAdcT0JoEeJ+P67Ua08nE5qFiYVa
cEStoH1fuwLbJXRGQMvhmFJOGhIYgp7hdsx5BMLnsavIGd2K85EmvNXSO2LHKJBkca9KXY4Pqcop
gwsfa9aoBem7uaroGxPebjwCCG9DekxGffi4KMs1UtzMLT7Fb+696FHqoMWPEitKuzicM9p581x/
7+jfG9m5rbkFBcXVESi4iB0UbS4skRxR1ySCmd4nL/JhQYviJiRz1lkCwhD9zr8xf2fWqCm+zDX7
3bQM92vyHgRPvAeo64MofKu7Wa8w/+7ex07vwFJYkwhH0Gjs99sCAudhKnIvvUF6048OB7tLJN31
lNiNME6e6MKOTS/+JPo5T7wY+NsEJXofi81OEmJpwr+xZVUZmG5yKlj+25MruIfxkATDR4GIAmUY
YUnhI50QfZoDQ6dRbAV2re05xBZdFuixPT3BjDBvqQMZAUjeT1qUrf8g7aFx8UHgJWEFBn/j8FsH
BOD87N3dqt89UZ1hRfnQDjIqVM6Y1Vg8byWMdeeOE0I5Siao0DFR2ogU/oNm5UO4mUHD5+QAYo3Z
P++AndOz3aBjssEbIqRfqdS5Qx1cXult194PDv57gbFJkwFYO+seDshTne3BiQRBlWFVS8yvqjeQ
+NfmQybhOSDb153d9QMAsFwdZ3yDZfOFW3YPwQ+0FqF6D3YUTin6DspmOpHqUWBv97OUUVSrJ2wK
A3DFLaenSJUUMVJCdQFw9bf2vrluNH7MvJw12sZEoVVntSbBt4h+kg5z+LZLw9MNiYnbqhxiXJcN
oJ91oECqgNWcmVzUPRSPEk6XCVh6NExj/eI8ZoOk9ndQJPrFFtYCizkXYk60HuB3Iqsv1A6yyr8x
2ZJfWGb9qhp/bCJttAfYTm6pHL9Vz+azVAoRo7wkYv92MZEh4rp9qLr75yD9nyR0ZtfOwr3Yk4J+
vcd/80QVhXh+gc9WGpqlb9CvpUTuJCDDj1OFk/2vEA5I50pXXZ7/mjxJ7Qqrl7t4ttTbnZ7FLvUL
o96DBy02sjXq9JBxxlLHLMLBCbFVwKgeh4ZlAkXzwRikGXOkBIR8JHYj2FM7DxaYaVoQQpiXpIEn
7xI6OCtCfA6CydDPRsWgIc/DJ5HWLUYxc1zca1/JCT3g80gaFknRwfU597Bv7p6csCUSqFIfDKw1
vfDXwW00QGBVzpUYeCc2TMpkgYB8Cf4JHSitrVVUsPySTS0iA8NqbZGdXFEcAqDKfkS4bSqPGPiz
PJCkQe1wURR1+UIctK6trfEctA/1kZuMgGGLv0mPcpfHBhI1xH0YTA9hqwezLc44c1mXwxxpvhrb
U8AMm3x/v/tJQLqVlqFos0Up5Fk6FxYZemnVZL9U2Qt+Z7oqxqNkjOywsxCUMMxPWBjXkXtXjxt1
yOrNUtJweuP2qMX61OTbSV+r/VRKYGyJB/+k2o+GXmY5HuESAxiRP7q65NxM+iI3evjCzWKa3qz4
Wq+SRHnY8f18YuHkh7w6VcsjEVKC6DxAbFnALzbZPZVVaBRHngMSDpfUKf9DPZPGW9VRwr1Onyob
3mLnDOrqOL7H43eIaXjHQvi7hZZ1PlptyHUNQpCrOs+2kHspa3W+ITrYkkXwoDtyRDiJ0BjagbCy
p5T/NKSiQ5yCvUL1ZZb81skPi0TcDPmq30D2WOL4K6FA2Vz7yXvwJIYVwVflkNaoOYs9+P+EMEEu
GY3CYLLfEI3XN5IYcIvWmuzt+0gVUGdcE7CQW5Wvc8lGGYhd01e/mfE7Ss7bYl+MKQwEYcVhGNKe
zlASE4wbeGKSfI08T/mX5EqEJ1HdTD8gYtmK+D3NknDtI8sROzBfJFrVji52UHe7JA8/4rBj4g7e
pnfwvdDBfu1+yXT2a2QnHjeJBZYP3hayoGbBAaVqw/60ozDf6B5HMjYmlO7y7vERMhkUcwtftiPc
vI2k+XN8FB+NG0M3sFYPZOp3xb9G9nLUdABK9MMqHxrVX4xt4mOyJ9AoL28pNfrCnZHQueLvxNZg
Ne4KAxJEdouzP5jnwGrM98OwAAJQclmtC0VooBnbVkBiP96A5wvPgcEJ+FAvQ+4WA/G6uz3HbdYX
USSe8YOW7yUUk3r+kJRhkzE8/j0357hcuM6S1Kn0GPR6ANzfM+9tc47lyJyM1eZyEFaLMER/LyDd
2zZihI6/mQ+Z8gOoaQPoTMS3w/glHu/VUbW76OcQMARh9eqX8LBO5gxej1KMbc7UqNl0LVtovN+x
6B9qMqsJKYpSPKDa5NdcYuQgOXrmHdvyflRMwaRa9XKoeOZooYuaroiIGz2Z12N/ZkO1mR8er0Fk
MeZ/O9tCC/rG5R6Ik80xFPNPQp3/7Nn1c4F8FtOV92zm9tPDG97h1qfAfxQbVH/ampjyxRhirXpf
ZMHFZwzdVU6xqQBAp6UosZMy16wW62qx8VtrX604haSWjyPVVdDT+DskcB0gwRGZMTtVZ/xyT7gA
ZczeAQoT6XEpuhEIwxk3T0JNt190T39Y5Fcn3x03N1E2AxRhb/KVYpvmUNlT0bED9Io7h5KVBWX+
90aaXWB03oRdQkk0ukV9fExypvPVR6gciRnebu/ci8LO0exQrAUECHgeKdphDo3xdbZSUdwUXzPE
4Ep+0bVv5ZjrCK1waC/V8MMBUOLKSVKkJDCrtG9fSQffxIXNhtxJKMkttWs0p5Y36q6b2YFEx8iQ
Om3zc/HVqm9W2HeNVPbrLpu7vRgzSF2pTTQkQLedn6+woEL7UTw3BVwjJWZZ3pHZkuHtAjJ8R4gR
NbuoHtHAkgDW486eSAaWoLOl6Kcs0vjYDr2tLafNbHrd4zuuet887F7tiUlfFYMHntWwQgLUstVS
+3DKl+9UbJTqLWvZJKGDgWKGTv9CBsF6L9juu93ntZJoEQ1ea2c7xUTvjzkSyhDrS3DaC69IJ4Fg
I/9UI3egm3icQhOAg/TmFrcrbvKJNPMiXjw9YRcJd9n/+K1WgrtB2KX7FMGnGs4xZR4oIMKUmdNu
nMwDHt/RBidMQIF/8Vmju09exgozrEaK3ktHuDo/5lqFOGg23TotM0P1iYOPRfwRzsnU+Mfkvx6B
SF4MhMZuI23r+Bs7fdJJL0B5yAKf7I/RHEd6FPCH+ro+9e/SGkaXjqVM+H3T656RXcSp4/+MBk8n
LhVqKfMvGTFKpR8m+6ckKEAgr9oOVd5s2F9J72c1eB0agXixBfD6Fq4drEmK09jdpRNdUAbAEkNP
Tf7yPiNy8BGLxJ9ca8scb28jkUxXfEfIONHGX9xpPvRBJgXsIrwKtGZhjB4GMnUQgFMRKiHTUC6b
pVGPw+B7IXAETDq33W42D7i9KzorYwSq8ah7TA8Lv5ZqnOWXMB06zRaR4OfIBPeMZd3Em6n1x/kq
24VYiqoJbTQcO26SPgfVuJrY3jKHiF5kIcvlaH2TaLg6nP6juMCD16Lfp5+XrkHnxrB+8n9tlx+0
SggvnmRVsqtTMRZjO10xioMNeKhLZQkr3t4un/GPJtbvpDWmZVFD5m/2zHQnfBm9ZsPcAxzQwy5x
kxUeT+WCMjuqLxKAT9GqUTuLZzE1QM9m6d7p/R224VHkXtF6k4nygTol2vN0EG3UgmB3EqnVlQOR
fytiZdjkquGabJi1LRMJ4OdKBpQb6wR8Y1XQUEAit52ve7bQhEoE6PTxgdKMB9I9gLm23LHQZ4UG
Pnldp1b9gEIZBrCYzCxzhH/z40D+YFI/5VZu9eWSKCB//SdzjAQL8A2TBFlIqJVuZ1K0T4gwnNMv
nyQqOW/LIn62LLp+b6vuKOlU8NDgEWJlF+3f6k2vPsBC1FH0W2lXOSboyV6EZP/EcPWcSHaOnEr4
/dD9sZ8a18AU7G3lyw8+I58tOz59MZFZM/srR0FIiFGbaPwbFzIeeb/P+fWKG75ilSvnWemHX6jL
EIzNCV0yC+xW4EfVHd8Mh61OJNiM6dg+RdmkrFdaas6OpFLOd6hE1qYX45CDxCDkkZSw0i/IMezf
zTEyARAS1poHz4Q3Ihkv5tfe/DbfnjQJWfPa7NLGLlZ1ASVVuRnIhghgysPXvPKX0vAFxUjak+/G
ozIbK5zGMuEjwdhXCPnHDM2Lb273Lk+yhuRVuY+A3Rmde84D/0B/QNA6m4b8LLfmAWb4EynTU3W3
K35M4K1uSbtlBjv0NRZC/x44ZsDM9E7T7Jz37te6ti6bs4T4kcWiNM6b3utrj+hOgXE02D4lye+m
BK6XqUJyIZoH3grk+xQvSSnNX6ei5AO4tE5rJwEWIKruwpHiWN6nYsFC2qiflvAUKYM1Dw+vgRYI
sEXRNTHNBdSuaek2dBHEGsqe1fs0fTeAKkx0XH4JYrSj3hmMUZLHKCEjihZJGWT4/C5Eb0H7Em3N
1Vu+CjUQkvQ449r7WPpPe94NsENr0ZsXeqUWjD5qcpLBD5S5w3dozupwrGnFzZ9OoNkTr7eWDOmW
sVgaARDxomYaqObdN2LpGFoUm9DFJGUfoct6pwJfVLZdJtwAcigH4y3Vl2kIRGwAo1GoCIqEjieB
UJ7B+vdXVP2XP28fsK3tmPJ07CMisyxWvcBkUUQm/hjN2nbZNs7HOJxv7q7TIEvxFJLCxrtQYEVQ
tAUEl6mIROWZ1Kx6iDK0XMjWqKfbz1S/y5IIC3mTmfkeT89lfhbMd283NP6upXfNFhnttofrau7b
2TuN6pb3wGy5Sz7iV6iIQdA//ZYasXSyXoVAnj7Eyy/qUVf9KMmWczq6hphvEtXM9D6zcTTNsp1h
Xtg8ad/aj/ZFNimpJTGw+xHiyZnsT9PB5dK5Lk6n0R9ZX3PcN20svxkesSTv3ey9RsTUUr8teIrE
nMas9jpthsvM9JHqqCQiXwod1gNTSTXhi7IcvaJeGu8ePQP6iPdA4UyN/u/kgggQTRmFNRS1t9yJ
MAhrWN0eqWfjSa2o1XGc0cGB5g5QoLmbOLIr59Y6eqOHn2NU91uRdtE4jhstw6frh6BOF21Y8+bR
nbJ+jPrNLdjlxuO+w+GOrk6jTEMxSdHwLadf/IOcu9+p/A6OFz4J8SUWpkxsG1ejcFHg51Lrzhec
akBIYtKxGjyMrqWwNor0U+2mh+LbEl10NAnsuD3+PWMMGDEEi5I4Fsy2vJrt0xCYfV6n3BkxMVrc
NUMeSywXGs86Wp6tbhinb2INvakbNP+BkU+9K8SYIBmZno3QzVXNPth2WU/qud6kMyQbQcTQx3MG
LoaKdZuNSNkL4Mv0ObRteICICsdaoGpUhYrJj9piYDzvkGaL3niwDqw/dBVQSIElu9LqfCTtuk+g
X2jr+8zRT4nfioRXX1fKXC1VFFS5oSdMRs7zSeGCdyKxa7zXhvdgrepOMMgIz6SQMB7CNNHyQKbi
546QCkW1Xf7zd/4937FOm4cI8JI/yrLq1v4CUWbAVKseED9eUl/Evwns6tKkuHR6dOFjWGQRbYIO
XXmtfPHY/kcGKH5f0vDYK0fdOPwirMh4GzH1tBMXQj13xVgLH5bl0lBWkMdlgEovL0tky3DKTP/N
9LmAy+jt9M+FEp/RJZ2p24MglExdFTz5IFpO+QKd8VTh8HA8x2hDsVoYr31ep58u1bf9Yk4fQIHO
bo7URQVnwGCYfAGJSQkPh9Pur4t7omba3LQBi1J+5/YZq3gITOpfLNPx1Whrqpw90A1g7eKvdG1R
v1sfqq211Ep6JXX6fzWfhdTK2jqsqdtKwKQRZd9HPj3Ho7TmjZx+Y3E6EN2DZTBs2Qq4TDuDIuMk
71ZX9kVLY/LLqLgupwgDEMVFNa8Maz2EOIKhlRP6bbLcdYx73VZqSPMLiSEaLYSeBHhf2Z7c7WWh
SvVOyi57LpeT7xVytvOcGrNmbOXwLdcfM0WLeJn1vJMDloFHO38riDK1S5jBAaGzmob4KOQOt3OY
KsGgt8KTnS8D/tBDUp1q8aiPZQyiygFzND3QvNzxtrl9GV3h0aHcAcNTv9KUm8H25090sSJk9zgb
FxdkvsdDONvm8rU/bOSwSuPBCByDNPn7kCg34dyhmAaCtGXQ4x77YMc4KXPKRsTXqCRu/Kr5du0L
zSBoSvdeyZuObp7YYvK3xghgO6rzNnYgWbtxKhq7S11F4YCk7Gig4KSWs74CA0IMbihTVfuWfED9
nJU+lVxPzU4bPx5Zf9puxSDWNhjSsm25wv+XIc13O8o23XSvHDmnoO4SOVB6waEyehLE8arwFcl2
oAEIUfJrc05ckSIOFrLB3PEhUn8Ea/iUOIOjigrGuCM4wOoIrXmj9/16kjDk4NMybG2TB11iuLAv
gcCjEUYtE2hw7LAQ3uWh9uOqelJh0S6Pgqrmk1tBQYCrt6eJSl6UWfFSKHiy7QOBEqY8Zbi5JKmn
JjCNywuOHB/uZn2SwhSrD4Bb9APduNV7TDPICIY5i284KK14s6JHsleyWcFRXUVJEaRFh7IW0PW0
SKQU4/MK6oDhEGkTfQ7OQJ5R0IvAABFTD6f67Gup+2ijLO//Qkz86xYYaF5QlQCl6dBQ6+XXGJnM
5M15gWBRA8rDPvvXpAzEboLHA1d0VbiEkSo7di00GmXzsNtsXOlm0HwwgbMPBWlmDn4b1KLNW5mX
PBamp1LTwrLxgYy4gwh+jlxsfBKKEosF2h9pfSZXeUUUHCPJlCDjkWP9wwBf9k4AKJk9W41M35wd
IIKe92GYyN7tosW4opYnHNyEUrgLsMqGWnhKeMo6Cb5V1w3SOGj2LOGYXLNqhvLSnXp0xML/N5kw
1/OXKbZfvMCvqdmMTkVV5s7SU7F6tc8Wp2KXB966Hn9hNRxHKxtBThdvWAKt2JBTnERvRsE86uuU
IsfLrPbQoQeka8cvh+1O9K9kiXjmAp0DTGV62cWt3YB4WqJYKmtst1kxlDaPbeHkOGFA2J6bw+JR
xLhUkr9D8co91idNTTVgSIBNh6EdnwB8u6S08krCxOk7KT3LoJRh049CVZMOuY31nKeq4YDkDA7J
KMOXcjhgM7xJ9RP2vzxjVVLhz5bm1OCm79BuPD1hBeHQWVA2n9eEHKERIKAsbKHm8URuV0mVzI9i
JGoL4w1RwG2L1V755MOauBl6pCwq3P5Uojgygp+l+X/cFSKKZOnC97RMBprgLEo/+3muuCTdJnDq
FjkYVWwtVvymB7Ps4gb7vr0DDpyPbUYQiGgvlTD2dqLzxJum/GtawfK75otf91e3Sfz7ZA+oPHW6
xPtCpmdqjPAhEa/sYu/OHuiDd+OPd6GFhUFNsTl7o0B7T7PCEVAeNjv6uspLaY/qNQPekBV+oVxv
y83uDuagpd7pxqyTKSJ44/tXcbD44akJxiC69DL9IQZLkLHmGRc+bC3B8P7/Lfg5UdtocPto8gvA
Vze0Xyct1c0N5AsQDqLTMh0AwZDueVwuMtQs7NCuAdjYbTM8+o/+kujPaWa3wO4j/6+WcycAe/0b
RDXlBjGrLAtOPy1fcVAQTsPI3Es1j6ga3D2xe2p94STRT5ONCbvwfzPHBcYcCQzlku19TrQKZTX1
ZuKCCE1DfpemQQ1CK6eXe2KScCN7yceI7Sh09n7FXZQeJQE3XG6pBra9BcjfmS6LFul2FUNpBRk7
ijpTne9qype7ryXRuo3pufrtY7MPsswySmNj9NV7PpWHZLRadwjlv5ZPHj0/lkel4qlRGc/WU9sM
ZFBNnzJIMh9kGRQs3fycj6o0BTbrbhvm8pxyGqwzmU3/2Vfjj9BJldc1wnurmvtbkD6EKSglTLzs
0GrAHZ3mvkuXbHbMpiQXG/q+2sNdStGHAEpaV9dENCvgmVpudtaUc6jcHsCDVAItbZpd8AGRH/F2
ydylklVJYXsAM8xUAB5jpgMTMN+s/Tn3STx1MDq0OCiDqyuyVUZxQynhW/ZG5+EDRLw62o981ibj
w3D1g6an0cZ+g8Sp3UZXirOByefk2X9+Xtf/Pg4Q87FWBpTemOcA049b6xXjhR9kOqn+/Ks+rvcf
wztj4IJ4y6dVi1vIrSqx16usG/nLPbjl/ZsiPYPe5JN78ogynrOvFL3k6iLsTkFveVqxwvkA9yvf
FbDJKcjNJrr8u9ORMlAsrXnLG1+XsytKW71P5F60R43DqP3zuIf7zYMRfSRx3k9IXPCpsW+OH9yx
LVea8WIMEAXxK0u5yImjshMS7NzvHmhd/aNF7rhMoLpOFB9Xfq1n/bUBG0+s1OR2h4bVfLfblqxl
O6L8QtoMf7p7/pMFvcBfTlIciHe/vptQDBDs9XEUFc6Xk1kHlQqlLgpxjj/LwZmKCcitzsTHCdza
270j2vGplmYVX6xO67p8j/Jum+Rp0LM0+u4sCzV/fQRflR6vSBdxBI6zqcIyZfUJUqZdTQUiAUxS
udFlVC9Yjal7GcFvmHmN4kMKiR552Tz5sO1q0is5OxJm2YdsWCKPG/1bqMVO+fyDAGF0Ngr0iuan
orHOuY+1RkV3aYXjlmPaUo/vuKQ+3u8qVmZFRUYZAv2ung6T88wZaEFWLX8rmcLGkj1gvtKO37WU
BOJG6tLtyk0bEeEU133bp7wjdr4F4P4oZMMxVyCpsU/5AgKSlG5/3gbKVTqXmygf80l5gwrxouPb
LMekXm7HBU4Z5ihQ3J5Fz6chx3Sk9t9gKLWjzzZaOe5vmPDO5Rx/styC7NydnVwMtmWF4qlgfaMD
+HFESICnqYpnkKGeQHjMu7Pc+v8Qzl7kz5SWHGG95RHXG5gTtcvdywB8n+G+n4vChMKh0o+63kQS
mD31mRs14BKVmBrHFG3vp/X+Tya6Y3MuwwgrXoMq9q+0ltOvR38YzmaZ41Y3Iruf0kjnivyYi9RP
zY3OadGsat1VZ46p9uKAJmxZwWR684WVZJgaB/FC9zMfFu59gaEGimTLIu0jkk065Z+rwSkDPFc5
1yGnOXCgR9BYn2AYNQAeV770uvv4mGW1I6qbq58fShf0QS1NJPEXuzPwQl6K1opz1N43sSzLBg+H
bovlWeNABHnM37cs1hEbNi9F3rx12itXMim18Ost5hRqcM4ldtEz7mjlXXY0tKJCQzvgI9ZNB1sz
sKGfQGApm+DL82/3G+vCOeMgtLuEU2R+/Mfgk8cVmDFNHCQ5oWTO/44ilYfADPwiw1zgiurB2bFB
7QPc5Z3xrPI1H6REYNL9eOo7E57VP6yf+pVVBfMDApUAUa37KbyGxdzj8QH8XceWdR4kevVMoUCn
gR1I/EiFv0d9gGvg6i9oeHoUTzL+kLGsOLw4fBVY4vUatq8iM1dxcX4o7478I9W7E5Y+sQbRK4JW
A4Tmo9hmiK/+psJeQKwi2oaY4j7Vo3gzCTnDSkT5XkxzJMgmIKwWzcUepxKs4/r/9FCMua4w8mIn
xO0OcaHSeYy/FMaskvqjA+yHJSv6FB1jFUjFztsKd3eTZyXUQ/oPw/A3LPK3fHD7qxcwmKODnrIh
PggBNKM9ZHlbNOpJBMkt6nGHfoHBaXmfHqRcq5GTRAJZJolmVTyifYPqoBn6q0tnO9N/XheAvf5K
35ZHzpzdTOnDT72yXaryu544na4huoAAHVyWuG5cx+xhSmw8qOtQ5hrlCldYO1d57R2SWLVumoM9
y/Kb/h6HXypdiCxmRVtZSGCej+rhZRchi7FIiIyPLEWJAN1ASoSQVZwH9H3vxcv6Qv0m5RnO1BS3
D5Fs/44z5FrIZ1LWXtmc61VF0lFRV4slSbfb4Dqd0ElBsUkWSDR8h2JT7JvCeZySvgwXecY6N6h6
N3ruoe3hP86icvmOROcMqIQw0iIOJGHfFgRigCl9vEdM+ZiCzzqO+qrMZSWgVfN9RT25k44IxAVv
8VnmlVEebCKtqYdI1xbrWewsXz1ZhPmxie4A9h7LHIsMNHsYM10ZoGX3N22a+4an9QMKAByEMWph
kfT9qsS5BurWD0fOA0iD1yJAsioOewfE6BgFpS95iCTxXZ4dxJ/NqlUkJMT8yVQ594ZYRigqXvKv
3fBHggMDG4uVf74l85v6Z/ANkRHBeex1ngCrUdEeHAtAtTLDkSnu1HN62NelHHXk/6QhGTfITpnW
FB2vJnpNkGveQUhbeSyUvr5SYEFkvj78QQ2fRgwVYBMX3x0i4fcQSaI4l2iGhtadpvRgogkFcHx1
2Sn5wZzctH5/kvhYs251MtGufbb1WpYAdJIUyRF5Dn9yZNItTvcQLj7hmWl/MhjnpRL4w/O1qXJX
RGEBjXpwgrfeIEX/DFK53YOP6P6STg4jiJgQK5PbjL1Q4s+omomqmribFLPvpXtdJ/nGw6YGJ1Nq
04Z9dvrtSM1dX+PiXY5IDlMt/bc3XQ5qJNAQRI9yhE/fvwgU2Mp/amzywMUu9T7ux6+WHBIMYVXV
hpnJxqSJt/q89UE4egKges/C/977ER5fbk6R5joHl30GBkw6qcnnZnMux4fDOUhwsWfUBGj+m9ad
nPRI92Q3rgFijGabMPRCjQFr6G4FuxyH4cT9JlSqanawtl6TmBuKcb38BT5kr6XeBv2eGImPGbNz
7bbZE/+IHceEbUjNbYun3MmY5KFpH6We6V2Es81HCIIFXDieHJaW4zxBkMCZkLMswDx6mkGpCYKs
5UtTEBK6m3Ppipl9M8qTIPM8/7Y7te1OG4fdk09e6tTvdxYRZjO/G0Rk6d35fzpHbJtT3DUA1l31
no8mCoSrs42wEUrNto0BHDsg8esF8K1i4ZPMiaWoKbeEig7mTmJBfJzamRC72k9+pmVFO7/yD+Cp
ArfzN1Z23v9MO+DcznK9WdJ/WBOgoS32mcQqTlhflYdZ4hfiRK0+hJ6hCrf88UKlcf0L5nKSxvOd
bBH5lWanoi08DZ4dW4b6zoXJ868ay7MMOD+O6Hg8aD7UM0jULY0cQPZbTZgzQvGEHDUTj2DE93fi
DRoujtV/DcSMUvdg1UVDQL9ohGXpxiT3cKDuEN7qe9GSIJ6JY0lnFajOAhseUXUdtwx4jbzfwDnF
qpBrc5OVagLHNFJ97bXqFaa3qqjwZLbizUpi8Pyi5tDmr+yi/yQSmpyL+4+mOSdBGY0A6rV3cRmN
Tk+/ipvNdeiqj2lkpZtYzEcRTuRBRNvAWDO5WJ/d9h1v/o1JRhcDZ6600vFZgzI4df1bfp65iiz/
OG9KjK//EelH/MObJM8Y6Trj6KZEmIGyumaWD4v1zOY64XRjB8wo52i/2B4P5Pupa7TsiqS6lR9H
XMVx+V8iV59ThD7acXG4z/dMGuuYuGjaJaxxRplzslQfCva+K/BetO9kmIyHJUUMy0BcsTjcMl9+
brRs5rekzA+SUh4pgUzxMTz98lZuitn0eisCUmPbyJ8zysuu9oDSpjjTsbQUly6UKzdiVRu1aJYF
aXsZY8GX1RXUpp/iPxY09bI0xor6YG8XGG96UXzzeIEUnVJcpYJZdaZytnF4dZ5FlWN157CVm0Cq
GdQZ1U63AOwFYq9Y5VqwZSJuZu/akJ92p3aa3C5iXaAgKxAJiLzSMQ5jFRY0S5dYMfHqfL9gLBwj
rGbBMUOlz4AJ51c+RQU0CACUf4Li+6AZufTxt/gE2zC9ru2IuJWr7MyfQaP0Apa2ls0KQ9PsjIsp
Fugpd8rSLh38sl30PbbrT5JiLCHTpuUJfbzz55G2vIhP6JZmHz5KOHWaKhrOLOyRAQFBk6igQXvt
OEI7/44dk2PFqwDurb3CYA1/QQGbp0p8tRWr2P4s2FbDR4vpygwrG5mIhqPODcCNGCrS7DPz4+6k
rSnLj7rooIgARUHcbdDrUtAw0PxtRbdMJPojGHJSsny1nHS5ADt+FQjSbKKGeQHHJ4Sd6pT/TkOd
ykMhezcRp0HRtHXmtSe/rmNawj9oYcnFGqltNNEKfPoZGSTR5cyCM3sYfm2ZlIPAJFR2sS8/cq0F
n4GMSeEkF/UA5GUprgwOOTPl65HDlyvxlZQiUrrceLV7BnRRlz+SnIenKflMVHMuNIsn+aQ/3i/8
l0ijU+wr0Ai7aSgc80fgC5ncabGwxZW7Z65gkdk8hdaLOFMW+kZQsthZqWRWX3dXrp2Z0WmQwzpK
mW/Vs8KDzWAQAFMAtpF4q8qqxUsP074NKlejNl3Zo0uOSx5hbpar+m5cxZQuV7gLW9dDtz7bHsoI
UE6YLsMNC59vMdSntfKIyfDzFA8nHcWZMNNUrgmwj6ORFtHq4xMRg612rZIiYrkhs6jSMAvvs25W
Mzq+bNVJMscETVFpFjN+sG6JT7Cpl4ldHSRl31p3YETvhDTd/hJtJNZBHiFSZ19CbPDlpVLa9Pce
XYh6vIX/nzSnTS3aQYB3ksbGIKYQeOAn3X5AtMeVnNnHq5T4R1+zusYfEDHcq5gZBtwNWqXTcXLI
DczsgK8+uPf3BlukFhMpb394UNX9LYHmgtda65GodfCGG6Ehh6hxDbIozJYXI1vWNis+gZBod6bi
MgdPlZiH+B9z8rGJ2yAtNwQNwhB+LLZovkkNzrNjKH+EZZJFog/DhswYET/uMuiB47VauFKF8rEh
0PW8Hn/0/nK9vGtrLGMLf4gsRMvJRSAApfHhCaq+II1j1qrOH/ls71sRbV+A40qY0UlOh82v2oUW
YWQM936NQowbR999W/DRhOUubOaXFaDWZhVjKU6l+IWUNTNuI3BZKXZQmmfizHNKmTOP9xxYrlSe
ev/wBuexeQIVIj1QygxqQTbzxe5aC4LvjDci83y+00/b/k+3a1qtXeQUehIXu28L1sAETGAgNNta
ae67xcbO80SWVcop6GJsaeOG+kgt/WnOcIOPY1WqK/f/mooTCAuifrDAZmRb2tWSwpujmBx+jV9Q
1VDX/w49TtmbRiU9v6/4IX8kqBtnrfxPjOGpXBUSM9FdOEjDGneTHXv0UW6YwmHPaXY8VJqhw5HO
Fq0E2dWgbDBt3glg+jbuMAjDcZcG9YWM7Ym5kbGkRPcDL53dvYFN0r0lrytHn7c8BcxPWs3HjTJE
4a5jOi2pFUb+saCddEUnq0W9oq3q2rff1zXWc6TFrvnajLMQBUZ6HoGfsqdj9IOYGf7bDtcmZb/M
/MpNiiotui2kd1TtdDTAe47jutwQdPDUPK4GzFJHymD42E3lTv7gGut70w4Y3K1YOOo82YIgu11V
bLm6xfJJEKfufrQxhoTz9KLMdbhR8LqoqFWC2+ug8prmb5i3AplBKO5xYjgUN2Cbc/TVhuPfgaW9
dcxBrIiDW6PgHPY4EsSMD2rKS4hJKKOD2ft6K8BqK2VHyNcoeXGmnkn2DyIlG2hDOXCwTAktLt4r
Q3D8ELN00KS8jRHFevvr2x5KQYNkqwstM2d92xeAmnfqrj4m4khkCBT9Rd6OGrF255c83pQneSNy
K2Tg7OXVwQaQI0iIUzdoFYaICHf4z8pE5y2qvhMOSyDHmwr6R8YKK1zIGEre3MFFeUDPuRZkeRyp
ljnfVHVoz+e2GbAH41M+Ky7830dwm54/7BcDlUaQR4uXhE9hRzTpaFjHCzu88Y5MtTkN3fYREQXq
VvuUYkbielLtuoIoXRl4kr3HQcP/pr7YYBb5h+obCh62+FhV6zVDD/u9KIL1+z+fDcDmoeO6o8V0
/vNdH1f4YT2rSFIzWw4YnaKy7qgYvKc+hbrFLacprwQWq6RzE6Ku78WN4GstZNcSBIP2gcdLisV+
bvTiAqzxXDsNmKyY79IHlPealP2nCW0U9/Oz0HYs4K3qmGoo2q6AUqmtrU6ZoCGmZxxTCjqu+UF1
2BmFyvqYJrqchUJKzI0o+wi7r6dF10lblVuXuDVSUopKYL+Qb2QvKi1I1JoBACYDH8j45wT94+E3
uFi2V8RpQIIDexf9AF6kz03oUcamESz25+sV2vj4slpIB8jmaQIHgeF40H05/0RAVYephcVDHScu
w3BFoEHtgPcpK/AYOcByxPTqyBFjWVjB6+30LIRP3NNFzeN1GBmp6jEoUofxV9SU7Ycpty0fwPNv
3jJmdwDzWqmNmmKpCidOw2RRzE924Y/AnaO6OH6Zb1o546zSyrkEzy/99CwC+t8IbFhAuZQIlI0T
ZXg8xyeOjszJAookgrs8RfeysS1upvePduxvRS0tVi+f2mZejOPwmXUf1Wb2yDoRd3HVIB08P5TA
/NBWTWWHOICCuU0SbTs6M0SPB7tUKt59FpmUAYh7/E9LHs418/UE0jFmau+5OJYkf4H7tr0IOdaT
HiRoZgbVmhmessdDRD0rUNjLSX09xnzMn4IYfqps/1eT8LpWf1bSLrejxy8R+YFFTqma3zFZo/aR
zmPxtJ6d2V+T+6iBnwv7ZYY1Yi2aVr55Ja7NGSrXLxpOx/cH+WIrpK5T6TemSGp+hPR4dk7UBrdK
oNJ5M0/sHHQwPdAWZCds+/Gnt+RcFgxsEgdINerd7l8kSZ+0WRXoVqnJFtEAoC81Ecrx9KVeDBGf
MUikc9PV3Kq9SsvRfmeMLf7Nj4mJ7vv74dDuNYicAYMjx4A/qFk1QlrgklkE6yVUs0T5bRR3tK4u
l/DYK4Idq6gdokJ1AAEPaji//5KQvq8nxGku8YQXK/cYdCp9EF2Es6Mya89wMJTSIHNuutH6cSW3
HOELMjLZfHZa6qWEvx50ghZmqi621tJmPOO0W/5RdSV4FCxstK850NS6PwNniowl8Bpx69BP8kwk
Xki1J7ns3LYEdH6lu3dYjGOKFvYhQyUoaI5csvY0jMikMVBZxcqc3n2QJuuPej6yl2zmtPGnfN1f
8E2fD4ZpNtB5EV1V/GA6m/RteB8W8Z7of5JjBewIuXPIQiAGfJOYy35NwkfgbMXuUactM9xAny49
tF0EAGljCAMsYb3wa5t7uJe+K+du3pg+numYbI8z6YZaiC83VJGWPilWpcRPPeXXj2hleucjLZEY
e3oTuDM+p8m6bhos/8rgvLGYsN020LNTqP11e3PYk5D4cqL9SdP5KrHA2LvxOQjzDe69LxtsGl+4
8yca0dUVPFty2qCXkYLgADruGP+i9+Kh3QTszW5libBX/eGks5YMFgvgBPcOE13tDH935bgSBW5d
gi8qY5FqtNI4l4wsOKl2lc+MRcEU9/xZyM0iab88s8zn97eDEIQ7qAxVmkBixdY2RrhfbLBb6PQM
yML5bOEkCRqVfzup9t9gX2ZeBtCEE2V/jtpNQWKKto9K8layDnvIUHx57od9jmHzPLrrGxOG7iES
AOi5on7ZtIj0HtY8Wt4vcBWFOOXuR3vI64lcK6+SRi0kaItVM+sZGJPiTCqLE961DE6tbRO7BaXC
rW8emh/9gwKhTWHc1m0lqrep5tW57HqOMOnFYgGKwfjrVFI34/KdXIIh76GZQpn4D5JjZtrw84/c
b5IhGAmKkJvUb98ZDIBP2r/B1O5vBou0dLcgbKpuA4ZqQQPwpQx10GLdtLGM5Xi7vgyNtKK0xGVc
JX4UVnSe4S0qO1jTbCMJvZUVaUDTlnbpZepf4Wao2Y8tAC+ZnGOPZYpoFw8GAz1Un1d4lEUQL/Mm
bwivjGBl22ink53Q9fPuvYIUjt4P9B/IzkASbhgMYkI2UoY4or5jD37DtUfkNhC2xxMTwUghtFSf
cKSQl2QUz3g44H+yWfPUS6jufUiZaX0wTPKqZuGfBuNF/GcLgR4uTORyJ+InJ2iLOy1+ui3XEOeu
VkwQDQurEJFq4tvz3qw77lCT1T4vG21ynck+keIH91hElILR9y/EufcPijK7+yszEoWcUVAJdPGh
itjJ/II4141v5Spdknd25O6M0oe0rpgHUdC8J0TuF1GKE9vmYBbr48a5H3yJmY/+2r+EyUFMgn92
VXlu4S+80X6PKuQepnj1siTMmEAUAOq9l6GojGJcVzfmh6ZY07HnA1wfVEL4pyrW19iJcSLfs+kP
JbCEuOv3iQrSHz6iUfDhTtio1e3cBx/3SlmA2IjuPg0eZZoFu0EzzzHokOAFwC7NpwmKMKMVtj5T
7xWXtxgxPRZYENuiNvgsjKamVum+loOSAUGHZAhnn06LpwQy+w+VENudX0ZlfEHKRFAWOUcMEgqr
6vC3DTOXX9EtXdb9CPxC45UW6xo06oBis18GxMIKtWNP0sWnGM4isTOah1HSRYkWd83yNHQwqzRb
9DyB8yMO6HWwTJxB8LLmSVDmZ2Jyexbfql3ZLsexg8lG4Zp9J3ju9HA8Jokvui9usHciUUeCagPp
9M/0M3OPAxWJTVKQjqz3KK2U0pnhZzw3Hbxfwqy8iq78hfLKSVrnHEYhOa+R3rf/xqqM3c3GSHi9
J7RKsJIcv7tV85A3Zc70dWDAb1KViMz7aPp5csXdGWVo+x62ueuI+/UJZydngMJXh6kZ22jT73fO
HvfQZrJiK60ivGc6Ud3T2zBUcFHAEV8BmKtxAwSRZdNYbZ35zj04O/YJqX+Y0PVnCE+6VHoWD1R6
3umbYqx5BwvwB2/plhunwydJIKXbpO0ZobpMfQXpknqivr3xMh0iLd9pfDQO/ohH5u8OT17yNFpH
JEl7bHfGWnr+zOngVhIAikcetm4Xym9lYk1IsEQxEiJtNa/2f8Gu7WkNXypbrN3+541DMpkg0jn8
rRRZi5L2gWIRvJB8zrMrjSdSQ3qQv3rnrLlU8Zzm0FKn61rGvxgh4Ev4BQWFHrBtVwNV7XtCQ6u3
59U2YxCjYQHG9j8UiDi005rjkUBVeYzUxUpjegP4+aSKOyj45PFcI3YomdO9israuUUET9mX+miM
X0JF52u3/S4DVqnRnKqxY9xJZjTSXSDCjYo17xRhWAvcSLY9ehNhRqlLQvkZi8m6c6MoZ8X3319a
iJ5z95wf+MqmogF6NZHALIISKR3ffF7/zB4/Hd5HdE0iYzYoXzZULaYO2d/XvAySaH+k5XO+ZeEu
Avm7n17DnC2c7DczxcjB9/tH6dKYJydVo3DuMMH5HywTt0PqgCl/Gt2bC8/DniXhnvw4rIrqSP3T
NdJkR4e7liiu9kPNHOSiq9dxaQbundK7eyW1+4wCMNMeyc21gOG0KhlPzHfJi6Og/2pOj3qMvbyi
1W1rnMHh05Vb6aG1eiCc19MwCHWGUcdFGNOzfaM54v9G/Fe00DGwECCoDD/o+/9wV/HdlDrCVFAu
PaBCfmryGORRKAxSClHRycV8M7tbgmCTTlNRJaN9FB5SK8rnApqA6mofmo+ko87iPZaY3G32kBOX
5G3cSv7sUMQBy7jlylqz7I+bOfoWK9pvq02OuFmxRODNGWIxZHnkm2L1NOe543yLuVXwVrvDcaHA
lGRw8yxUZ/WVt/2MXkMyX2OAHS8K0OUIRiAk+mS9npbZ//ZR9nqwRdGBgfnBqfIsNOR7zshmZkYw
2shnnVnO6lM9WR1USkXHUlYfeHOy5uDHpNnJPoJI+bnDo2aqNUNodYaSw/3YaoDNLArOy8goVyY/
HHYEjIk4dfAm8Fnci38yg2aZNigboXend2lyx4++wf/NzYWDqLW1NXpBrWzjDjgOWxT1+QnxVHK1
sLt6XAtP+AzTRgbIrdahxpHwJRV9s+WIeR+h3x48elPSDlS1ZSWWSV/L46Evh9efHKGpa7JeYHAp
qGySpPRARYaKuqvFZkXBG3euJaNXpMfxfdjo7rc9hm4HRg+Z0v2JLnnuZ8jb4fiQEmALPWeQTAGB
ybbfGHzjsyB6lm+OStyxz/jDN5WADxCMDWFuJ0TJQLY4rfbozYcC/iiLWG6Z/cmfoGU88zhY9rKy
+kChpz96TsPOk/dvR/X6mQN8SkqQ2r5Hlgqlh9UdbdOGzWfHz/1p81pKoDMQOlhUfmCJPptZwdl7
H6bYoLcXrlLKK13hC5m/ATTgqbdsJuIGh2PPK/f3p/phHdLba+jUodafckY4kChPAkwHHS78kUVR
JBBNRydiRAHjDbohWXr9Nr8hD0jiDUxoKsKRi+OFx33Cqw7xqTmUmZfI+bLa+oiQdt59ZUYcdvN7
QV6niib2BZLCkN17TyOg39cLFtdZNr4Yq0NauI3kZMJ04KZK76VSu2ak9uF+C93ZXrd1+yENHFaj
D3is+poyIUwvGEX2CmqXmBNXzGf2WtnDyfMNIuFAsTuyz8wGE/HwSLM7FsohY4x31XpeGfFj/SQz
IdphhtvNK15NAGcuoPyoyZT2etsd+rj4Osa7aYrhiLbFw7ojcgrmJHmixaznEjeo/tDYqd1L4tpN
wglfbN4ZCzOI0yorffRxQW0Mo/vjO93fN8XrcAgqqstMx6g3gLYVqqI8rlFvoQKI4ff1ERfuKL2V
nXZtjMXUEdxVFnSQtg4P5ixy8kjSG3oPh5TfVkbZe5LHtLaDfbZwbTPCTYXnRA/MAlqXp98g3RvD
IPTMEjlHIBiUlcWnSdq4uWT8YUbVuSzILLq2YKhEyjl49Zcer9i9ilOOt1cwdswSMbVaOB2GxxZa
AigW0jvteb+/gspALL1wF++c1URbtZHumoHbDZHRZ4WPWVan5rk9RmGjciwT9GsSkRuIH/+g8PJq
ujqtwREiWAMeSDLKbOEfPBS41qT6EB8fYj5z9tIck+I0nG22PLFF/74BCcFAh8pfsjm7nJ6ZFsU7
OIXYCPg9j+CbA1L3zz/pXmL3qucmINVPA1jYmOiHx5YytKhH9geuxw4pV10KZRdNZpGz/uXvtGck
3kcpRYKwb/2Qq+oZDTNPdErho1K71IELhJlaLzOGfhkLuDFfeKizD4OSJcm8qn/ye3vtf4Mgfe5n
UchbsSUQmmDpU4/98Dqelkyzek+NlCgQK7D7XEr8QaAkgLWd8Xk3eXNvfAhuLrjZ36RGYvu5b3e1
EusNtVy5O1eUVONiTMzSzvTMlZclFE/4FEnOlwu1i/vIbUjiLA4ryYJEzuDum6uIx/BdVhoGSoeF
TW+kVnSw3PAQafkgFtMjov94aByLbeq9XLZFmkhadfaYSb3dVoteqSp7JzjJAhk3Zsd/E6vQztON
VypZeOkMYJr/qyaHURDWOtefjppRE6COm3h6rDu6D+rdkw7YTM1c0TeJgXFXRoT8IJlvoPJEbsg7
79yyuNx7GdK2C2/8rkwCq6GEgM9Zczyl1b9O+oUuejcETL0mYF+LSU9zJXETB/UvindE7PYZ5KBh
mObK/PkI9HrmDZiuqWZvM+pFcONle98Pm9A2+fdjlM6Qx6MHDhSUMiCAa0qEEkJFTSW95hdQVLai
VbjSXxbqA0kexiCwHDXYRF+0A4Xm6zGciL44f61xXetA9Djj8Jb88N+OfrAXLzSqoqYdkhT+gJRy
t/xmSzY2dzluIFiH4tU+4gbSVUmvIAZjjYjpO1fdfY5qsR0aMUOPioT2cg3ti1L0Ccvz5DT2ghCl
JfSj/a7PThnjuqXE2meAAdWD0tRjmiswkwoqqQ+wDSfBxPhUAi5G8w7wouV8a4M85wEN/YVW2xyY
ZkgigN2zfUV1iqfBuU1VYzjX84OGLh08HIz/QrSAuu/feOEwfhWYxkuQ7Jclu6vIN/9UraQFgdoH
fH6LK1zCdUyJpA7EVMoKx4Y1htTQ5Dp1znE+Px0SRB15pMIE4P7uD4Os3sxBLTLChls/H2RQPxfl
30XGcYit9YUKbIu5I3oXd5oIIM6KXaW7biWYOPsANQUddwaOZXrOf5gwVNETgqLVVUP6JDMY3y0I
e1cnkHhsLifhN5WmiqJVvyp7e6fy7siYZhTU9iS8S6sw5wr1K1sZqB5k06IXUK7De+FpIcSBglyB
Z02NX3yx0eyU/jCdOiMUJiArMh8DFbNTJsJU5vS2IHIowMQZ/u3+XliQaSCDK94/lDMZOrkTPD88
u3RuIIUu8x1uRb7B7A4gD10kAL40JW56i98If7k39Qg3cD5SmkSJa+GxpZmG9Xjl1xUUUUnNTK2T
aIcOClXZZNjbxb+qLmCahH7E1b/QPq6UBC9fnZQJIeSIs9dCtQbSnc1zQ/lWPKg6g9bF/4UIBpr0
OwfqFMY83XUfeWW3MWQbkfHdNi2CEMQEEVvbfpunSlljf0P5UhGx6z9GYYLJaW8VrtQvuIpotkZz
vCQ+3sN4CtxqK8QBC3HVQjAUSh2WMAbJTM4rCa/4CTIVZT8yT5tigGf4VZyvLi+fNydohQ0ekThO
jTq37D6W65UyZOxsARACtA80u5lUgXMA44J86dPUwVrky8uqRy5jRHSoVklR1EydER7g4HYQqTwS
yJoVB01jWzg2wOFy2y/67P+v0NC08hzBYSMfH/ub5dSYsz3GO2Ap5de2qku9Kqzc8OXlDOrdDY2B
+20s0INUo5T5Ro/ibwZ7lftMOvqVbPNsrN6nYQuqGLWWprxX7brwVxJaw55gVrUb/uuDEWeF7/Vw
frMEq/0dc0jhc7eDG+nYGZdXrbq4Dyh4WPt0L//zrYRG3w0LCWQSQGajUzt9Q+OOt9nT1+cyi98f
TH9AlhvRHgV/gvPS2SMAyEwM4Fj74SXFQgHMLc6azv9w3YD/BdUR50U+hCWZyasqsAr3sNYh6Eu6
I4QnlneJnDFYhHZWoYuuPhrQ2KAc7TOoacqxk9N3R7tQ7YJ73PSVzmggwkkCtx0eCt4i3cURy/oq
XqYPt1z1uPHX/NpLgdOwz4M97MVyTJ3MHUVSTZ0eDR2FyDGFeE56HmRQVm6sq0Gm7QEmtqg+gFL1
k/Vbo9Xa3P3E4TKmoMu+p7JUy8iNnxjhdsV5rjhRNDNJZp0G0zi9BQSZKytrLR8S2p32C6fphUWS
FQmlY2ixbwO/BZpyDMSopB2JYn+qZxL20iNX0KFnDYAqylMeYxElPurqsY7nmMJMCnjCHXlWcxJ8
MIP9brEYnaJBjp58ZQswwdnB8OAsmTMLDoC2F5sVcAX+iqy8NgDyxyKReLxjNCtKBNvGrLyMnKAX
9Sxf9fG09OC65rvIdTOm+q6vlUK6h3HtQz+Zu7tr0rNrLxUZUGmBW1uIQUDWBgK/xjWNXIZjp4Iz
kxDge6EiBnhZnAnR5vXM/dK1kzD5wWM2THJ9nNj4do5y+KO1x7/aP+nvwJk3XpUVTj+AlA2JdsZG
l6stKRduCDTmXU/LqyWDxwD4WpVxCMsknrzmwiaV14z9xH46g76XU7MrJho4pDPQBszF39bYddjD
wPZXRS5jcxLcydbuHP+ipUws8kZxP+FvnRFMHxBDLMPYx14+WlpaeIPw7h6BO6vftT5BR80Wpx+z
4PiihQKd+1LifqJDAVVWMIenNdzJKzfXzXNIBzkOeYQTA26O7YUVeFH+0Fg9Yi80czpGIaogaTji
YTO7KvH60n8jXO6ZELh7K0Yt1rPKYksphEtCZEgJSDyK1ntqFgpFkOeTL+G/D6hBKoq/V4TE6krr
+bKoY380kEpXYGLec8rPG+uX3J2f3tlZ6zeqj3Y+pF4Lk8AT6XEr+22Xfi86uPbboAQuevjqC9gA
4/hRyJzZXg0sYNZInUAuKrEjP+3iSQPDj87D8vO0tLNsw/hn8F3AduOvsi7YpaVrpsDk8ODnGVxX
p9hOv4s1+trdVHohubDIKEkK/ZJRHtOWhmAQcGXaiqutQI1IjwdKu1MnXy5m+snMzbW5rDVvsTi4
r5EG0CLEIFcr1ClaCMVVI85p61oHrQ2/3O5YasELwwm7wFPYPYD9yua469z6X5iV8sd8SQg3EQrY
3hj+CUS4JwM7jIln5BVprSRM1Rs4Ifl/9wgh8lkzxYVREzE8mqEJzr84Jf28y7y0exSDLh8sM13z
rZoTrjLEzLhyLrBK44L5EWyes1lKIZ0lCZzYP6WxoS2OzFjUUuSjCE12xaPscyGy2GzVYCPmar39
PFklEGxHKjn4Nd6YHev/YIkBB1udnoHy65MJFqZBQE0ZRIbXFHyJmhGdHV9qnoTM7HNXtmQNaOtB
081Jam8gyuA/7x+mr9HXBCStwf8nPMZp61j3ruLw2fnzltX6uvkRtcDYPgrqK0s75gDwVXq1aGYW
EJN9kfNpq8MWKfw3pRzO7g3iMslSJMp1T6YEuIz4QDoBYh+4U90Y+r00NUu8whkAIJvvAJVUDMIs
2XE1YkXx82h+NL58Pi2uSYldomKIAvF6Nb55uRRW+sC/v7jmulDIaBS+GYDVy8x1zXeILJqVr/YS
PtfwWvBdm1ow6gHATRrC/V2639etg23idQb6jkVF8WrBVJIpOqmRAxtIk7DIcGGBSspt6Zo0fvOB
twwrKBtzSznDa1vJ4+zQ7i1LQQHu5jv5pW0sjiQx2Bk/guZUjyOWB6wlXFR0a1r5nnZ9zs/H3li8
MMliqtLM3BgBnWieW5upZZNsUf5ggOAx0V/1Uga82fFHpb+DTer2O/yv/3ALi77GaOGNTCbK08lR
rgsidAUFiq9tQQYqLHAf9I5oM2J+uudFNwMr9L9R2+++kqDG9c3f4OcfoWtWZ8Ui1NfmdS1ngj+E
QBxddvYQzq310xtFpri3uSAkgaPrJviSREbepIt658Ft8OF5nxaON65AgicL77qn9ZX+CZurEFE4
7IzhJ9AhkFnfp9zNBXfYwzmTq0t/4HqNW4BHvoDkk9d4VTdTeeVxN69NWrvoKJs73LDtkSxRukBW
QFql9STvq8DHrqZVtb4KfA9+NrAOoMk5Y+i10JMiNydpi6V5iCVOK+fCEshziDcpkgzYp9ZjHMam
g3jOQg8NSpqoC1eNb8M8/rs4rnWA30zWQfRIsw+fyy7YFbjO+P6v76RgRFNLGTgaIfj4G3Garn/B
7vcCdMOkh5RznGksxdqCLmMEnoWfSMcZy/V/KQj1W0Xjcuc04KO6Doeneb4/Ka3Ii1M1k+xXogx0
9PEt6eX3e+rfBPs1mwrAMcgpuMx1LvMQtoep9dL6EFWJIFNm7Y4zkFAoVRp2GMm3yD7V2A5pO5tG
ZWYnGrRfXZOIyjEHIrGy+ah+YZjqd+ScqoD9exDN+k7Kz8TIF76g4HitihSyHpT3pFTxCa3LfY0H
DBkTUvPi0ssgUvlpL/zS/iKTTMDzYrOPUkDziqSOpxOsopMqR5130ZWLzSZo8TOqJd+rQ4RlTV8h
vHtpn8/rn+3ldAqCmNgXXQF70iic78k/n0+Bjiu/tn7iJBnpa3MkEGxhl9dEs4/mCyOWahdL5NWd
n32mFdrLtW86osR9V32UVOMbR90rrlzKW48Fll4NxC2ngA6c2BR6ruQ7ym2iU9XNbkyvKV98o7H9
hD7HtkImQodmdhKY+YZHAun2K8Xmddn/rYEo0sJIW3mEEfMdu0pRIBhoEGTu/UnYRplEUxpbQc7T
aYZDB/T6z07YGbDh4PGR8gSsD07wbfXEtmuFL0QjBCR6kfoVj9W4Qx+qVobgUaTrACk2vrU3Ip27
ss9lF1ZMUPABs/GG5EdUvTZCmGeiw2As8yIQ8zE7EQDVF8JYXSYqGhg2clPTw8shpDKUg3C8Tdrt
J8V1B83m7WhSEesWVBDBPDxL05BUjxcnQ2b8E354WGr520EBUJnGVrcuhKqqVr+X7eCj1fy0A1VB
3MuOgqqAAYoO5EQLl05qeo2jsqhUpF1mG0S6HWSSkh1Rxcgu3hM3KIzKMgyEGwtPsFNtq1y2oT9h
yL6DVEDjZlyHDb9u7AeDBh4kb48sALBw4XrkTZ0zcvW5hLRrTyk3EDDrx4KTKQGDl89JkoPsqJJl
shO/J+uQkTzYkvQ5aP2PbPoE2sriWXW55bgYP1jtrGfrGWdaKeS9fbl+1lwcPguomaadFceua22D
8AIukAItyNLFvwZi992p5O858vSqfPjZnoquFq/u7qa+Nc9qZEELe/CsJ80vz/4u46XrbgMPRfE4
LkRQsV99+Mo0Mb/4SeWL2dJ/8mWCKCcgO7qiLowvQkoLRB9itwb1sP6YkhfhSL3Abk/Hy37xYn4O
DM8xgpquYpIlgy0gkYaXKnIXi6G4T+u6QdbzuKuaKgGTf3064rIIc+MUPujueENYBrBqTdIdNRq3
BlkA99zmrDUqubigISFbXr+17X+JyaYkhgXtqLogA3Wt2rmHP05+1htatLBSv3z1Z2mIU2DUTsc5
IwBy/L2DNNyN47xh45DMRqZFF3vNCxBh1XeQZK6UjU8Mt6yDSzYodoWk05eKJCuMQaLKRv43ZMxb
hbGh/kLDnNLKrzZUoyga3ARBEci3cifd7Buqtay75iE8E4QWqf55ce4+j1csxl0h1JbzAI1Z9EBQ
nOEjqet4XWJfqTmgRGEUU5KIRAG3lq45NjOX4VxoXoDMeRMP8JBXpOxHt/0RDfPKJJ1n0jnkMaqw
aXfjo1ZJVvaELZY8koAGIIak/8lbMqbyP6+XMRE4Eu6Vs+kPc9JEQ5xw/e0SEvx1KQX7R0ucrw8g
hjDWgGFyz/Vbsp6Jk+cPQtOUCKJtK1vBOrrfc0W1yEHTVt9QQPRJZWzYqtda0dIIG3D234Eu3SQ1
+u8ZCXe3WnyJpB84hFOpbqwVUTgjbLfHYpxvYRwoLpc65Yon0b4ozigFTD2gGZz3w0II4sKp9Tys
ICOHhqPP7CxhPUPrSjVSe5xUma4JyEUDvrMYxuqjKymzJaHvdC2ZGNjySTeRnnwI0x/LKh/5ZDex
V+CMYKE7pLGloDrtD2K2rOxc7+miDCnIfek+IL28vFLk4phBws72DYJb1z6jpc2ivrTDtijcw527
9Wo3c0CBdju4jdsUfAhQBPPN8yfITD3U+d3COMJ6TsHv20XrCBY9cnvH65v8Z01vpKZP0PB3et12
taxkPupuRst2wERh8YhSWn84Uel/iNp9/5OHvpiEs1wXjJYd0rO7A5CGJOcQLMXj2sJHzx/zwDcL
0BOo1ZaPVgdAyfSeUAlvrsQq4s2OXotAKNLVhrAWTJlJtCDfoWW2kkgVL3cHnfLIQg+/Zo659PiJ
DMnaCXIoOxRZCISwaayx723L+BZJUaoqBsC60HAFdxk2IVF3Vn+mc9OxSUqZ3t9AcYZ4SUfdIQIM
9zDf5LFuNuGx7MkyoIjGVOWjP+a8lQfP3eQ5pQyip89lHj61l9UljTbejrZHGU6ERnuq5Vn75Pyy
I5fFgWx/KQDMqvvtkuKuGSsF9FQlevESbiTUPcJvAg72H6Ix7GWkdYEm9IRzBQswYX2JhGudEXeR
r/C3GKBdaTrq4/UiyELq+gnE+qFSm0OH3swwgXF+n+9D/7njF82Tw25qaPySsrvZ4CC0DruA+G8S
auJc0LT5psEl7c5cqIydjqextrarXu3zIpcpYXwjhInNVB7itiokXpY9+4xJAusDQash8S1U4Vu6
lqcbYcEr9xggwKMqNkQFGc5DYPj8lEfi6B3z5ZiB4wWrX03vHc9af6BQ2bYmepxyVZqRZq8Q+16c
H5898U2vD8vUAe4iu0BGjKJoW+Si7ZyJsEyZbpg7Kg0ZLVxROXEaahdcqJb9+8Mt9YF1z7YVrAKh
FpUYb8knj2Jw3TEwZ3ij5eD8lNVAolfRH++gc0fw6Vfjnpau1ZyE/VZPQx7coJC+xBh90sccrkLe
wPhCK8eNZjd3gw3fnSDlzv/0nIoHri5Pwa7W0cwCkjDan45Adpgg79RksfN3wO4VTonVxPgtd3e1
TUvuWiR6MxpkniumsKStb8wWbKIVwlPb+218jkEdKkKa4jF4EMv1c8Z0WuUb+7cKRQLUgd2WWhrv
H6nKHIV6pL8WefTyjmuCfSukJ0xDzzdOYArX/Kp0TWUfvoEX+mOnPffWY/JfmPuzc0ffSLwgifJm
q/fr4smhiBPggUKTaBNCjaTFtSSgWotl3GziyEPsjqICeErYvM0JyBezWD8B5E33Cx7uJcND1jKD
OP71GJ/ENZbA0BxmVK4RPAjaWDT+/fAkIqj0i9ZLTCVY5jf58OaYO0Pycib7DTnNuSe+tTpRdPox
49L6YMMmzNaCZVIpPLa50xXi6Y3/GhLVRHE17x3dl4um3UD8F8FnDyWgIB82TWcmqLsKfzKB2+Xr
aaECaMHRoHkH/HkGhxRWDDwFSK5LRWWIn3jTVEJt9icgFEWl5IhRFZEw9kjNocnGA3y+sXdrVg4X
PMVO6mQa+3Uqv0w/EZck4B452cMSm58uV8NLzSQ4Yd+BZ6ET/7ehzSGggr6DL49ESlm0jwSq8c9/
oSVqgJoZ/T8lDoZcjDvsloy1iUiI1WBDwhiQsJL/AdMIXbfZO/iRBAkZXly78kOqzU6yVhY24xQg
ML92yycWA0+YMLnqmwBelPPP0OfB97yG0MutzvKLvJyeCBSSdsE8gWQFsrQ0efi6UoH5nUYMDIWN
CF/BVsXiZ3DcO+mAOV3o9BAx4FqulRt6FAAQMNeFze5Z+z1Yz9STfAblJ8nO33KBgCPyIOi2Bejs
h6mpa9agx2LIa1kZlrmpDPK9NCXcUUovEazNGLn7gZboMSuRl5+Ew0I/CW0o5OP8R7PyEP8E215b
BJ9bm/cONHye9qw4kMyg4LAkyAlWgDv8IMrTnRDeqpFMEe7/91BsClX4fmYglOis/s+iMyhzyyBy
2SZxHkNunjO627WSDqvF+yxpoACS8eqaEQDn9gH4kLnom2KZBYDXJI8UKoVpBNToY7C03vUKnrq3
yWl//VslSOsExekuLoUe6Aypkh8Es7z7PDWOY8d5g7f8YlorQsxWQOdBFV4htgXwho+3jGHT9GWQ
i74kj0Jn/JNBRpNwNojsdZgQ10Tn/YxTiKMvex8usWKGBTlYx6EKxQKAK6rG3WyakAu+axnpyWlz
l8YUIyIoUUb4jH6H5KcSx5Mr5PZxyWHunkRgvd5+75ctVfiM6/lSCNsVIXYUSkegph+UU2EKiAG1
+lpsymZ3JonIEn8ZYTkArVVr1WvjU41elPB9yg/Uy+4rC9J74Fkmk/gNlbe5IB5/rwxIk2O5vmvZ
sAurPUFm3v+Wha3XNYbQ/V6530c3IuafxKk931beJUuygA9I1vWueoIKymyCe/2hpaGVS+6NwzMM
9uf0kLmc2ADrTHKByBLlewWmPQT/2ApAzVITLRAKdtdaT4lKg15q2doVxA1r1tbRDXzIeAymwwEM
GK5Y45OnroFjyW0ms1sr2IsnVSgzj5/AuqpW8vEMouRvkNtQt6JgQXxCiWjafY3fkDbkGpn9p26F
D7V1tnl79ll6zalgWunXdFpHN6JPry3i6dz2pKFeFQZwv3mCoDqHLwUI3OQj+dS9IV6alarBRUL5
+n1d3a8Z8QuC0uI3JAwC6mwNApBZKKaFtYi4Zh44PmEEoxIh4l5tsjWZRpAITcr52wTXW/7nDS0p
FZgFhXoX77qacwkQvqhFbEpbmCgjBw5AIlDPS/11EhxwmKk8vfi4989r77lI2qIZZPDayWOGQ/SR
P32UPdWC1wE+sP56IN/s+8CAiRbqzy0jMD3eVTft1Ay7AcZqJZRpoqIOh+EGXXc9IzKkKi+ZJcW4
ffXc6gNtEasd+ozQmN57HFPaePeonAwtQNl2xYRo2BWMvmeazFrX6qIMhx3uPd6srIz+fM+Lj42W
a7cVUbBI6wO8b9YcBndZXHVtdal2MzBkiipqjAtFNPX96IIsO0dXY1kLs/9jthgV73NBjJIVODX4
KWqGz6KS76ajuE1JSDkh19BUvIJPZQMUAeCvED2t6o7HM/QUIod/6D6FavlSqXDNapw756RftYgD
rXOkcUckwHshHBusp5cCHhKhAkla0fTHiDHBHrnlqqKFYMHXS8sPd3QfiKX81RRT3qUpfEmVpLLS
rZ+KLaJYoBd5vxf9m97UKJE/JHVBr6fCJAdS7SuA1Q8LEA6n9HJ8WcSMiJ17iFS5QlOgSpJnQF2L
AJLK68lgLh4DYkZiSl7fc5M2P40KEEER4EVVN2Mv+39SqbCY2k4Ia78efFh8HkvtOK1lomrJaXJ0
yr5QomoLlwZKeNik4pHkhKV+kvgZw9x067HpH9h5CNdT7A4qNYK7AS/xiJ/bBm5u3SNEZ+hj86XQ
Ss9pOqDE6tFzSn+Px9g4WS6yslCec3H8L6xz6LobgRViVsQdwSvtQ3k8d6y+qUGi9wA8sHMcPVMp
FRqATZGamTmzQ2oykv5KM6pXa+qTiSwkY9Lvha2fL0g5E/nXe3zU/V223lqV6mbxn9evwDM4m4Kf
scxf6LdITri98w7lJogIVXs5L6+q3gew4X377D9+KeIlt6QTxw4R1PUxUqBEHQBwhg9gS5NbgP18
bS6+KvbDshQsIZ19VM+QciMsWMwiRvcYEjH9846MEFFD59UvjE66j/JYDGX2WaVSWV3kh/ZKQBSZ
1C11+ffHizuYGmpNGXsfBsRk+5JGuFeAoERa5RstFnznksfO9cQ5eUoq1okQXosyMccyW7xx0VOJ
vdqNAG+rwT1zRcCDU4s5FWteHR9xm/a6qXuCpuYVFuVio33xAi8Xf8pYpWrDUEfaVklyVdm4me4c
kibYfEOW5hjKcUmSloNF91hXmTBRQvoI0OjOwLzCT/YYs6VxqDAIiJ6cFfMLUCbiheb6acta3Pib
D4OxceTMAx2gcWDT3yaf/lXTDktv1BN/KZCZr/8+2/pPNujFQ2eh2+okewaBgj+r8O0Z7THXtMlO
hkNn2fQ522FYh+nYmsKNMMusT6aHBEnfGRVhvJJo4Q5+wNBKEK7XY5nhYf1rpfZav+VdDBPj6/JL
8yabu7sE/KRMlE4y99F9ir22vTxx2Rb4eN7/VLQY5jRkeHyf5iGtoO51wK6RXAELtE5bjQAc1qH6
uEV5tZGiTw4wzFo4HJeG8ZyJ4nSTQlLLkYU67PaA3gHs6djIHLwnfupl2MQjUS5Yux4sn/fVeLOo
QrJVTVhPa6wW10O2NBrRdaXrJQ5EC0SVAXRX1TdrKxmrDssXhu9oNCZbY3omPcEyDpm8tq+iMtr2
M7X0iwZk9oq90J4sl2GAk61PPx1fGWWw0Afjhk6NlW3unGFimsuYTdWFrBGep5diuY4JqFEcrpg4
UoRo557DnN0ZhWbM99c2PHOFFQc4CvmKgOcLtE9BBmDmBucwwjYwkCVGuNpzKGRDUikjroHJfy0D
K9axfXa8wSy6lX4YVbB9jxUMju7LEOdYq+5tQx/F0RefjYBSQc5wf/zOa37LWAu93ETsSuWnpXRF
e6QQ6d32tvRE+SVUaRn2mdfmkp+dxi0m9biF4UR9ilaSsR1K9RpuQUva1ApH/JTOo7496x6Xeg04
3XKEDou8PegjWvxY2C1KwGxvzZ2JLPWyt5N18SZAjgkH4kRqgVayOQiFvH9iJ0ysMlfGn5uwiUTq
cx3pI/k1OI9bP2ZjBqFH7oDvw2ecXdPuBGuwOnS5rCNtgLdYz5dDp2fHxh70C0XLgn1TXWRKepFc
9Pu3mX9CS1VyJHZ9SiJ3qmBWYkOderLkcjWmTIXlg88Zqn+bI+J1tekFhcfqk01LDw1xdvvdR5Ez
ZgB3jeorGJxn4/3sJZRHsDOyBD21vPrzCcTXKYHlpDBZCGuMECoZeaX9UmTqqzAJ5EOG6YWq4rf4
vjgPluQl1BKkfe43Buc8J/wXE42KE9yxVXA7OlBoq7MYId4a8T3/QZSD2Kpm0AQ+4GhlGaFvBCho
arBxyrWb23WAYwuvBN8brj/o8ifCiqZ+P+iSb6SRsO0yG9QaK8ReWeivRMlm7LIld9H6fPJGKBcK
KuJNnq7E/zuK8+d015I8vpn5+5oXfO7jQb1UsUgBRi4A0R/zSBKx/fqEBEUSxYn9R6Tqxknz8RGh
sGX6IVZvn9gL5feB0FNoXuBYxHkb8o7XhODmsixX4/jkLdgzpJKsYFQXZ00OUBWgosleHrJNG3bd
wWCQU/VdJdCgZnIkH/tdU8If0RZrHhuUGfMTpqNOmSGJnMh6eQTm88vLR9kkywoIHKSu0MKcjzWx
pL8KnTVFjn3TS66gDaD2xLsUcP97nddtBiHbaCzHoyW0EPY/YbfozSM/AmtmjnfCI50XO9SbaYTf
bt0hzFB77YMViTPzrD2+ubB+cozZ1X/JpSYtq3KOKX/VsIxPrmxu+UioXJwbuOiCC1zJulY6R/M1
p77mE4MjJqy/rpY2rl5nyokKLF3ra/XHxw7q599gXuY+k1jR5QwgMmVkRAhqviEeFsIg32ULjBRh
xVzpjKEVm0Z9EoV7O7A614lKYMts89B6Y+mhiRY73X71cKnpBUy6tI4f7CNGkFhGZFamEP6KWADr
aCH0xBUhaVWNQFpFPpc1em8GlHs/ieE0u4iDJrhed7P/PugBaNVzIhpRWzeyJPGwPXRpaqpPVB6M
mNJhXMqH20KDxxu19ur+iHAR0X3fmMwTdeQOgmWACXpbUiDw9V60ZIbTac11YozvdilIsFZ6+ZJe
ljUr2yvyQEHmmVUOoW3sG+7v4EPNqr6TGRhAT6HO35T90UESi5VClwj1lQqcOjONg4CaZ8akiBFn
ku2fJyEtYVKbVK3fiLpQBO1CbY+Oqwtk/EFTeLoW/9v//45npAyYBAwBmCBoauiuL9sqFVNfwX6r
LXbRaaGJAB+EgxJL/3ut1ToL2IBblr/SKoJEAxCvTJOwwpIiCMcJB8dyBhbRvT9CbftBohl9MOKF
SO1g8EkGTlkpBb15FWgulq8J8BO9SUXRQDIXfR4nmFpyuNnb1OSoadDJQgspO6Ipqmk6eQ9Llq8D
i2m0njcIjqtKEZoTlSDR9jugUeiw1/YmyGZirbdw+uvG3ylrx8nmtTIg1K350C8F2hwdMzSx2HWR
8MCT7P7HgYjo+XQjVOSpgUsSC0rWHui83ESuAwKOlv7Jh2iDdEX9IhyA7g11CnNc+IpwwPw6xkGL
FiTWDbvG9aC8wjfvMZJNXfiXvAsoILdW6uTRKVU8+UpiUJzp0eqNLgG2c/I9n5vZL/Y8Mqwx8vjw
KZQAxw2enzw12NV+M0n1uaNooaaSjb84zgcEtzC18yAxbQT4bsx9ZbjRAzTWCsGry7RAJzkQy/dT
knJXjrzOSgraj2zsIgzREuaQ5kbd54g9UVRwK3lSA7ZEAm0Ta/uMou0iRtCf/aug6tzUx1aj+Y6h
O6XILC6n2qyIehN30d25EIcqkVj2wVfwOAAaB9psGFIVp13cIdlWbHbZQV3iX/VH4QVj9QiPQcVm
Ebl5u5Ho5myeKkAXxBJ6NndYhed6+idJZmTzWpV5HCgwEiDrEuStBe8U7L0xU0u8m+l1uypYZuXO
C4/Np2KokfRVIi4Y7V+xBIwpBAYW1Np54/+wbu/N0YLaHcd3J8zj38JYxqxnB0DngCXrWFlHkelG
O9k2v5dBrthjIRyYbup0qc4eIKHKHzrJYihJrdQ8Xw8ujtCeM6TsLzkro5wttR6SGoTrDUHtd02/
RmaQ+PsAke74PMrci/viKiz9nx5/GKM1pzn2430jHJc2qdS1hOYjG2y7ewa0HN4fHfJXmOQmUGMA
TO5aNAaY1Hx6E/xVSacspls/ZYXGolXEhL2bA1IaGErzNriji3wYa36k4z+nWD/N7C6y63rxDx3Q
jWZFxUKHNrREFrhxuTNH91WoOk9DaObwvziEQ5+w5drQ3TzwfCXF3gr1mni05F5AJEyG357Ja5IG
NDAklh3+N8UMgLNldanffUkHVYOgNKJiK2I60YFeU0bX1QeQwQqH6xfSH7vuD2CUmsjTFSor833v
CmhrvqGN5S/tYp61nlsUt4KEtRB3HPjG+LaEd1UUCZRr8oufi8Rznl1x7iEU0hJ/UvuKLKvefAnU
ZM90VYpjZNjAOu2ZhY33PYf130+L/5/0YynyqAZTRW/ojHJUBhonzfiGhaQfiVgTSLtRcprNWE4U
WAyYJ3fDtQuvqKg/ImH/DMMQgOG6B7GwdI4U5xQdSSCScaR+ODEVEIqYVeCcGMjSmW/kuI3VfT/3
blUF4FsbOmu8Eu1+JwkpblK2MZ/KYjTFz1SBbjO6wBrUCpr8tgIS0GeLtoWb1fs4701oQ/LsZaPi
0y7Txwow/9LwQrJobJ7rb5eJvGiaqDAdQVZWB90Agr4itgnK5wV5Xoar281hiAnQ89ktI2iP8x0F
NXNOm5eWX7QtY5EeXsFSLMoSA8FaCNuvMzNlMEj/goXD9r2325KN+u/hu9FK6Hgr42ioKo69T6XZ
ux9eTAerNGoEQKbJNkzR2qTLXQglvc0Sf9229gVN4M46aZv/ZCPDTLZhZ9CjNRDBVPdHek5RDzAC
tRpbxthFsAQyWAFsTGkJLv5zE70DG0/kIlsxAH5PRYjadUeWylXxVCtcCmxtSYpT/GEzYaFOqoO2
Ww4m4SrbKKzJH0msbVysbayylMlbMdrQtNPTyLRvHw8+MSvLPBgb5ZckSHGP71KiHCAXuNfGhA7p
WIhQe+506BJMs5l4f0CRzVoBKIjb4s4IggkgvcqVvi8vu/wGBdsMez13DGghOLXUkVtfFB7vPsx+
8e9AfJuotgcu0SjZGgMWsCL3YJYJOHe7X4ZX6wAav/WHKUisvxSmXMy4UNgcW32qmmkgUX+o2nkv
NcZu8szzc3FXLo+45xNtYSmi3pr3d+VSmoQ41eMie6z62Giaaiy8fbeB8ci5u3sAZ6js+2IN+f3u
X9kHqKbarf6QoLl1br3ZkMcf7zC9p/TYJVnE4zIdET/E0ABqnoWoWP1A0872PPv5ujdaNuC+A57H
h0/Aro5xEGp/InQ0oCctUQZEBc2eLMtgTNL2m+gk4Hfn5uZXAqvynu8KkTbjsJ9VX+O1NoDcjPvC
GwMTHbuJ6WqzE/89QQ/C+nme8yG42l4qcfRjulUghSUJyOF59G7EgbjyODggB+Tyyky/k4mAqrTk
BzfardY3xw1qZqnPllS4GpitveZ9WGsqBB5OfPg7L/xEQjsF+iPNOpMM/HxXMKAC7A977+bvjJz1
lAb8vDxANobib17pzd7+woWwSNCG8RIlePvs12R70Rz8TMJ8ukWtdF6jnHvnL1S+FlQl2BB37gDi
gDhLczo8r++u+5KlnCmuVVw7O9h2F7zFslSmDrfMShXmqBqRJzBTF5BwYwazF5sT3qmXjjUJM7YR
X7JUDkPkkD3v4guDp8TpXhyofkwbyT6bOmk8WOwP3FR7KMUyYDy8vlhvGkFnznqPKaBVvLaC+E2u
XCbUUqXGO+iPRCTdLwlwMCLVN5U4SJDWFZbb9FleoY2OE7nCKBoQNEDGhqeG2CJvSBq4sSzcPAry
qavMsLYDDfeySCeIUYurpBgszE6T4IXq9rf1DhzfTYAxv9bsoQnjqmM3fqdQg7KjLyQrf8PVdUdv
HxMkax05ILW5IVljLZfV2nuIzldWED6rbwwCzYTqolDGI8cN3Jhdz7NhgSMNPeMgCBq76vC7My83
epohfbIpyDMHDfsNX9kiVZeDIihjBYziV+kk7Fn45MeV/ekVf4hXcRJMC8yaOFaQ5F/Hr/Jz77LK
HtWZEvvt6V8YsWAPLAtT8x/dDZ2AtIUGTGPxVrd4NzT9slLDJ0YlBbZTFD2QzHlL0ermTUCsBiR7
A454V9WUDi4Q2t60NNPxC4TyUfQ9bM3caA+QV1YEeJrObnotzRrGq+QS8K01rv8zcp2Cxw/susUb
DjnPdQfynajw0R02X0wFkKrypT0FtSzEi6MMj5LQ2Hse5ETmbVeWMBSBLxyUSSzyqRyk2BL29AzV
+lKxvLfANk8w5QlDHgnYxmjP5IlLdemJZP/nZr9jrR02TZPbup6bHnBSL7xJrF0okmlnGEukEQi+
DDZT/p0pJOoZU7SP5jY/U9OvCnun6BPf4CoZHkQU1FGV+dDR40yGfpX5S/P80WfBZeEcj8P/5l1b
UsPKvx7cO7r3zhpo/df+3+Icu1Md51VJem3KP8KR1k7rQMC+7rKUDLX7uJ31h/j9HPFzm8Gfj7Kf
q9tldRYqTH0MhPGC1OW50Mytq6a0pGVuU0mQTKe80ufcVgmZ6HqVEJai7ViOsiSDXsEiXo0j/zKa
y8drSZrBKF02tzY78Wui+pQiBf/liF0iEsg/IUZSGWzS8OcI5fmz3y4Zd2I0jxhYRj/BC3hOMZ5C
TVdR3ewc5Agmg8oKscw+6sVRwgCS4U+dHntfMfbUmWTnt5gfdu9R8XrzBiEmAH/fbkhkWd+D9lyF
f+jNQX2jz9HQCJL72MGjJp0xankb65gR4KH9f9R1goy57RMvzGRJSCh+AMszpR2DoFsGmUo0lv0g
tU/jKd41QLShUwegWu6QV4+FT884HQL28yOTgJ0QpAYgIvpIZmMEy/nOjJS8mS9qh14TJpMTWfAn
9L9+/K7Ru6zoh3lLmY0t7kDvfxW0f6AGpyAm87+HzkK1OUV/YLi3Vdz6oPpojYFQhDVPhwtV+4V0
kxF7yLB9oEV2Hw5xX8ILgknK+0ylRSDpTSy4WpSUSPgVmltretEkgG0vy0Oj0akKGS2uXG9n+0rF
5QTRYRJdTMoBjAk1txwV4zfZDVrz+VWhkDu1GmqknBzY2ytCN30xO7O+0L6Cv5ipxBNsSPx86K6k
AsiD4vJrSe2LQQt4Y7ObkllMLhjZa83Zk8D8WgF5wXoKNM7WzetMBGLnDMVed96ymGacnPNOBSvZ
gQD/XV4cpSdIVdBXne5ckmcN25Va148xnDg/SmjWWOhMJ46gUHTiKDb+OOe8YP+ZqJqChwY20p8J
iPzObm8cTr1s9Ys7If56ujbHRS4u7JO1Einiszfs3111qgMqbBss06D00AqBg3sj9V2pSJMyyBob
2iK5ecoTA7tavecYKr1ZzgZJ2EncUiI/rNQITIVyi4AkSSQ+YuJy3Hlu3bDQ6W/8+7PPgSRsScr8
8Vmivb4sR0hdE96jUWNttO4PPjPNqiZmcOLt6z6T6NSacxAL+IOdXk444XMpmd3RKWulH9yYUof9
HSynCgPfbttG+zwahVYDE32+OfRqgHkbEq1ZsNd9T5k4ErTPli7TpNCZjiYjieHra4pwyiDwP4zz
/LtOfdFtpz+nFTfHIPgD0R/MnRcamoiUL9GRPnRr86Ex4U3SZq7YLyvpmtLU4hVlSsvTFECQzD68
1ZDtxSthACJm4m27oYpQhVeSFN49zkt+H7LMzPXUp/5XtHaJ9KTqwCuEn03vJHXhKlRT+i2iXR87
Zh5Aym7krjdnMQiXT+x983C8MngKRoVDAECkF0am7s5I5O/9L3UD2zfDhqGWpeIV+2frAjpUJnRf
mI0ohXwDTNKWP25Est64SlOgARUfuIfsWtIoKkUZ+rFuAYlfqKBJN5oMo6Yy7aoJAcii/i4HNsOu
gyQL2/66R2eFoqMzUL1pQOd6kNA8l1gwq1mALvBIlgL3LfqfrYFdqAhjkegAjVaZMuQ/uot5cWyg
vETlgjZaE70cALSfYz+4qIhuwU6CNMJpzNvXHH7MMq9vUeymIyQTrKSSQqLXGluCaqg7BgZVOcXa
8OJbed+3KVvIe4hUq1hDu8Ep2rHSRrONznAqDqxvj1hfxCuOLxktlFHGaQs6vDNvh0J8Iii7D5Uc
Y3MrpsZKNaX0VI10N+lHIY5qpZZ2OcuL/CHQyQhTXf5R8Z5gT5oUN2lxI3U5ZANZsfEuXfoLEAtY
3F+r0gjtyn1XeZRXlMNDo5m9G78Ot0OdGZHlMB2mSP+dLSh0IfUUq/h7YcMVCEh9p1FwZ/61Af9Y
kdwkU+B13NjUO3izxSb06m+FjKJfSsEkj1aKuRd8TWWrhxZa6ldRs5uvlxjepbuRkPOMkTukeFz8
v4FaEoaM0ajp2NETDXN25bg6oLLL94lh9Ij2kmM1CIPbodsLE5ddT3bUJqW6g5JacoE/tojtN6bE
Kwr3RrBFH3ZDToz4yv578nD0iyr3mJ7g0k3Vl1GQvyhJ9AMFi+72JBG/KzZ8CVpybIXFIKS8i8BP
B1BAVkxp/2rihZU8lzQd9nzO4qYw1UxXQWBcxiAA5xqJjb/s5tbdv1UtzmiqZMhQ7qEGpYV9IUwJ
KMKHtVMmZbho3qMqLTd0Pp+shWn6AmTQ0Kii+exS6ZSwYaD5/S7n3jB5BCzT/469Z1FaPex67XsL
B3RBPdNRkrsM3kaRHOb4jMPiN+HZ3U7WDOgjDqzdNYK6jJIZc0xHeo1Biejr1f9BWB0A3wFFtoMW
WTqLO5rz7sqXZmLKFvgt4hYQ3+Vehwo+RNlLHLry0gz7/246EpgWi2Veeqf2rLynC93Lb19XGIrc
zjKn06xqGnvsk3vZlabJe8pcaBP8LFMCBA4lN5ZEe/vymmKVrmNyVcmtwGHQ1DScIzoxRMoNPyAh
5rmA2O5zkVjVEym0fiEL/Hm9F6kS7tbI0jsLtN5TMmE5HIpmsvdjNYhJGl4khqoKfMCwcOBoJ8Kh
VOTpWVU4lgmP8cJVDgSUmz08F5vmhW095TnKIzigvHbM0aiv7TObCXcVkgpWBLCd2gIN5mkBpt/4
3VgyeEtMtweRW337lWG3DiOh2iPxrTFswqOeJiIElc9PqVrijWg72nBrItFIRcpvYnK6ENTrEC+w
NyBGoJ+aEV7VcEkdG4BxQ4arZCDKlSTzc70ULGFWr6Pdo7McwMe6eD7go3uUVPxqtNMzlJYGpMA0
2kbz9SgvwuIM/H9bL+UNhUnQceifHhTV99GRyv4lvFkpSgPFD732X0HHHrq3LZMooA4shGugA6NH
KNkza7w3ejbg90OmhjeXEIdKf5A5GvkM1AY91plH00aF463T5CdTGqkwNP4ogb8EoPb3XxTS7DPo
1Xkuz6tLpeSwuv8XgssBunVZi21klcjwJVfF/i0MifEh8G7+DYIF/LzKOYGSAM4j6ReAHjSzjE/L
ee13e6kQ3cTBYoMyK5KUrdMWJqqwJPsZ/RYXJysuHkYfiFwDK04odhx9tFxs5p0hU9BGSVKxX9kc
JHS+S5CV6y85d93lyIwv2o9up+UNKJ1NFk08TtvZsEbzUmsyIqoFmWDnLqTuQuZggtwG1ss8SapQ
WWt/StY/aXGvKkRrsaeZ1rigFxb8DIXtv9ZsjAd3x40d3mV52gsBvnuQD87fBrxOd38+VJy7EUjV
p2SX+CXuAwvH8J2LHcZs7fLO5V3kA75WMEVl26LJ+IRdhnxxF6cZlnyGpP9EjXW6oKpqBILmZg4R
VIUkLsDC1riwwKx6yaX4qqhWr5bYA85PLD/cUjMnimhwhcFYWdwmZBhiwMwNpy2OiQAdZUo+apLU
telD5kf/RAtlEIggOkPr86msFdsYTXDQAsccdMOJBHqb7k2zSll42aXJ13ejQcjOlCf21nmh6Xwi
f6nFWJHCSamVMRRol83Ssxd7RaJFjHwrOharOhf6ae2+TN5/eCVLabB6R6l6p1sQZsiIa0YVEHnI
YcSb5pTQoZFXKd9dpsMSLme7K0AaI6AT71tRFwb6XC07Z2LdE07WAWfAfNBj8J/EWCPirTjXAOFw
Ai3AeDZiw3FTtP+SlNh+tSM2aGdnhJc38Zk7Y6bx/TlTCQQeq6Uy7PI4s2cnwTp1oY4VhuZEmfJD
YyPDLWWhV5hVjhEmwHq2N3FIzFE6dW6z+S8y+6rmxwKuNxYvbLb2aUWenCIgsMte60ZxMx+09plx
xTiCidVeVN68q220mBB9Q5YS7EZWVHoKc+1jLNIkfmlVy9HXodTiAtW1vCRVKOWENKP1l/IJeP7u
7mMf6eBzrma32MCKPCS78Gt02dCgasrODSgrKmH9zLnmXYdsc7Z6kXCPdmLpPVSXZxvCpQch9S6H
dyUEgufGgfeDJ5Mb56mJXh+9IbaT3HI0G8G8iSk8KzTUCRqkc5KbB/F0JaTeO94GgYSNsBAIW3O2
EDIPZLjwEnKZbKkxgydMQ1DAyPMyiGL7xgvnJglzuaVuY1mWxr0FgApHV7CgpiXXzLhnLkAnsjsc
pBMI+pQkU3XQAWPtHG8tJRlD7ByMAdEQOsR8Y09GcDsaUJXHQ1Lx+byqfnkJUU9u6eUWvXWjPQgQ
K8CAzY/tLF9yv6xAGrRPOTrogcQQtWOMlUz5E4bAE4BmIdfcf5Px3Fx3pIUtR36NIVelJhOr6hgU
TSaeYokQ2sraaXr08+jhfM55dZnDMcL3KLec9sKHKYEy5LWBetbc1K9j06HcUxVpnBiz2T0GcqtI
VtRogR4WrGqvxuZRiKtXbl0jxmO+kHbHc0kjtqClUDn1g29XesOK1Rns1UwJXVs1N7rQUp5JPK4t
EQlPEbOaJbxT9qHHnzTLboF+92Z3MxPFi/dwPFZPe8AOBex3m49OAqtpbEXOT9wFuBnJNW/34hPR
oVJdVu6MWzScjYrGEUQjYmW4M9jUq6nj7o8469prGjFj8uEYLy1pyN/BXvxNKMezesSoPlf1WBLq
jlMk9FnB2euMnlg0V1goWEHOabtmos76KouEUFVjUSQCqaqc4Jk7fqZ1TDOUHKXqfdxTq8ZGMYR4
UzhSXzYuWNkRMqag3NleGhvN4fX0PV3RXf3R5P322/cpuOM/ywIRl8gZc0EjktRTgMjqtb3q1xTu
Lv7Spd1fI/A7b1Jq1DVcWqcrWMas/Zvq99qRWQI/AvJTv6eio/Qg3nNe6qRlhjA3+ax7uPF9MiT4
8FASW1DnrWvr815R2OrySsQ81eMzy2epfTWpasgBJVSD138CKzyCg0K2+yeki1SWN81bvFiAz/Ve
XkD1xdG18duilUQycf7Ee6j+cBjRbqN1f1EFh8f6NVLoRxndJvTQq9xBEBqKX0mwEbn0aJHlF/fS
yvGJgAZz4bkjFI95EGBGo7j8xNqzOOIU6vQQSmTzukeMQIklqPA1gemfapUO6pWXJ6+M494nyE5a
g3qD1oaHZciVB1nZcxjGbeuT1m+7xjZB2K3R4Ptq+cJ/V8JLxBW0AeZYS6u8ShbGIJLzD0HrtzCb
EIQXcDsiFDq0xkuveZDciNQQ/DPSAADgHUBEPjCoAS0PUCnSfv6WMEz1VZBA7LZomN4KTnQ1Dl6I
3dL3uPo4YbumVoXn8VOE+WX8mLZgPf6iBks4Xr0S1miFQQMTcylSCtxUTbU2tQugtkoWzKuSdwfc
Al0xRoZZmNVPOKHSYl3pVwHaLS7aGklCJbQfq/BrmDMqmN7zp2Q7LzKDbzAUd/BvOGfVltaXoTYY
ATQ2Iu4n5DgWIZRBSk9CMARsCGmHLfDzM3+d4qV2p7c1hU5iNEWfGRP5hR8Pw/qnjXXSwxv854LW
/lhMaCEKQn6mvNQNmhNpCp/1ppWzkVtcMvX4JZmST51WugXRcI0FcJFsAlOF7/okaYHgq70n/phi
+fE3UCafAmuzAR8UfUTv5M65r+MspgxwS2Kz6Vc7baFVr+eROdgF8mGTUdxcXwfZi82htNIXB/pH
BQZZM4RTgM6Qz5CFuZjSUR4tJaK1TiI4vCkhXl0A4CQ9G7A53Hx7XpHIhDHmb0KcGppcAJHyvP0B
aU+FvpqXgHpspGDkyLVxA4CoVjszzPB9mIwCGlvvGa6AUP8D6NQcE2OXiz6WLpBmAc632k0EkplA
iT5Gui7gbn2DHmKxRsJMlVoMDjhcqclVV9DYecMZDYHwxPiRundLfPxgV0fZx/70BVmTxEADBEB5
ABoAqtCPb/k20G6SmxnIZx0wE+asUoKSbCl7ppWtb/ovgdfb4IabGJr1qd2ceRnf2BJOUdVIFhbC
v1P31OaId/JR0JCxrFcEgEWPWEa2SWGFex1gbXfkSZg+jqNxAByG8gJR+svFOw/fH7fTuXttSqpx
hMq2HkTSPH/FbbtUdoLtpFtqTya4u7aidd+ckiCj6UkrKSRLSZ20pEG/BHa3bFc0GD7V+/mmZXEc
vhwzbw373qtrMvG/9rbcLuh7jCio3nebEtgP0hQDtByHqBgj+hiZfFbrkC6gpRMGf+HhJiCnPJv6
wCwlA+l1EQY1t7g7J7C1mGOk3GJ8SJ9NwmyeQ6xZE4SYz6tsUvKWJZxbLNyuxZwayklj5j+T0Jxv
NPBdxGEjM5ysrSA8UNb/C4ATgWgmVMTgmolmgKgl0sNwdVeO3zQ9Ee5RIEMmY9m8+1RiL9Hrlwcs
enZvWPQcO6wIQXEZBpfG17EPNF+nD4UTJ06TeZZrOAHXzO6hYWYXwkHSRdVKx47QmoQis2nwTumf
msAu52ZmLUpViknx0quXG4eEIXa9rInzOJ5X3tBpXm/AjzbP28EjCqZfyci7WzkTe2xizGSu3Sg0
WPu78DhfS/DO1ZyZTiooXqDX0I78jWrkLHVGAH7q1YIaNrqxhUYudwNVuh051E3HZO1bDEPvfQm1
YxsmwQVVONlIxtwQXva3UpULa3OPiA8fpBdeuM8hss+XBk26xm1kelie9ryIyKT8yPXQpcFROFZf
SY+GkCM0rq8ICzzIYKyPUb6buIsh8HFF7a/0HZ6NjG1MCOIDQqnchukTg/Urh6yG5nvK1ix9JKmL
Nj1iIrBQM4bHzZOVNl59jS7IbANCz3zycJMOs9WsOWB0xt9QJ/2N7UBTvwZ0PGrr9/Ln447dUPBR
CgvCvTxCINaofC60eyWzoIzjqP+d5GsuzT8VIMDgGJ3py1cehZHay6cU/Z1tsz4xPzkeDB/MaVjO
8T6oC50Ux8QqHtf63ITdvb0YTp+R8F9tYIdYs74cDL7jJ972UmAwzUCjomEkWSnjRhJoI+0t2hv3
6CKmBEzJc4w06n31iSv8GXEiMxqcbjJX8STSzOZZM+Tuah0NYTSstRNSTFLFIG1I5zZgaVJohG42
oRnV1jPAJF5I5fBGXcl+5hA/9J8+82pp+rAOxfRDv9f5TzvYuWf1jM/cv0vt7vdqkJeiqtowlDxO
gX2zelXkMBb3eKYUl2ZjjvNfC6gm/wskiTstW8/nlVNG2JeTPmvju8/Mwd18Go9StLAw2J2q0RH4
hBn4/1fzr+pXZF+TdAsxA46W/ueLazTcnMKE1/kH6rv8q++RTNOEhaqtxJ4iH4qbzvwwg0npUm7y
KlIqdPfJ85pdQk399XFzB1GNSq6gdHswafNsxxMtgRlFqgtO2yXheCXtxijspseH0LZ7iNJ9SjBJ
kpWfTKJ7KQU1+sjdNxvGb69f0HfPSAuMecorTEGIZdAGiELXgRpTbwvsf3JK5CFKcx2gPuzOWPMO
/OZH5YMG0pJGA7mfXEZILsZSCEtnN6Cex78pec73O3LGkIOkrf6kL3IIbJUTKycwrp2i9NXy+Hda
0eGJbti6P9lopCPnQGCAZS42fP8ODhjIBILDPZPQkXtfTGKswrTW5bnfaZ+PPZUMMLVDxP77lSB3
fvKtScuYNKuFrEYU+EpuZQfIeyfOXjT7TccJp5Y1yFQvqMkfrBEe7sIWMyeaGZ+ic23tx3wRCd1X
+s1kvfIzLLNtqXSlCXKY/Nix6kxmVcGtWAFcetlcZ1iKTrGGZ3gIbceNahou6ZdxmSaY2Ji8hgTv
SiX7s39pL002uHezet5N8FdWS70WF4kA+uE8T2BV68E1UMg7mMeVYLRYQNRFO1MbxBW9L4WGv3mw
64joa6Oz+tJjlRNw/VuHtg97RXsDQMnXQDXbdNKQ9ibuDpYeC17xzyw/2EyY5Kn1gTF8q8an09ZN
GEVCkAdks9UFPz49tY7U5DRP1QIIPhCZu1uakA//rCXPBS/L4hcLplm4MS63dPl9sdtB5lPWIjJw
vm49BnwXKhvfNtCOpuQGH62o0YaRxrrEIBOoed5nLDvuc+pYBP6yWw4B9bDF3evT6MfXscz0ZHDO
/cnPZ2WhAbrY4dym4kOyNqyb9vMIax9G4nr9/8gKc30AHjcrzp+0+IpgjRfqIJSRtkXDrXO5UyPb
Pjh4YBnfF8uwL/dmAer/OTzzRt7B+qoEHSN2Blt0jpvAaRFVIjZDeE2XLcxJLYtwlV/uJl+rmd58
68XV1B4HbW1xCHnvGpnPAWvfQ/uq0Hb9f+5n4JiMrmkDasux+UM2vEKSf+PY4fQ9zQ8JTuNbKbti
KPyFMNg5TESkTRRrds2Idd/rHrW90fKZ1/FI/msy3GAdg7ZNJRpcCoC9UIw+rxuGhxUNaY01DFHH
GM7j3pvSKw9ixBbCnpn2CIhGOthA9hZ+mcxCaD+Ti0qS8ew7e/DF7kLwkd1eHFPmNakoVxSK6olY
9lLO76YPT855A5VvfBdPdZbe5rINhVFckRHjkRApPzXdcNYGCgBguXpi3XHKPIJNv4aAY76pLON4
a0zeTYPDnnx/d4MB7ocLYAKXxPEB+uxPaiiBQ7Fuk7YszZ/cV9Oi/6tvSxAi+pZdH5Mqm2LHd0ub
L0+W2zicWBZ/xV0JOb4VUo4CoHLfQZi8jWKEJCG7LnY9U05Z6gcUrpJ8wGQTS8Gw/XgzusKmFBAW
G7FnnYBN+Yk5dFHRHX+cvsKYmMUizfqp7XWJ7+DJeHQnwSfs4UUe73GK9WItdBKSiNpkv+qHi5yp
uytosby5IJEtzsb4nNg5ZPRYiEGSt+vcrVON3fyu6D+wsl65/oNd2STMf5tP3S3LWB9WdN17UmaI
jvOCRLbpu7WUbJgi2oM868GbkphHFx4omFoocBaMhijftGue4W6FyFIuUUrlPwSFEkxwLWQ2nR5h
MbPYI6crXOUlkmw1Ae0w59Qmn/iqv8SCjhoSPaaaxCNm6e5FcNx71ehmJOt/3C+nuBzxjQuQKAxq
6KANgpLpnwWcLyjAs0RZasvzDo/s1yHFPivK7s4BIApPjNR6qTqvaasc6jOhqXl55JgXlzuEvp6j
8XsCGwiDzjNhBzlSe0YZoc6+cNMtdl/gpohqEUa+7THBPW706DEWa9yjP4CH1BaV6JW6f16dybe6
82YRZxgEaeLJMjI2xQWzqpwyV5JjA4vXBEO4WOeExifWL90WJUoOJsdsLKwb718IGAE2DI2sRDG5
K1nh08Le9NPdID34/LXLvaxbagR9JtLee1ONMQIPB5IHNJshGz3PEBx2zY1sN57VKpQP/vPp/sIj
d4bydlKYohHzJK1Btl3zA4us6dpR3/Br7K/T+yey/cLY9018z1NVkK6HXqLe6MjtCIBOTaQeX8/v
EYM0ouF24gxUDy4jdYs1VBRcQDlMyKAm12CwkOusvm23QlQXbNupJssBbpUKUxtPZIfk9HY9mXVF
fJBqRssHiYmHwVcqS/ZV4i0S12RqbpU8AlJMOx8EpgTHR0tklnqj80Bq4PbjASjSt3ldgjJprwfS
X12Zmd0mAMHR7wdNMs9iOrEJmL2EZm2HFPbA+xgj3UWBoOmp0ifMnI7rMU5WTMusofN6Qgc612Y+
v6ngIPQXuXPTEyG3a6WLUCwcrAky1pHDxoHExTCk40cXHag6M/LY/xIGaUeaScHXmC3lBnSWSXDa
pBSbTv6DfUwxRT3W0ijfHvdUEpTwNqofX5N+rXGBMpmmORbJ6dXcPtPxE3MajfDRASzLI+u0v6fe
D/OVUx6zvzeSf0OwkBcDowCnZ/CQJvJbTQFKbhIIJXN/AXgp0pWphaEbHY/ZnZW4IbG6eNAnu9kg
X6xyPiY/o1lW4PLclt0uEoRmURY9cws8Kz5kPUqTu1Lt4HLBlJpHoZ3pNwJIiZVWH/Wjtlld0yJK
4eaqAMWWSLqGmHLh/zGomfHxbOxjFl2Gu+zOe1zDEUDwfpV9gR9FfJ5ZkZxTkdDhe1/JAF/lBypT
GCsxqLbDkrT2itaksVeZG/RggNi3fbN+3BFv6EmB8hYBBFTygXLVg2Td4/Q4ElydBr0m+rVzBht8
mX0rV6fj7XPnsoGN/+XD01AXq1IazIsr3+KCk6T13Z107U83vpXSzaJCIV+xqkKYaa7bTEQPOtKP
OPd4K69gTRjjMJibD/AvBP2gdbYiTMzVBb2GmGgXjO+jzLarAxnpzplCSOYCUNR96l9/kNLwv5ne
pQ8aAXlbcHUlBm93iDrZJpcGJDuP1pl326d6lALsHgIbBHqlcqe65X7MxbeaLTnNnL0PxiZfNiUG
/RVd0E2+nkps3ZUrkE2iBukiXV5Vh0Vs49yyF25DYoExnwa0pUB3/qNEigfAKOrCRXC63RdOtkyP
XKInXnzkoGl6HQdYyz5T0CXEwrOb1bWDwn0jtyN8oarMM4phP79uooshTYLuuF/5R4N0jTZBO3aL
BGraohYtWbeNCPKNsb2IGVFr7uFurMDbyF4sZEj9pF4aiGWV+syHznSqtU+eBD5W1nIXFQ2MwnOg
DFzLY51dE7Bzgy/h5JiT3jA0V3ub69JwF/xE02OdfeCA34BDMlIy2ZHBPOPLl6lXZV/syrYRdCVY
bVN98Il7MHBU8PHki7o8CBzNqiFWvlinlNung1AIQjE/PAfjXk0DZiWnfaZaqQxLHjMwWkG6+xe/
P5M0910bcsxcf877pGwvibHKh0GuuEaoUvs6w/xOkeGMgHoRyu05BVmGcExol8JxRTSWfXEAjhGn
X54rUtx7U4mr29CdZ8o3iL6BgJOKOgLbexw2aCKcK7ESeztECneKYMs4wejoCORc8RWts+ILvydN
mqgGbY6tDK71YaW5WYTne7T5BJJb1zFwwnHIz0pLPlyBlwYMA5eMqsp+oJf6ALvmh1Yy8PoNrPLA
7lTHzc8uc4UYL7f4T7sNQEA7whNdeW44kc77xmgqMwvBE5gKuTnSdmxiTgk4nb8wc/BSr5gx62Tp
Fs0oxqSEnxr/KODG4OOCS1mpIqELywb/f0rVA+D1P6oifYoTisZGR+uJTJfkUm37sIv34VMkCLME
WfDhCBFUiz/aFpfmXnnVWNFVZmH70eWTHGFD0i2yxue200rnlMyJpnP2VToO7EVmfdSo1hMMS2eC
IFcam7MjhAOrLtIERU32zdKpmLLTBHF7wbMPkhcAoBvtkqKfD1mAX9sJTXReHYVE1gjTeppXOvD1
00TxKQ9niVa0ZhuY/hXTy3ltlAsA0ETNDj09EBZc4h9TUoYAn1xH2pyV4tRugsla5lO47pxvDE8P
0/tJIZL6LO+fFAjxngSksXzb+lMZBuRJ0GC/Y0lS6/s9oFUwdncA4YLPugJt6oauFXPaUwe40r1n
FhUPWAQBxKL3msjW9y5ncHBCJApTZmJsx6IUQZEVFIe5/gpIUFAgx0f6SSSqPlsiVDEyzbPCev4z
w8Bo8k+d8KP3hQj6wUw/aXtN+3HsidjcjD9wZiOtdsWmn59iVBAm32MN6ZOVxWeLkoBgHODodDYl
3w3410tynJejamQpHmEGNjbR9ZonD6nbTItefLZiiJj2CN0ArwjskICiji/Lot99qmq/FET3I8sR
6dnfKzWwojA4SE5IlhNF9YGikg2xIDvRnZv11TslL8FDoCyInCfMB1L2gwdPxk80jGeZkmvt8oVo
IUCpc3EZUZ3hgkkpv0/Na8AgXPP3bBYHWG/l5UtAcQmz5oNIkNugOCilfcT3WBJXP/tt3KCwDV3B
aJhzkjerKCiQ66QWS0xk3bJzmBMynlGoyldsqA2vDJgdfBKpPHGhb6/fZTRyHiIfc6si2uGgbRHP
OXPzEYIvDWuSagenYj/mbTCyaUuX6wgX2fDSabAyO22xxy4Ag5sFaGvbqtau9aa6S0WK2dxQ6lFa
PdZzazRo6ze0Xcv0H5bFpX3mMCVyHCfzs11qhccsD/2/DKI3huFi/8MFtcgwSAGIwRZf3JHpCWla
zid7vJ+ITy97zKBkqYG/Hpo2wzAwp5ARDtVRWkL2sFOHtOHXQpBoBOH8aFuq3yLrFce19RGWjbI0
BPf5z9B4L3Vvjvk3vE6dsBWQ/U+HWfa0LuVTiy11PdzzCbi7PPTC4e/8D2EztJL/GQSgAuLlDgP/
+3mLPyUALoOINhViXVyfoxyv6AXf2NoSE9i7qlb+dw8GNbyEEDVz7oZ0BADgd5anZUkxZdTP4G5s
vlpnefJ9Ws2jCh5nORmykuIITm6L3o1yWcf1g9WdUeENAxfc0kPjYsyIRpllPwGkFQeTkfVLEA6P
wCzCzoWvKQuDJgqn5PcY/mGuZ5Q30+l9uOrcgAelscZZn5gaCbz1OksH+IaDSVOi4tx49CcOPecb
kK6HNMUJBYcvpQHJbignLGEXFUaEHybkUHJ/JZvMT6b8/RyAdoZp4hU6HAXUXHLydEzyOIY3ptlo
32VXpmyBLwyFegp5HCa4OH3o04M763moa/jt3bJXukknwflTW3yiJaDN3UpPYggBDkYts3sl+c9j
hS7sdCgsr4qqnLm6ozofmio26aoC85Sa+/9jh8U3g8AZxxOD6d5vJB8ifH04Pzj9sfeVRuZENq5u
E/Ukox8hg+IyKImBFzmBHObQdNmSVPHM8yzNvMqZJsyIQ1BOQl1A4Jhv3PPrMqDKZ0fM+lBP9iLy
BDCZ6p/b17zuwEVD3TO1hDG/igLA65lK/+6spmsb2hedt3UDh0bUzUCDdkIVqzFAQw1kk6Nq10FJ
Mz6aoXCrSQywC5CbszZX1ZFuDExgW8vOtHcIi2NTEbdqlCLdf0SjIbcCqHIhb/CSD0LKVlZMQz9l
wjgDdzogGWpugOA4Ylc/mwf+TCz+aQn7YxUWFGkTcK5X5UzuaCV6chWQc3jCanqQzoRA1c+4+0X7
ksrxkcXcRqJ+gj1onqFOClTvMNxzRjTMF5mxz9KiLiJ2lYGf9BcIltYhvkEumHUX2/WzPwNJNbqH
v/GfM1o4zD9BooaPnUefolNUMi8In2Apnfg+Ynl8I/RVhyFDuv2t5og/O1OPcrgyi2zgoIY3KB61
zDDRSi/bcDS2bdEhT31wGjtTWMi2nL9FRT4JSmSS/dp7X38/CKg0NhlC+a59AuQkhLQ8HR/4cuUI
Ozp+a41DHY1SJGdCZSlQpam6mDoBncY9Kpg1VR83G+O1B8YDkAn/fTWdlkc2uhS85773jmtALUuj
UFoFKex/zqervmU2crlN1Sfftu7EfR+dVDbc42Q5RySievK6WYLY64Tb8qezxU5RH0BMpCItvAFN
+rfz8PWBz9Labl7Hgel6MRJKKC/aYTOMibc+HrTi0l9w5X4Q9sv/5uPmesWX29o+votFSiPNm7rK
RzjZVVOlUdqWrJaVPHvbWpc9u/Cn7depQH1p875bGJrj53q7aJDEMahHZk5qX1MGHjZOfKwKCOWm
guEamPUqbkEn1W6Qb87xiDaTYldTw63L5q3Wf97dtCPGCExSw5cALckM7leoPZmkLiAV+0Nwxm/U
iiq8TamTJWMIcb1Nh0R20AlGeD1l3PWmXt7xsLaZ+x3smYwyAMRtsCbS2NX/4LQ2JOn+AA/w4FB3
ZRLe4z07ZIiOuuYVx2XF1K4Hc+Nh5E6omvgmxCgoA2xN2tFz7npypIjjwMyiVX50dDh6zXEawkBv
Xr03nwHQEsTQgFdyAzcXiwECRlmUFFa6aLZOJEC9ZqrYdeh+YocsUbF2QHmr4ddZN3JGGcQp0AmX
0pvH93h4furXnufNrczZ3W9Rke9IWD1GCe963aamtuNeKsRCZ7qYDRRC6OdhHiwckXNaG8qEUYsE
JbBYL+IrOtAWrupMODlcKS+g1reifVCddwDMoO1JAPCzEBJnsL36p/kwWTQfWLc0zvQ1NbawTgC9
wNF82Olwh76e3jBRvTfOT8UnC4/k/8Ds2e3wHLwB1wCBTFILzYhBQlt2Z1D0WABjWZWR7xiaYE70
k4KiKTGJyAtkS/yRASgpFD2LTwIpUhUkjX/970PKONxUS3KzyjBbX7ZM8ziqgz0SyQbXurQEZyKs
PakO6+xUfN2OKXWYesJPZChpbVvsaDZ5gdTkCMwy/onrKyrxkNRC8nFeiAxxM6vj6b6XMwlfDrq9
p2RCpnut0gp3wrlU8nqNu0yAkTRMvGhfS+/9XX1I+ZxuhwepgjZz21eKm9bvq6W6Nr8sUDqHFztA
tO6jsNDkfkB4ihLjTIznWkBHTPSjbN3mEXJCvqoWdskQB04+aJpQ/gtA/vvVoNKOOKy2wCh1hyjV
p6oYNx86a2qJTplxQ5S3tMSdjxQeCj2qA4bI80HqOYxw+rj5R8JLnYqAfSWqC+FpvSXCN8l0YVcT
UIfbfXcpBPh9wHGhVb0RcESutBKnQiZvSrZwsk5me5Ak05H7xehkGNHYl3ZN9fAkeavpBqKWtVIC
K/2vwR7kYx6My7YQKdTmGQXZR3UzsaxDUX/VcjNKwCpwdBksNmZNdmdsAhfm0Vy/ADTZvTtQYVVT
CWi7ehWYqZP3H8/LynkZBmoxoSNaD5dPSNepySSxcsBWJGzkOVXiwo4VdfpmpC4y+z26Yqlvw6sI
h8kjw6aUwvdIhB2vql3sk0wvbWjwiCztuzq2Nip6CafAxc1fyZrVO6mP0TllXNI05URHhKaOUi3B
R1g4XVr0rKBa/H3i65IPpYR5w9fID9hVt/Uqvqxpyd0RSUIRb3ikI8jUcWzc2jPX75NRkWoUFqJ3
c4QPCalZmiTXRbCXFrIE7JGc+zd6CnK2DBpPXJvf6IMktQiuEl4YmLzg5ZxesQVOW8ssmbSGaLK9
5ySl6ZDZ9x1t0OH4df+6tjSZsJ4kcmuhqJK0B1/4rA1ZDV/Wk24PXJOqW8HyYMtAx1+YFN8+g/Oz
WTzdhF08sY4lNI1b/+17WO9dltLhEIeQCFYwkWA8HFtAQpURR6LgbTBlW0j0jCCescf1zQR3jUCs
6mlAT0g4Xs580H7Di9svyiOUn3epMCeWxha0KuyL+ax/FF5qFRXHq7R7y/gzMEiTDThm5lGStUcg
YrGSTwOM71f51LzKPzhq+FBExBwDMjZmU+SPgsgz0IASgm7vnJ8boHr4pRNvsbnjKDCqVPI11YHo
uCKpGruHnWKpukK0eIqKh4T0yfIB/mjXv9eXTiumnjG0DuAbMrE9gHdITPnz4hICXjg0gRyuw68F
jlFADoqBxFI+u9Nmg7lRwqxG5iQBSwUwGMNEqYYPE/c2v9F/eoeHPlIBvr2+hLRJ8V62IVcF6ZQh
JOvqVp9eTi6JV38P4MrxYb++ojxYMAUlEvjQKbt4RebaORWQZkh9NjqUlroGbCwuAxHCqFWsjQSK
XstHFYmbLPDel7wwbjnQL44q4qIKqKSSaKCt6uT4jI6o5BWmL1Z2JWF/Gf6WmkA+z2c8GkjoPAF3
vstpi9091TNHDEMTGivrDNI6bVIbdp2jSxd/mVFmyRj7B5O8hSZrcsWV4hbTGQ3+bY9SUPmttwG+
s6v2VThNFbPmaD8r1mmTAJfU2339rTdjfVCpDXZsrk/gb5vT+Rf+3oFiiGii7pnCOjGUvJg7TgbE
ROw9wc92hDKH/4Ebsv+VwHvtJ/jiu4D2j+7g6e62z1T1c0gFxVCu4CizjKy+705cM84SQysRnMKW
VCJTihejyS3dcfQR4nsv8pO+gvSa9+1eW1gGXwRNkraQLqr7pwmQFTRf9YjUdWtt7bxQHPp6Dyun
md76P0iz0E3p30woX2mO6wBe1bhKDIY5bJ/9lqOnijVzwte3YTuLgZWnLVWPc6wfJREMgBMx9P18
9ZDAm8WsL3XFYN0E6jG+4IYL+VffdXGCSDDPE/BdcUv7VdDtMfOtvbf42r+kYXe5gU/aRjOtg6bu
hx6EcU0z0n5cOORLpRe5+7r/FSm3GFkuCtSk+HMtOpTrNKkW5zAANZGFRRUVYyXnuiXBYNiTb8UN
7j7tbal4wvw38GSXK2AAvO2ilnFNoxbZY4m00+obff2rLeaX/kjY1CbgkUvFibZmxGh12jWeO2CZ
izo9hB3rToXjE0q1h8wR0Wiq/BFOcfN2CK8HIjObF5+ip/y8ZYRh2Uklfe4ZqWBr5Dr2Ol386bEF
bWwcRpvMxkmXz+Wo3b/ORHcRU8aYP3gNg887Y54FLkHR+Ao7s/1/4sQRhmMuW1nTUcjkmETKa7/D
wS8uutnjALwWtqm+J3C+xVcgbCzYSXQ/U7oc/MQ5gTR5L83qhRFngHwnvC+asp5JWsIkHLaIK/nM
D6eW0zGVfTzk2zNTFPsdEYVdMyTeMfzorbm2WUDLcCOcrR50P/tnbRB+gyYYaO3iHGa/8BMYxr/W
2XVZiddPQUzzz0b3iRmRZaLTHNl6zhezW7PcAeoJ581B9i4iUH3T0HTezvOyWsp82I565FYgHLS/
Z9w+FkVasMh5r70DI7gDSpgwRFhTMAlHy9JAtcKJpQyjaxleZnoGSkEDalsqhRWKpC7VPhR5vO4u
bf1VhaRrYPVJEA0qV5Bpdi+r2WpcGzOjp2NDDQFDsmBC/ggq3jTQLqIsR976qjnl3AXOfMFBynrh
i5z0TelmPoa5NLoi9YNw78ezcYFQ/i+bhTNmUwwyBx8NWJxDnTw0Df9WKLx6gZsME0jy+e+sXCSF
F/JRW03HJMkkD1K+oGRLWOvrBk5uzTE6dx/mrOs3TJ6/sAlYAdfVbW10j7D7i8xeYDcORV13JGtU
ihGqAarbnB8OdeZByZVnixadm37S38bWlLGTLzHRKTYc0BX7yFGiYOiTWZIGuXcY9VN0/8HSqBd/
RZJ7Jl6Dp9tioRHJ6ak78l69TO3w7SGxDiEBXx0NadcLwk2OTPAG81KMnCPV9UCUTepd+l2vY332
lbS5GNoxKkl3utYiLKgLitChOPVfTmShs42RXikEUeLBnnLs22mGPyvXUgWfxP6zFJL2aUvRPRPd
VE8Q9h5fZafRUpRznF8e/lK5I4nS8zGe9bzhDfygq3hlOfQcwSaHmdZLKsaM2VF6WbIF6W2bSogL
amj89E7indNaA3z91XrYS2056IwedG/CBlIhaqZbBgT1BAB5w/SRQ/bv9JBTCOzKovyZKz+WJ4m7
0+DXd7hA1zZzqngX3htACnEE7DMABLzStdGDIkr/8t8PbdawsyraIpSjmQNAh36lHKjBG6svlYH/
nvArLGoaEEovx9sVTmoMZRgCzeyFx4il3AFvBa28U1ZGel8h5NA4HKBiV8jZdYFmWzSeD/2BdTJ8
oNkA+I2SGbM/7YW68cpeQSwXx0BNNpP8mh1odlbA7qVzPX4ySYiKxwOMBPzY9HPrXYLaQv5M1I/7
xrKUjbmTsfMwG//qKbZlVC2jM483mO2mupL7KSqMOImKWiks1HQ5b462445XubrIYJQBQTC9iM1y
wn1f9aU68jub26Kr+pYq6wrILAuqTo5iTjB+P3UM97Zi6vWS27ixk/GDvsL8g/8DUsyyfZDz3DuH
kgtINjWqfzRsbf95I1gxQZzvvnBofHiESQ3/lEkQVCNGENvf5G/vSdR0AQeAZpJSBMM4mLsxbA63
1yMlz/1IokV0aW3mpZBTaHrhnJUiwlLj18hril5ID6qDqirsYj5jhRGDeF58M62ecRn+yNwQoCZL
uzP840a4ewK8a9XQ2w7Adx7fB9FSF3svubUKq6a/1mQ9XBMmvL3v13nB7/zmR+Ypbcd+brEow/A3
MKr/1yic5Tj5RBkieLNv9u9/cz+ykzjYAD6ghJt0uZAalRsGqldjhn69LkzKz1zdpwOy3KVZVJTv
5uUqguG4/70nymWnOYYENzD/5EYTOgnQRs1VN8XrHFj1Sn43CmIW97Y6lexbbtzBHD3/DhNdb4PJ
f1z/FwiQBJL8qCsxP0vit6D3gwky+QUk6Aeo5SZU1J9GJ2F36b2mZ9brTy0Eh1sg8FaiIMW1Wc5A
06LdrqcW0XoKLj23xRRmkKoiGMiRhOyMa0YAL8uj9J8a5xP3NoZMqVVvuzgMk8u4NV+YDLSzGCS8
8Esc3Bv3IqW2wgUcngA0xcLdKaCigwDNFwulWFVmqZ54ISAvLEzCqq/UZi31op/DcuJVLHBUmQMf
mkJCHaDyWmbPbVvOo5IHDtJuMYMwsjwyJqyAm1zydBaMGQnGU0opWPezrNxaCSTiur26hmRu7Wd3
0KHNq5c4D1XUwqfkaCwzmu6J75zPtguq9/J+fe2UQqWKCTgj3aPHdCTR+InLoQ+56pQs5r4TClql
p+xBiPzNbXv3DXeTOsuzEFh0BxbyNYk1vn9N5AHLxGHw51jPKQQdz95jiViPL7AMJaWIOBI5sEJB
YR145YNwOtUh/qBeenHJOKfQhf+kaA6BEsNFG4bpioZEfeeNtcWcKFSsU82aXzRtuvQPEvBcLMAA
YsmumkoEbSpGbpW8oaW1uoO60FqH4QgHrEo85cOwdpcggmGFZXfDCjrEkMpzQLhGGnu2yoErdgX/
E6wJGj10oh849rHMXXoAXRo6dOhm/6uVqan3F4w1eI+3cog1XKbttjuVPALAH9igfGOIQIDMtphK
JlUZ/meyOc9FCdLIdF59ZsDj42lH0XwUSTu5A2tBFULFoGneOSksGQW5XoicumeuVssOWHssRqFR
6pVOux//Pi+AzIhayRIvol8p1nk1yuQrauGp4HoJuvPZUgw04rW3QS4Kj0r2DEXsXRKm9qMlF1Fb
NSKp6j+V0y54o79SOt0hZiz+391Ap6ABWxa0IL991e7SMIM3DXzhHZFX53LRU9CSGqVr9md0SHhM
cdsa/k/3fAzpGLB60rp7Ey+0LUopwLO8ibXVTGQymE7LIfBY8FyhQ3+TOri1TTX1ACuewaiSiI92
3RQljlGFAfKIMozur5sud4gO2Ed5DcPCWvVzS78jxauVGKgUfFOQoc0Gdp/6oq4cw/IeC3f/1IkT
iJ8czvAfWpxkJwZe9jyqOJDNmB1JWiv5Hy5HC7XPKrAhsz0qUeN92P9YEHc3dkGww5Q1eVTppWEW
G3STBQGH6Bww6G2baMgx+WRirIyqhYsAXauKqAmqnmgIH2OKH/BGlhPl64wszA4S2/11I00EdkMv
T4h/iC5Zl3cH2UDTxd7nMI1qnOd4B/U6WvbGlj98rD+0ISvj+O660DvGBoSskfv2Z2bQlNIH9CDe
gZtIwkNZsQcyBRYB/YaHTnToaSkaNeB4UqV7UOQOS38MEbfvWFhf0RYv+6oIBRz2hfJ/ICRnRfAe
MuVr2EflMBQTgQ1KKg20OurmE6cBRYqKuQ7OcVY8S5D6Nn1nXHFWfHVu/pmWgpDGVTy2IFfdGKF5
c+A1fTYj+Kb3kLEGlxdOfbeOU2bvKv/iBXMm62wAt0sdup2xsvXyT1o7h7JOnE3Sr9hZb0gwjs/M
EatOO7r8vEYNFyWXXjY+TvmsJFee/R1aYfpkXIgvLkHmG6oK5hgbODgf5hO2IhIIo3ja43ls0TDH
B9okIUoukxskpIVSZCUIVKJ349pSrYI2/Z1FgYINfUi2Te5vu21+ceSPMulJ1tT1exQpR3NxwXtX
bcVT5QdDzy0oNdE71qPRu+55hhLJBzzKX5ty/lOXRHLuNG+YSf6VHdPQyYY8X96xT2ZNEVQJtS+t
4mG8uupkL4tPVaSmZEXPbVKUMnrEhdTpOolpHm5eHH/dCGolH7S8nvC2z8Rg+gTvu4IHXvgSDqHQ
m+dFGPFG+MnbH6sOAvBJowQwgs9Gm80nl0t8aJgXoLNsAVYbn230ZK8t9EZdgfapPOvIqRSMY0QN
9TrJjF3FdzBN/pNFUH+GL/yVEtdi5ld6Xvrc8EUr7yB0s4lpCiPj7DolUIdAagZG/oEc1GUclHQG
rXImrWoZa4yq7Pjc2aMRyEiwhhQLex0Pd8REyxu0sJ8bpvMKDtqWcjbtf4dkVBHu9+iDzSRo4X7e
kKGCOoLHgCEO/wDbMRScPQv3AxJzlZBQhcFZhnyIo1Ig64fo3tj+9FTzPyjvxZ15UfdfK52mZoT6
09Nt3w1c9rdPBSVh4a4wFggHWxXlbq3EfOpZ7JkJt8UTxNLndviWLapWnHCKL4Ay1nIRws+iGIOB
8k+sZEvQp12zCaU6eipB7PNHeMgBpwA7X3ssZU3aGB6r8MeufoAb2CGdNmvUoMUy1RsUYhLYlEnN
DkwVoF1aIBrg4BZi9vE1OWoBARMn47L9lXsiJ/vcON4QDEeBuas4OCJLX8ewDzpt1xUYgYtDZZo/
1G0rBvOwfEdjloG9Gu0mAudso8q3SiLW+tPdvQTpC5kpIOuIxtjvDNPab3rZow2WOHMCyA1PSX89
hO4jEPy9icPi+HQid5CuLDZdpdzNwIPJRNMUbwsCTM93MLHPu3BgCk/9FL4VXLhkT1GdMnmPGqoW
ZEGvnB0prEhBfpvrAPIpAAQkzcqYN3cdQSiMfwqhdwHvAai6CCKmNlln9Lkphlyi8rOsxy9OcTPC
Rm7uQuLxLFa3Q9tjoXHGOi4aNiGXOWLHYxIgu7RSNOR6COs8F/9VS/S9AR8Ta5sthpmQQOiOF35L
mXvLPOrGIYR8QbFplcI8PLrWvJlI8/MshIgruhKlygUG1ww6FHu2XMOdX73oK309CEOmRtBGeHLu
FnroiloxCN9vT/cYdTtK2dSsdRYw8kRezhzFK2pUZCjR1oydazEw4wQ1us3pSK6512bWg+H+2K72
PnmQp68QXGiD1OfJLDPgpTJaGbAFwOWKzTnMOC+XnFzWXNalUuA8EYXp3befk0NTVM97Jg2ve7il
6uqI3CrDYPIR75DFr18n+tFrRjrSpc+aAHpBTxCvSd4kQ36PU4w5dKHpskGFPiLddiF+OaJ0j7m5
CmUeUGH5dVC31DZzDcqYtepLz8CMR+AiokGVL5xPlZEuI1wbzs1nsZWfh/NIBbJUd5gn/nJd5Ntw
2MkWk2jB3ou/LuTZWEdeZWtMihLJGNVYUvIZliBbuHnQtFhYiUaYqLJNjHrp+5I8LFou74Rskc9s
bGrD7bN9vH601r2RqpF++/JrTXC4RhxjOufSA6F/lkHYgclpavubmA3ddADh6kcx8qNZva7e0qHe
PUxBPqBtJbxQC7TieNe4HOMzT3BAIzruRVNrRuGVJnZd5TvCQ6ZcJ6GiG6tNjO0+oJwf34BT4sHM
sLNJUShhp2WrO6sh4lbO2dPumQn4PNErhXD49vxscBtKHWLWtnLv7YVp4gxWHK6GadNTN2EnALlm
+WtrTKfP14ePxHsn8ua/WfZ4ZZRCTO3PEUAu23zfykmHgyqKtHCf3ioRqNkWl8bRv52AAiZamaiF
5rfid5YHwmTtSigv/YPxNus/si2ZUGlgx0ZJDhYIVwoAHU59AeH/sxHJx2yseF9y+6QBpDKIarW1
vNUjo8MygLk0uR0guckkftOqjz75tucB31UMAoFN5ohqXSNnFaoTLjXRt5F55ZDFmniIimcHyOL0
YzITabiR+IEDnQxNxLA69VjUAUaz2s7aSke9FN34FGi4LWQ3c5yCat+S8NEhWU536ZpAv/Bj/k6Q
jW1k+lnLr5+MHcTmKYormeJE1yrW+TvMtYIWl9kZ+uaPMj/yhgp4HhMkVrzGIAtholwvzhREMpEG
V9iiGVQE+iXOJc5lLS3CpxRopw33e8Wa3Wfjk116+oBntaDNNk8bx4a3Erhmit/JdcFJhTLSPgyz
KgtWL1gWWCJK4C/Mo/Q8jSyxGHTS78RPjxDqVzNYRhCY8sPdIWDytrD19APtX/KJfGCk4xJZRRx8
0ah/Kp+JriutUDsACwakX9BznUn1B0FUynWbkjCR5eeCmfF/eklavh1+XdHDifXFEzIr9C4C7wnG
m6S5ikJuE8aBw1szkaBl+68wOX0IxAnw1iwiQoiIWiyK/AD27eF2Sj0fu1/0L/iaiaJGhN52Z42Q
EfKAPqO7rt/ElQbCgDxP0E+KEz1/AdgxTqIszzjlji3GhOvRr6dh+X3iYuTT2oz9SltSAu+OzMR6
0NSnIBJolNM0+Lt+UKfBjul/IqCQDoKhXfdECwxEDZOO8zDG9IGhlyDGeXv+IO2NJu8pegZiHRRZ
5XQfqmKVkYmU3Md3E4DKlpLQmzOM6QFZadN8P0Tyfev43sxAzEWGpfxyP2LJYPRT4Y8RwLXvwr72
UbytirSA6qC8KgTs4flKmHeUeP069ViFk/lTfcG9Lny6VQ3xGpZB3JVlgx4in079PdVokKwr2cWW
HYZtpyq7jyS6iFhluRdTT82vroU07jdU2dzGFzCVlL06W+qsj2RNx3527ujbspwv8v2+pZruqn2P
6qeZuTaK3LD2FbTQw3h7GauAQPtvQzS6k+WmobqmlMQatJvyxY+zA6T7XswbBoY0M83Am7eBC6MJ
NQY6xY4rFA4PF+pdhrXvJvwxJwePVoUUSMza7SJiFP/KbUGZN1lXE33eDZLftrMNze6lmFGk0Fc4
YME4IKUMD6TSpVkFI/8wx3HQH4nnVm3KyNZ9ennCjA6eKaP4wQXDtzinbwGCXp4eHd+b1Vi7zDSr
JGgCtr5RTEPG3bBWOKitfcAEuIZdCmCv53+j2GGWKgApqqBaxa4po4c12hgM8/B/uNMO9XiBH0sb
hgWzY8IQXQA3wpkM4W9ZaegiqNCe+Id+iEtrh6PZqVhGlaUk2q7l9pqDgK3GACuUEuU3dT6BHNr2
dOVwED2vM0l9R07V1QFpy6nkK1M5k1mXy0oAF43Jhs9petqtCa7CmZd4EZRjtwGKtiuUt6tgQdge
0X9k1a8H0zhA2ZneLcTbmPFqEvcZG7D3xyVJuK/4tCQJ7d9EKzTyFT5EAfgXulQgio111M1IW9y3
QzQ/hdTQsyZ3yl+rvHqx03RYjWjKPb+OXElJYCnN5oMp2t5SXgJsSjOPGHYLHabRj74vA0Ousi98
nicJawwRX+c4TxV3V41lnrsgSyqDoTkmlNGW1n8THKOKlT0eZCZZyTBHr88DMIbuUNBAQEltrmSl
pR86am2ytUelp4AWuUxyTcIsSLBRPMxdlaBX9rhw6dI3ssjpZ60iYhnU34fJjZjAkre/TDnd8Gl3
kYttBuhZPz+m1BSsfGA732eu3ZzZMGaNsEb+JcRnqbZ/t9/eZkEH5CkHTh8HVj26WdSYdqgG4dl8
mrnTZoYTztyQ7QH+mB6gQBnavd3i5ZkQettbfgTt8AiqSh/hMbJZTnnz6EYxQw6/tq83g5lWXgdb
TYG5DXJYfh5r6ZcKvBRMPzQ+57deG3Fdd7zdhRlYjF9XHq2bkCljbKERlcXA1nxfZNtrTnkXHC0O
CumeX5xypSFdvG3W900PZ7AqGoUrOhZkBBGYgnixPwPEDCFK7VHJu296f7J3DEhswOAb3Chi49Jc
W8gXVjyeJLP/fvb8JWKTfWLaLk8mYR4Lsyuv027ZROOHBp67T0lr63RAJAhr6XRCviCgAcujAYYW
34VyBo6F/R2TMw8NsTvL1HW9398gFV5XLI69KOhjek337cfi1hY42hcg3RFvOtszxblaXW0ncmMH
7sqDVlUAwGQqj3JIwQMiHS0jiUH8y/Nd5mkMpIrQ5dh4MXm1dGZ/yV2oxrc4EKR7Ik9YNY0vikRG
OSJ0JIPbktqhsuzXqx5OS7BSbxHv2boQ/mo49FRTHIrY+VnitW95gEi18fFC9YHM6lAZGTQHenfs
905PwcEXxffRQeTI1SHeENQEnqZ+DALiDU2fuIeF49720fqerqAw6HHJH+vwhnGZPV0kQ7mnG0np
ks+BSGjvSlVbV+67Dk/APrGgcnbL0TsTTHPanvzzHLJduR4FmbEVSh+DB2n22jJJUgNQxjfd9JtO
cdvdN/azqO3uJQYJovykefYDGloeqrQng6qPrObSqn71BnO/7dxM95jhpa3HQRLqQnBwkeiIjgkt
24FKb+oa7LpPk3p0ZpE4j4eYgmMCbSzdMLt3ME+Ymg3xEOUhPAHspWpe/rLx28oKPtCxWkjHLkRO
ixfDKAiy8Bdn6eEs5kOuly7xf+Q1W5DqvO9zvmZAS0ADsSJBAl4U9OFr0PBM+siVCyCDZfOfzRHd
7Qe8CgEKeGJww3RrwpOwTCDkONbQVf53zlMUk0SMtu8qC31arqzqS/mcc5ATEIgjXuffFQH85Oa+
GtItWzS1kCP8+iGinON27SmIKmyDrNkg3ErEsww1+TPyqxahg9tpj388wABCNSAnoxGpXgIAbyjV
30F+orUD+s7a5OoEErr+tzFvk3du0hB4KcKBx80I0uM4xLFBhDeUvcdqgoXwVjeOGMn1QaiCiLRC
HngzoVb41kJ1699OsDI5SdwnDuvNXZOdTC7+22r6fJfoL6QOhRRvmCIRG1mbvwZThRzWYAaaaM9o
ECT6UYYNkJfHKQQKQvV6+hmiRxZqXvak5ZASec9esvxwulPQaVT05Ac4uRxMt0KQTAix79KvFIjO
0W7p2tLoelASsqHm1uCnYyc0T0BK924zy1xgIlnJSBhPTYC+F/6W/+3OhMPYC8Kdj5GXEgXasnuk
TjC2FxKqYHirPYdFiqOM20iEzre0qC0mt5qkZ2RZIl4j9X65AiYN3IQPDwc8pQWYveT00JvpIBst
EAk1uXSv9f8QRLkInjvJ2xZ2awojj5xJl9ZS0j+vIKoLU6bP+/FpNSpAHj40FdNOblCqlxtABIEj
1xhoPGDzS69Kt3CzvPYbtaTess+/rQHgbrHNpRFP7iBRKRXyEMyyfswyXfaWTio1YKtnhxSMLxz2
YmF7MA4NZDuYZ444qI6fwuFpjQzslM9T4fP+CgbROwxXCFyTpYybTKn+FUlfCQDLCn5NhvXTqDuq
zIV8wRwoiHmD5RK92w1j06LPYea6aTiCzqRS1orElAmuYTfbujj+O0zK0AHY5xxf5FuqMw/w10kn
s9HzNVoimX1hBx0QF5u0J+4T2vyY46nwNX1Cnq6D8Enba4scp55VtEYidIPEvA+gFqrP36nWa/Lb
gB3qUXDFI6sJDun0hT1NONyb2v5DDDAOtpVlGPUBwaI3o+wrwm5UvX6Qdxw7VJfCbQ0hCnqrFqQp
hrodKUpHQflTeAYBkCmbVLPkbn018nkaJNdKBzKOEglekf0bjz2JBV1P7WjdCZRQBkFus7HKCG+N
lvpDyPKDk+5kho1mQi5ZJDX+dLYlstsIA2t1yvj46hZvbga9l9Q73TTS/kY4cAyAuiHYZu353TIk
lSMW/gEAboODcyeyRaWDdCnDfu1NqahcoOCbWklPYWyrJj2TePI2WKsC7nWpJI3qOSVkp+VlUCwX
k1b8aBeR6BiLZ42kmoJKr5cjxMOzhzmmRRX4ng2+HKdp8ryJEhwA/SZvRWWAzPc2g9IE97r68EOy
r1QM/hL0TNiN8cVxtL8tLmppS061FJHnGOPkHA4mtdiTzdpTy+9CumS6zk3q0/k6GojLNyYOTC4v
e/d/AACvEB04PKnrOK9y5PAxfkh+qnSDvb70TrRZqXUTT8m6bc11NtG9AWWpqOW9gpEs1if9x5W1
LyRVFDmmb9bKRcxPjJssbnSP/PcoWTESR+9AAIyXgg5NFBm3T8Qe/PTG8S2pdaSAOYjosZRe8do2
UIigC3gj5dkleCvFK/zErHD79NOZnhH9q0MM/iOIfv4E/0ymchBdEYNrL6ATNBOijcwhvb047qd0
r41oVBhEysujlimLLaB7x2PsKmLYfJNbYUAGV9HTZzY8JJ4GDR21ZtIAiq3Dv/1C5ByXTJa71KJQ
7ghNvkpXs0Uf6BmWnZcOkiHOZxodW2Zn506+rm5WRxhsTNd5qIXYo6YMzrzfdi2SOZsbCbvW3hTW
bK0u5LpxJ/87BiCHE9yq9ZfCccBkKgocjchf9/uWL0XvfuifgEuV7Se4gVnYPSSFhh8JrgtERdh5
4sF5InuIkKQtP9nEwNXuDY3UdgaJ9XrucvmjZud0T2nzKJY1tTxvC04L9p1wKojwZB4DCMYpgX7S
v03TsYqIhP0CqGSonSL7ko0cpCD4xIQdlIPE1LuOnMcD3pEEFdqqHXRdxvXWsXoAgJQN/8AKyH5w
N9wCDxoNm+6SUYmuQw3fzJoasB/vi8605I+2QGI5KLXmX87jTSDbKlMNnAKYYo174XAl69at5OwO
1Tb6hfIwGRi2cueovZDtd7rGDL/0eI/d+uS7a/yutp/25h+3X+LjjmFoRwKLKZqI7WcjtiquStfK
Rou4VBeAYnV2bjDXwR64CKI3gjphDpEtyEwMagvfNI/X3qiX2TtM08gDFKhMIf7TwxdM4fLnt1zz
b5qIJH32OkWFkNTTUKHWH6A2ZNygXrJgTO/mRRlfaWovufclr04bRY74oR0vgekCsZ14GQlResuM
gi3DNX3iJDikmcVWS4SFPH+pqFeP9N+XXBr27dJX6U+Nmg6mOrd+i7jMvfo2HXeCBwSN73HV1rW8
IKTli3GAhUrFDAhxvBMRe6Yc+oc4SFTL1Gt7nzcGo66sCxniIv0ZcgY2VzbpQQuH/Onv2LhJvUKJ
iKMRtVioOwOY6vDX5Q6nHTqQ0gnmot/ocg/lNN90vsbTqVRiAdm1FXYN8AgIfzNnl942/eZaue3k
8UMerhIdxaJNFXDAqQAWhOxr0Q+qehRlpmFwRcAM8TsYmX5dkwgEO2s2DcGCYqQBHWK+l66TGLLT
uq4mohFifDCjt5NQbmQIYhHQFms4wB8UUvPlX6sdPx+bGiUkYV4Lr6CW+BgW+Z4bVUBc+4E2xm5S
pvrs2p1hTh/z0ekWjka9f+Zmu0cnenIOgrW2KL9T1saBmwwSdR66Br0Y9OTMp147mdCPqQln9jcS
eaike6yr3CNvKv/ulTX8o148TWs0W5v61QeSBrBIYIElxvPykYy5xNOsUWwz4mkd44Mh97JtCNHu
0U2kk7cgCdCBaoT3kXTcSdKwa2ZwMTbR1+Xb3XO4xK30Eq9iqZ58eI5SiO5sq8nauA3M+OCuLHYT
J944wm8FWJqEJ9Gf3hICDGTW/bH4m02BSCk0fiuH4rIQ0H4LdGrsJpAjiHbQiUp+bTSylo+AUKo4
7d9QlBmxtEQTRtNNEr0zH6/m/585Wv9/qNdPem/EbWVwx62fWPDuy/TP16c54WTuq+7QwEaCFZd6
52CgOj6gBm2j0pTvh3q2wq9zY9i76f91LX3so8OiJcAI3tZjmE+j/NMznDDNwsDKIcP/Uh9KAeJd
jzGTH1LIfYXlxcP4+JVCoz2q8dSE08SpKyEzikAAMyE9rUKLgRo0Z9EKlQZoBxJR5dP/oJMSmG/2
yefEP8UGny+Id4o/4+8s9X9yeStzOLtfkH53yS4vU1aoFPKqxN9PSVNReoaWI0l7nqq920ccbDjM
e+49XL9AcH4GP6QR3NLuhuMe/kManFKWJFrpYVR+z+/gb1uwu+sRGdkPs/i1EAUHLexuog5KuJvH
YuDTJwj9cem4+birl7iUsFJpyVF2KlRZrHKaXOxoFzC8TCu+yQaaAtKKHtoqLlOlRbKKZ/KJkQ1w
ecbCijYT4h46fyRu2nmhEjk6+j+Vli9j1vgeaqHq/N2sxkMPzl1kgH7Qbic5lKPJZn1ir5GIfaFG
EjOitJ5sLU7y0p9uPdsSIoXU0RiDe/9l20VeT6J962Sh2ld64ZI+Z0cpwLz41Ewy+nUilTipfwfm
dtYhtFKyeIl7dNgKGcipT+c4n/kWLzZsuZgoir+ylHYkFYV/SG54eh0LV8ns1oRXf890cCR8sSM6
JaCzW7DSGWVqHs9z/b2np9d06EBqADVwux9pFc/0UEGkdidW5WTHsEVE59SiJ8BeuBhshdxGQu8k
i0+e+tRUTG1kwSMayDS1lIsPu3cYcvoMxLhVY5zH4TK2DuQ6xzVEu6PmIGk/h7WFKA4PCFzjK7GY
bwxgVXgpsWxceTk3CAGLVp2Ba9DzCqkmaz2tLQm/Kj96Q80BsGYcyITJkzBtL8AD2AgF1ZfrBC72
VOO/UT/nl1eDsvSn5QEneFohhgQiyOYTJufmp9HC667bB5d5D4Oq/Ljb0PeKKEVNJsG6bS9IDMFQ
/lI+PEnj8GcF4YvR6mDYVi4Asz/2Sqv91XW8iDsy1EE2aRayhGhiUKQ90lXg/W43218ZI1dX6hDC
o5cv65DZL9qz4vTiBOm53u+zfr5kjF3fcB8cCJGatO3g0KQ71hAhgkZpEszsPuMy7FPyG14h2GxN
ei61L1grWBSU2O7ozsddtcIpWhe49N2xN5MpQO6NT1zCXXx6O/7AGMguvWjbKDyKPMHLzC8wkWUr
3DanMrYN1UsTTW9p3q5K6V8Y9PpjCFSc7KLrWcRZluI2qrF7sLNHY3wIzCabEoKltQlpG+E3ZfEK
LsoJlBKSkPAlOrX4KpoyN7SdLEpGjI1uF4lg58Uq0XyxbtMoTTi0mftb7vHLeWB/Y9ufLy9P33UH
A93495ZnERQFG5myOp0auPcZvT7P1KWMFAVdrC2wuAFmyOIMxEg9p/8Asd2xYBd7aRJNdgwMixGE
htVEBra6YEmvsYw9rFAz6KThI3FmUz8lK8Hq51bNWj3Y8OEF8g6wodjmZU4+4DcyZvKuU0VHUb6L
4xUCsISqJpexGx56Izd7pHdpssEQWSvls6vDcsfMGhfpLjR+Wob2J/aYkiSgbuSCj8bXf0eSFttL
JI20qqe5J3Dyl+uCJ6MM3TTx5ra1S9v7rJ1M5dRDllBSTIxPw2XnYhFJujM9d9h2xrouSFzbffiq
jRoiXIGs49IDjAfT9ogOifAD55PY1WhnRUMO97s/Qs+29t3dQfaDYb19tyQiVAC9cKHPN+c9U/ae
aRKxBeN4WPeYKA/kGsjiO7LI8rzbwLg60gMc8yuH0fomKIS5vSIxay8qb32sgNfiNtSxZMNNZ4nW
JPIyhXF4qkCP0ltQphB9J6HPIkEECpLpG0dRWGlUPPnP+GRCXCCyM6mOf07x0Q7LudTOO9ixtwHz
209Jk6/A29WckKMhLU3uAqHz2pjuXsiUY3zm/yXerULl5EIovSVqhXtpfb6UhYefNclxlx32GfOR
iqUeyiTBgb7+M5hgD4dE1KNKjMrHu+N5FjfZ1DC4T1KiXmift9Yb1f01gx89ZTXQaa75T/oXSq/C
3Nak7i19eORYnMU/wqG1X7ubsB0yYcgrmf6AAA2BF6wJ/3p8GT02TL7S8PM/WSWuFs59Ifk+z+Kw
H8Nzm4QgU+cEs0bqNZN4JD6CUN92l3R9w6ZiMlW9BiRhUaelnaohs5hUo0jRzwYV6rxh8dSDbvjl
V6qZusFyRsfxBDuvWrgTBcajmMB14BY96dxlaGmWSwdCYccmlk30FoVhmGjGMkzsqvLjn4eVPCcE
GksCMGkFGxP/26YLQCwUM78268wz9uaztWlMlK3mtc4vxPp4RSvR44+nURBZ2CxU8KwHh8d/EVwM
SjA7xnnvptt8+jGLWiZs2IIkevmiJVQhvi8HtB2q4mMItCzkDyCoMZMBmOeGEooXhWWHjsOOEk3Z
YN0l2AQ2KhyrdQnBKzrG/o2pDeYcVg+Pm1thM8nvs1+yc+9vMURkwkg3hQX5KuQKQqBr5toSvaxY
NJP8aJF0rxMZule1zrE6N1MxYkzuN8gbVhUnjxH9Erokj2VyQ5H4BgU4WuqnPGp9pYFxB+olv2/y
/iyO2Pl483+4hfdRQY8wQsgQ5l7X2MeVqlEsbmNsDSiib4VnBvYw8oBwkfAxZp20luVu/lYFclS3
9TqF/CNkl39xnzGRWsUG9gUhwyLx1RTnOQw8ZjywrJ59e1qyONsNTaknWKq7FirZTQ/12eqT/Vg4
Vrh2yjedYtGbLAwPE2EKGNBfj5XrrbTtqOkhhSO4eGMaWICG275V3sNxlATetsbDosEbHLDTXTOP
y/4NTRU8jpxIWcRU94uiaBEwyH3NQLzxXvRDQQFYIzWJibffunw0quYp7Hb4pQhtbPpXDi7hnRiW
CTofMOz7xcZNXiCN6FwmEjDrSqabklz1jHMzNh93fKC3L/zbNj+cB4l7VPK3PvBAAz+oGgLIt6pQ
2rW4+aBG7WrmAuUHB3iNIGL6PruXzTW1m4SZ4T1iiZdoId1E1sOiAn7tXLk0IwZcPv/CS2NUJKKq
b8PWDGTzeHLyFmtZlxC0nSk1DSQ6FhEHgrLKU8eV4ONQkoo1SwP0zk9s8Pp9yeS9VQCpxOmPk6Y9
cUJVP7eeCi6PkSH/d7ATnvl3oQcG8IVrr9Jmdc/wnEtBGSNzNiyXK6fkh5Rfs/CUpWejkyYnLy0x
CFQ68bgHJVa2R5Xx2iNB4MxIsQQQ+F4JpcHgTP4menbhGJHfDM+tvmUohaCaoMBfceENH3k7CPM+
QPkC4Te3c0UHFRVI9F80gpB/gED/2hFH7YjGorJeHWcgAFfmugIn6BQhW53mPTWjCPvWPaAMvlhO
xtwrMLmKweaWudX6jIdU/fiJqVv7dEaWked+8fsrswYqSZuLayvjHeKsTMKOzoqLO+XM9DEmcMb/
NxbEnlP2JfW4KtI7ECZpqb/2Oa30hPTMCKA6QWESngRSN/gZJcQZEboIZDJ2eMwhBzaWXsAUCviT
VWDetSyZV/2QeMWIS91L0UYmh1Jij7PVI286R9ulfA2SCfUZMHIH/WBQKApxeomzLmEMDPiepg/s
6LG3XPsQCsEQjYbTVfE3xQV89NHFvs4Zqj8q+31RTw4NPFwKzkQadUPIfJ1T2xlRqonDQCROsbCr
azpOoydqRSIg86dz9bjqO/6vnOZymcmA6XMkt+XX/N4bK5q+jmlRakFn4n37Tm4T64WjvAsxgZO4
nQtBNF93eMvX6itQj1lzTP9QvP3ccOREgQZjlGlmZSey50TxbRb+KyFVdLVnpMdroL5ecp5kmDQ+
X+1JMAMTCinBMgG0VSGJe1CuXxgjlZNbhRi8srZ5St626G2k/pZNGN+1NfnTnNJ2siR5Bkp4Y3EP
mXk2rh8BRohMReA+yarCBmSktM1kzTKyRvtmXNHEDU9yrEaSvHV5X0s2IJvYU7uGSleetKeZhFs4
8mFogQEmuL6A1oer4knGEZghG0Q4vdo7nN2mvKF8px45VrSW+TGUraG3mzoPruDt9D0vI8e6yMEO
m7FE30/FEPV3PAUzQ+T3d6awSeu4XaTvMorj1UzGmQDnHu/yhcLw7JXIpkOm3wRlJ+sjmJdBd9ui
MhiypNwJ96S5rcI4vqgC4TMU/RHH7TWivpz6xOmJZjDzMKptj2rgZWJ/o2CZU9luOptM8legr1yS
26PWEZJIM1nlbwJ5cSKip5HN9Wo9tJlEifYdHmqY19WyYqVlHEUjD5FxFxFfPzPsqxcAn3cjPqm8
J2qo7OUVC0HFikxP58KFjwqi7xNTe3D1EwdTK4urHZjUs78ZPbmlLzE0+UDYNymBb28NXOPW5Ydt
PP0sXxX455uILO4QygGv28EyZ9mBdR+gDNRmAGaIEwTHKqi5RmjV1sJiRBulLXEpfd8NIjDXpv9z
Lg6pS3Hf2T05Pvh4kxwXZRKRKIyXoRzQuBImqr0ard+hIVNnsK4f8H42uWOL8juDBHhr9VUWbKgv
uQ1Zt5s30Ns1rpIGg9ukRwLWZEvR7VnW/Fv7VLztoWpcUYfZGnlyCCCgDHdDN/aaX7C/MS7uUaO8
ETWsx3lMymP+/T7OpPrp4TavHp0bXqk64j2w+9m3aEyodkbjzPrJA34rUciCrAPLGfJjRx0weAr4
UtQG5B9ONZgPTdMUbXm/ObWhDvs7cgdSahfgv0exK3yjyWhgTXUiKFguhRpYpvmnMnnK+fj8a3PO
idUTpBsZ8tS8NA4DN5w8g0PrMWFPb762VRx5RQm5WLndtcZ3wtAXBqefyDrZqJLbAhzoakfHygBp
zzs8DC/eohyIjK9TXeg7wtBWlEJ7IHLlRcJdbpOFo948/DWYSMmEJJ6SFMrf6OjGEgFLaUWmH1gC
w8yvL3s1RBUOC+XA2XeQ95EbgInhH+WMn7Hu0mZLgpaSlHJKHrFLGrpSxORT6JKJXLEMkuHPmrqA
z3IQlPQwrwabfo9AtG2JSWrvVOct0dx6txI+PSIXi3G/bTSTCCPZ9YAe2Peb3E/nulNLA3v2scAW
QPQbXch1t5tHvtsjkigTUDqTG4pfINRdndNRcmT4wEGv2+D24eLWqnyWEsDXUnG10Zo62g7z0xf2
qTt7bcStj1gZ6FvVTI2OOObUHejg8toM/9rsv3+qlpVM7JNeydd3gLAfzWvVHlW1TiRCXVAxoFYL
CcHSrelBePwI3tQj7yiEJYzhfoLPppdQX4ebSe/bt2Z9/emDLlyzXJvF/v99RaF77UM5mIuJyk4v
ONWSZ2/7fYDRgX3hiD3s7JNNEaGu2mJevqpkWEi3WU9wr9UT2S+QSi2DY3vVz967yG3T6G6CAAIY
A4CTpuVGd3916F+QZtE3ET+fhHlM3zNJ50kNs6LbdTZFf9KHwlYQ4MLK0JIo+F9oy0szef4YbC3Q
DhcluQpMB9uMPFU7mWxP9SvrJVx3UD6FMpICQ6UYbon4osUAWhXA5nwcyrv+0yxkWJd0wsdG3MUh
UDJRirLt26phyHUzH5sZ8r6sdARe1SCW6WidKQKinFs5+ANAhZbYAnz7eE2JRf+/FG/QXNKr1h30
JKpR7RgFgJ/kJ2U1yKVgEVcQOsNFpzSZPdy4CFSY1MMeYxz3co2DGduyQXFHk1ERYQCzYX03NvpO
WvHbFdED+0vp9/ba4olLq4IamCof3zenLg/rUMpeoa4qCj7xdZjgXj9NfpXhmMqTnRE/cZ2i/73E
rZ36T0+6/qFaFePAp4iBAAaCyoJGhqkndnL71oJNhRquvKTsJnJ77/U2EWcHxuda6RQZDmenc5NE
7WkaqCErbLEdqRmjlCUDJ/R0Xuz3a3csvGUx/ztpX2WwvBTi2Y02M0o61R0zFLuPAZPv0UrvNlgl
vVo/46eJWyLMOITsA14GpUImlmytDSMv6p0PuOeTnqmaFBECZ0SkHvzddq71SomMf1pwURSUPk6+
e1917APdmcME4dKOLU8mR3Kdjw9WL7PAodfbgPPBVX15AHcxPCEvnMt6CcpXGsxtizKdip9DgSzC
gLclwqreQWl03fXI9qO75R7heQrnPQuh2lTowgQKzXPyD33X68mhrK4+F0j/kviYD8XzwMBt640K
hvoDAYaNK+CZ3TOxSCSIPhCPSpeDxvvq8C68PFGvb4bxzA0jcm4VhGcTuLbJrbx/fNTwq/QYpv8H
41Eh/8SjcdavGyxFSPVXNB6O1/Aa3aFP0uEL5uBqtoiBnEEcj/Tx3qZeb65gPSMkmaEIZiAJV/Dx
aVcGr7Dvd0wxzXFXJ5fv06wsyf9wlsL+rmsYIGPZkAXhP1L6Xbqb/v36uHn9MRQ/Tnmd5tPo0B58
xY4rPiCAzsSbCZHGcNowNWjoEDEzIXVV8P/tKJAc4Mzny6kvOSvtk4vJX4Tstye/qrhRmkrivlGl
Bd/NsOPQNWE+3nvusYlG55F0CKDRdWb3vENICrEhPmRlC0Jo7ZLWvc3AeNFKKynOXHge4/oKqUHJ
CANcaXs+3HjcN05q1PcqH5lZQjWpNBAC7ktLZT5xNBMCDc0yic2lXbT84GLZqIxwZpZe/butcUik
OADvDz/FDCeM9RblO1MZblmBCZZr2BgqtfUKA+Fg/FaRlIYs4gifyJKm7g/5FGbJ2BBWsafUreuG
qLtMwO8Rz5BgxB7+K7HtzRPimWX3wZdJPS/OJpqo2ad/ve7fnAJiLoB4t+n2H3TdIlcL9x7bjXrz
bm9P3VHR7ykU+WkD2KkcmGj8cNbTUh6qnF/kz3ZLh2V7rTwx+46vDp17WHNNYeKOO82dMjFERUoB
5TeTqcPb8mKdVpq3MIjOk6ZDT19ttSYuo/8zzbKnc+iKh6jJ5VROaZKwHKB+9lerTR9q/i5LAfQh
FkCLHI0xqbibtE7H5RDmNr3viLi5+Pi1OCC7nE4egasvYM/DDaHqIHGfIk6zykW60nh37oQQFfbR
IOzUk1t4Q3y0sV0Z9VAykHN/Ehv+gtxIwRnMPtf8bXgFAu/DR0sXO9eEdI6TPP1axDaZPuS8TbMn
ibMzuRHEc5Fm9BnuyirSwYZOIQByWUvzrwTG/ALYh/gzpo2gKV725nkUrmHzYHiQPe07Ya+p2vtm
iBAG1Zn546xCILySfGlkFWJoI2lkG5pXWuMqk/ew3Aic3x4jDp7g4Gkrej7arENVodG6sA08ZXK1
kyls07RpogUBkDtUf6X35B2IR/vHd3eYs0c1rx3E4mBgenUSPr4DmgFqvlXGcDoxuk3CccMJFzKa
nAM1AOh3fB/bUztsizUOI5Fnfqzo8zSsavrUso3agYE1raeJ0D0eiYI2DKZ8inswQeEkkAKLuATO
KvZgMicoQqLzhhnnUwA9IOkCRxkoDbn0X9/tlj6VMilYSHFHwwkgKBNLV5iChPW5tzgYvMwjYD2U
cZJbBxTIVUMgarGo4mryxYlSd3U7XsiMTY8LijcnyuSlQpjxOqoPGpSfqOIOkzVfBcrAGt5KcH5a
osmwoKW7YIqIq05aL1ggdMaFlb7S7/e9KqLB7aby+9JeaU0ij7xk6tgLkm7C4oXEGr6+3ykn3kcq
Yna+Z9vPcljXO02jo7Bxg6riuOIQb+O1qBsK9DMZA2379nUCvqX8njUwB9qFDawQIQhwmuC/r75G
IziVt27dJueddMOrc0ozLCZS+LF4IhfuMnZxzMQWSsTGN8SztxFtpkMBbG9w0hkXMW9vgS0izyMO
kFZOCHlUQ2tQvQ1fpflZSuHnY5KHe8jTw05fiNXJyta0SaQpm42KP14p8uEpdM60PoN5zWn67Ne/
JUHuzGBqkvFQ0weD8RCUE2AeUeaETZ1m6jqE3Xlq4NCHa/q1Ifgaki0CEwWtFSEOXyoO0O95iykF
GCb/StN71IKr3fXUYZ4SVV/jg3wCHo0OYl1aWcUO41FlolheLCah3n7gqSG18i2dhPfpcS99gLNm
Zl5ELJ4yHA5DpUqPg9X8PoVt/s0deCRLPhLs+1PJfFj3Q8pzjVg6kzigSMYPkxL4FPgFKWbenMDl
C+cjPJQ5+t6lY1yxfYHdYvKAij0nWddy5x3hWwLqC3CjhUe/XvqzfxZF8gPGA9wGPwNYQAp4cX+h
Fs7aQEQZyRrt0MJ+qjeNkw7Qw/YRR9sW6stdyiTFkJ5dAsxyAFqKclHJFPC3O1kIsJvDQwV9TPZA
4SLHGZb3LsFoJNX0PKhXPZS6r9la/1/mj3p58c23uQYVH5qms6jRX+MPjLjh+BBj/+0CI1oIo8kr
YK9xt7V4zg7Kp9SEsO7adok/JRxdX5tsR365RH0xmc35TBn941ojw0hP10BRZHzUNNuVpLxtaqtc
06rEbDwuBIISyp4zVjdWOtVe7xdzaOi9+BmP4rLr8Zimicq212AO9C1wRmLu+LCYY6Sa19L5oGYX
g1FE6kJXsrwpWxNZA90q1Xz0IqxLkVI+CUNMPSTcpbyPg1at7tfE9yQ512SrklSgiuZ+JJxND/e/
2SDNXjKprfq20WSooJ9omPSsyW7opgKPb7jNbpDHPoAVdmUPOWZe1iv9v36SVdmpS1mYs4SGfomF
AUINjWoEHTou1BmSmI/AVEW+RJNykmvjxBLpkGw4ut5hiNf1Kv9RAZdagj6yd2/tKkwLhgkLosT+
PukuvxPQO9vt20BhQD0lzaGOhwQg2HFNH1Z6KBA1kwwGemajRnOvrH6MKwoQDaQhqeIwtviSKMgP
C+jPHidc9qFo3HtTJPT/LrxO82u2DnbrW57sGY1vWc+SeTj42/5Z4L6gm18NsFn3Dy4EY3y3Nt02
xx1GszdqY4JlkhQpWth9CKFc7bMKrqYTZGAhC4Q/uZbth5dk1WFy1sx7xoBPuml2o2MZQqNLZphG
sXaUc49ATjZdQ7A4Nx1lEBC0zsPqVGb+e3twgwZscqTzsSPF9xtQDlqrB1anPuzpAHCDNyAiW7xY
2r5h3ppuWI/qbsnFX8bmtwt6rvtHoYsZ2rFPKTVFfbtJjHYcZBN6SZKMDQ+1quq/6F22HM2uGAYv
3CQly/POmF3pox+MWTd7QIn9devCL1+izaSXHl8+NDr3yKg9OnTSbmaI0R4s6mdveH0sWmUX2ecd
aB+N3r3GbIvmhiVLvfSzmIgiQOh35fu6OdE6LFLMxPn0skthHLmxmymk0xA6YR9Vn6AALgOiTKY7
SBOXkCVoKxcdWbt++YX1dE5ayLScXvfPRNttgCLoZzaYHVQnObDigT2BzbJQCd8d7my2pXp4rzb4
cd7hqhcmYFs/NPXc8/YS9ubqSxQElaqTQtHkyVqIWCTf0D0hr5HaDRtPBpeM+3mBworlkZgqT50C
ewHY+LU6Dvy8tWN0fgh0/3YKR7hgfwzPuklDq45gfsiNTEuAV1HaEpBRcJdHT5L4rD3pynZpvoug
GJjiT/lGyPb8QiPN9PI6PfcHp7UiLUFLJDUdieTB+JU2K1lXVB+2Pvbw6NdFpjvl6lkynlq0SVMI
neO7fL4xnajr0HLvmtv7Y5why/oLprSf5ZB/FrAXmsq0vSB5cCo/7rk0OS+Ehzxn0lKjM/ogeivG
UuxfMCJ4+o2qdtMQVrlynERYZ3DUBJM+qgaNOZIQLfGTebwdO1G5PnoH8xYyXIlcI0ZpPZiJ8ZsC
P/l5bWUilpbOtKq/gpe4ojIEI1e/0IueGMwesrluMYyMYbu0IPlRItOeM49lokeOwjx08HHco3Ir
oi7QlbODK2rFWuhixSVZi3fIF+ZA21efZEK3YEslUKhcedZkVlrM0VeWRwJtcxAOSBoxNlI38HTY
5T48dIUZGBaAZxBLGsOssfH1/4AOHj0lu7stoq9vP310K+VqVqLWEl2fqfkxIptVUisAvrMxeLfZ
7dm1iddh/REfA4n4N7JqzakRiIilZNK9eW+aP+4HV0iJZB3QDzwzvEwhHGfTJ6mhe9xc5PZhy9Ul
orXAw1aYLum+dArjL2d1ylE/rxwKXIqYqcONxfNF1CaMkM3FFcrlHGaBUjCmXe5Swfrk40xigbpm
5+vOFNkwgk/iIxQm43U9Arkx9FIJGm5MbvL43LcSvHK+Te6XoJCywVACBMQNL9zTizkPJw6O5pih
2B4xCfh5b8sFrAs1MZEpIurrSV04mYvChn1YB588giRNim5hmJYnYhneIdW0LWwwJcmXB512h1t8
zJCgQuGhDGrPwgNX/qo33G8GMV22vUxtWdaSpLU0ceb80PBBRJ4AymQhhXgFxXG9XoMqL+7K3ZJt
jEV+BOkJtcItB92WGM3ae5hWbhkeFvWWXDy1R4vR23gktQ4E9RsD1aL9bsMtuyPK/tJGkXfkA748
wcdph5aAM+3kPU5wteObeRArruq1SkUPkj96t2gUOQFTnb8GRV8U2ojP8l6PeItafZPFArB5KULd
eLP0hTgy9F0aOEM/ApM+SKehmro8W/1fiuxD+F++JHbpaNe8wb94GSggDi6hxAw+voYyYrxxCqOD
0ABKqSD2r24Kfac4BxvsPUFrz3fspeZqU5QAYSoOFUtYOzKXyNTIxpjcv8ybqkzcG3DS9Hdj/ajH
nhwZiGo+AyjlgbJEcR77JBOjPJ0usrxHNN9qyAIAieuabrZEbub9Y9t2/W2XgH/oETO7Q/lAkD6u
UA3MWbvxg5XotssrwgWTf5siRJvSI2Vz74xdcQbMmixFHecFldAL51+foY+dI7UwPY2lz2YXliLw
whAD4EgailELdnZS1EUMLbr6WaMrjB8kAvV/YpMaT1y4NGzYxAkoBVq/TSwLIIY884ZnxtqQVDnU
E3LHVPuPcLpXcQlbAe6O7ZtG4knTjGD5URs9ntoqiZ3drxG5wvWOzGcCQYv5jzpq9RP2hmUTmoVb
BrOaUkcTbPrTt3GCy/0j+/Vtokh3pOkA0FQUjClLrqS2mdhyVq0dMZydEgFC7vcD8zK1GgjnDK7e
qv1DHY2rVG3NleH/m+RP+iLzKWdurBfgLVndQbGoT81QXo++TBwORjVlRSXT3BfMbY2WP9yKQK1/
xkWsowWsqfJC9pab/qEsM4XJXVQ9P7vmfP+HaFe0nYQhaNdfIsVJor0/YqYxUCXvmAuyT7FmflnQ
Qvk080Da5YbDMNLoPKv+fT+5dDPW9kdxFzfE6AtgOI0Y682EExKCLy9kO3IaN1wyxWkz2CQzi+VF
8sBgT/QC8jvuqq1ocPAtI38wU1OENxBYjPMWTEvIdcigzID1swE+xRKLm9jL9F+4erzSBF3GKE4W
fwWRW7SItywE3jGrBz8NfoKj5e78UIIPM3tUJ71uGl/1FHTu9wFtHbHjCLS2DPP/+jO6M1H5kygr
ym/QKS/w+gQ+Us2xAR8PvwvMHWgard5cZk7wQ62y2JfGggu6Z4Y+u5d5/AG3nayohMOsFkTYhiGe
tu6PMVVut+bDAa7trKiRZqywkmuQcSsoJbKDZCI98Nd23ltaajIG5XvnuKNMj3ISGKTShcYPjjML
uMeCyKRQm3VlVgl9HThUu9WJPBtW67scB0pLNy4K0lxBvSpiiCs2HPqagCb2Q31OTUDcr9a385U+
Tan4+ETKmxE/GA2hf5Gq0yVcMTiZVHASQ+09/SYZ6aqHnHr9TfzfICXF/zp2oyNbaNRsarfj5JcN
9uXs6tR+IL6zzjeaJyZSOEFSwpNPjfTHFf7gpuzS89TpZjgblAxvB6BLNxNZiNe0ttbM9lscsnbs
FTDDwOwzfpe0zI10JD2FabvsB+Lqg+C8y1cyxHe9zF3QGZyrdMuBYdw4ERSaO57EG137QHpyLIud
AmcLdoK0KtpA8cObTfEKdNjl338bjjCzPEKoC8K70UP3c8nW2gDSnLEzXRPuszQLk1Ia6kp5I7Kc
wP+HGcLgiGW2c/lBXNP0dn4RwTa/rwsDX40tyP5qumwQzUlOSsCrjMAWgNCia78VkGluanJo0tdF
WwcuYeNzGcomRTVSkmHy/VLjKjHZS0+ObWxrepvSD9TO2q/y9DL21X60xf2gkY2FD6IMji7KtE6R
3b8w1d9j9bNQMxcg7YEcliFPMmsrKOTu1jt9F1wL7smqJYCfDY32z3kWYfWKt9D9Entp0yZuA/nE
v0LtCk1e0dVLjP1ry42Tp5VP238njc6zrZB2u8Tl50uFhCxzWtDx3yzBnEFwgZwQmF4nABeM6gfi
2DbubPkeOiqlSN0RtqGHbvF9XL9ehObpTLhYWMuNeDoxCgP1ZL4qIKn8YzqP9Rq9c2UMwsq0iQ+R
4f3B+55bs681AWZaXHFlJ9AsejJyFcZcMsodJZ51l42nftWi/pAQrdTQjSK7W4y5tu26hUaxmWiv
TY6i4sWT2h/z6UECtIiIHplPKAtqUus7yGwK0kQ42aB6CS2lQTPqCRNHAUe1G3dTczrUVoTHxwoh
so7P4h3SP6dPWvD+L7a/jgzJPQkgav1t0YncWNAfzMxYEZTIB0m+qyBFNyF418oCGEgUw/gZUQxw
85w8cNsSVH1OvjS3v+8LQ/dDIEtu1e5O1ZA+9WI1qNF158R79gH1TxfpDCdz9CfUisygsNgK4Jux
rUcbb70u6luu8LHSHErvo5BtA+PylqBxrYrPn04V134XvPfabF/KQIWNDbre4+iPQxGo8gPN6Vgr
BLJlNFexbfdDDW7eoqq0vEngSNlB26X1+MHNlsEItf7QKYCMMSJUGSeyms4DgOU09sYBPtq5dP8A
w1ABB+okUqSiwnNUvwAJzq/gF5VOp/85U0uOqz2TmhTcTsITYhjdJDkbzq9lqObwziqOMhpNc69V
7UJDV03F642TRvQ/xaGQPEi1cHy5V4uLsG8nXtSktH7DaIfw/fJPNpJq0DgCSkyNhK/ygMIuTrYR
2B5Ny41LNeBemwWdUwLpEz8JHcqtzJ3k/cQospJmddtzLnxV0UB0ArddGDOmxS3gNl5IHAZsED7f
mJAFhTrQ7NZT1Dk8bvNx7ABjwQQBIwqnL55wTZ8XAmmw5RJJVOlAs6nr3bbKEaEVhGPdfNDtiTmc
XfshPJSyXZ8o2j96K/Brw3c5pJKVR+NWuSUrtoTIgQl+Opf3mr1w2iW0I+d/7n7qYk4TOvUcaZJx
JhrmwT+OtuWLQsgIfFBXeC/2MUk97PLkkY2tmTUvoijLXYcG88FGnd5VEVZwz7E7Hk2ki6UTyZe7
zGQ8swJM18k9SKr8LBLig/Aq+XmuxOx1n78ZgO3jI2Y+Ed1kn9/0Lbv+IiPwZ+C17FP4z+hsz1TY
SJEv8zuNpiaGdKTtYWREzUVmxF55VDJZOR1z8MMgXIGzu2Wms6jyYWBP1vd1hpPLXud2LaAsUP+9
cbZxWnrr840n/EsH8G9485UF2B0vKTAx5vMwnNquiW74oAxP4di0brO+bI6aDj61p12dSSAc0Do9
HxAkAwUCHEfmyXvuUnwsl3Z4zcCxdi+hue9eA+9NPgyuhq82kLCWMMFP+cVTSn0SIF3TI27VHrgD
1W0xQWsrj7pbF7eCnfiPpYbb6PWlCJlD8rJt2gmGISvLF7BtcAUYJGAn21naC3zYBRF0hIiQ/M+g
TQD8e2hsR/ORGzxxfwTca6evj54qYElWihdIzA9bXy9RhNHysN6JV5S5gpYrGEDfYk/XA4gyn7ms
vuE4phhd7oRXbJJFtjqXVrTg+sCQOt39AQkVGLolBUT/PQBS0HA4oCbqvPZSITuxM6mkGb/NsrPS
j3bhRyzoK+0rclkNobz0uNVMN6mOHLSWq8fQkDK/HSRj9wOG6ilN9NfvEl1DnhE9p9VXSlzk2qit
PV3bv84odO2u/pmAXXjxKXYCl1/y+tjB7PynbkkCLzqH+6qCaOYLXUB6b8Z3zEtvUbsMNtPcF5Sw
OpJ2d8xnBfjflgj97ipe60y+w8XRMrTh+qQ/uegJ/rGcjRt/eAm6cBZkWh6RWZM2OWV/bv2w0i8P
7N17f4A0SgnPiy41Os0qFu3VyLisQc8UHGudT2HGDsNRv7O700pCaPXMGM/otjS5RcnR0FCZqLQx
gN0mQGSnx3FAHiiz6AM4URTP0fDwDDx9NpXrBfAl5lEgAvvMUXmUki/q2rQ8XvU0sLL1y7ShR57o
ukeNXAQjYZkMIXhVyNHJE4DX7yk6mVhDTYsRYcbcLYRiHo8Wx3erm3pv/+1iG9avlE04LVff4wU4
u/rP7EDnYmT/6UghUVHg2XVU2+X3m1mdQMKvG7DbRcdrN/Yep8oaRhTvULl0l8fAbtEtMh5dzQ/2
VUH+m4GjIrj2/IVgDxbxp62MKBroVLE9bRA72HIvxhSqA3U7RxvSVC6sa703W41B6f78T8ouG8WR
NtB+n0MwjKRd7cuzQI4Gp5DuDnmXeozPkk7TGS4wjQzyfzkJXkRPjuDHp09+kSp/e4B1qdd38oO0
p9pkpFKdnAF/dCdJuSJvq3wJ90wMC0q07v73dhCTcD38etNHbdzrkCJLovHjV5XnJGibNk+ARZWT
IOJDjW0l2JSvLSfYTWOm7jBtbTYfQGKu4ta0fzXVykrvanfolN2EnBUCOkCqf6Iy3EXDVBuyjdSY
A8cYY2JOMGg4YHsa5MSkdVL5/LjRSAOlP3awMzAFgJI8is9qf7vD1ICbQm42zUSJyQw3UhzuDNCI
dmFzHhj370KwhLHE6w1drhfRO4cCdQZW8p0wOLtiLrRmajqxI0Xc68q5MiPuc4swSrUZI3WTjEVn
rROju0Ybr/IhyW2CirjWTSC0J+bIZf8BygQZW7X7hFgyqlivko2L/qs1EmNFTGKOfg25Jb9Qs6q2
0vs3YPuemxjO+fUTndrG2w8cxAOLN47WA8uBXAJh23eIan3tA4CmCFYL3uX6iTNe70/RVsVyHCb/
3P7kd/xOEHhnga3DT5izIo0bciorAAhnbQQ++mCc4ttbtqYjL0L0/qLvmMWL3UVHIf4AsEuZX8HW
V5TYaaCWRwr3VMG8yDhU9ubNeXO9f3lvXnahKYqvj+i0RFML1VZIH72Cc34pBLclKcEcprHUbBh7
t/+GiivLdrkqLhmjkR6fciORvE5ben9Dy5hS3VYcBK3TFsE23EDz0msJIMTma56+Mjw0Dx02bWXX
lPembBwT3hcxOwyNcDano1tiVBCoWrt6aUxabiu8pmrPZ1FGuXNwtKPLaXeNIJebxFTCyDTtJmeF
qyML92IgrzFN8WPAMYu5MNmlhBAxJgCs6fAOxvkwYvwO7Es3g8Zdu42IJ0Mx1O8LWVYFiGHnJFl+
buanX0+AN37bmFlGl17EUp8C5FHeBA1XBPz6XzIp1TicbNqLJC6HRWSCSrCguFyCgafsofCgikpc
Cc01m8kl6IAnhjvmygToM9QVdPSajxKCTMrgQnXPkv+AzPo66DiDbXaZ4EUSHqzzkH/+pDtz1jha
cBH6gURLAc5mV2XHqf3O7yF2vk0sog0xKQMK6RrEo4M33FxSxW6PgILW4lISxuc5lp8Tlz+Z3RXi
Lx0CaF6K2lFnWIEaJIN8F8kA+sMLGFpRuaUXCtfSp2bTCnsdSAUSylDw4RcyordQ7OdsIYhV3e7m
WoH0MNtOcWXxi1HKpQ8cqgj5UaCowLSmh3/O45n185ed3U0gdbbG4MbfTfTK9Z0qpXtdi1fjjY1c
NNztzYnv5JGhlZn9CSitqInM5o3/WKHvGNX0F3px+IISN97OMGA3kJZinj9N1segk+6WE771TMCz
8102r+6LQS7+JyH1HTyYnCBrXUCuovRqq9712+vK9ksU/efcNQh1n2rGrcnvk4cHcpHTn46Bfd/x
EeaybxT1/sTdyeIrZPGCXcp7xRYmeqt0GChlZna50T3rZ4z5Nf5bhKBqpZe5/rqmd2JmkKeMydLY
PILMgFPm4kvpI1uqcxhK5Afy/UBuEZwJ9Mwc7zD7+9cOAaev5sGen0wyoSrA+Y3LjudE33jp8QNF
UGkwAFrV+bdw++pb0G71cXCtv6cLC6PTSBN8UV+xWaJjRIYxH6F/z1dQtre5yo5djBXuoV4/CMUb
UQBYWKdMT9GmUdap3MXs4giq55cdAYSCSljyqt0BoeHnfVaPKbSNcF01YCi02hrrYvmWLaK2qPWb
BnRpcDA6CiyNfMqU5nk1Wbj+2DNX1NUVev7S8tIUqqBFTA4EM2i/l4GcImreLC3Zw/vKvhzY2mXH
yBzrJLLnHM2zMcYNwzY/cIilzPCjG6RpG1CPY+neZXOc/UOhDpp3rHEVqKZ4pvJit2VaMqNYrNLU
Px6/wVS1oXkMtyZRmw7hh2RSWQDXwtUNymVLEU35kKnsLClumYJtDREaXONrcY0P7BbUKufKkvc/
7TAqau1Pn2jBm/rBe4OBdgjq6QaVXdHOBnACqFRI3JY0fLTyehgyzzzUEsCNQl+uJNXXB6AGr2bC
LitQi9okdaAZCBO4+vBRfze5EqjR12krcXPpta1/dnqYElg7SF24FuD1nisxbiOSZLUdtrh45hUD
0/yqYF5l3aKdrpMPJSRDwvbXZvjW+b+UzFPEmBAI4MLTwryO2/rWOra4TBOEKLkI0R2otWLyOFUi
0oRCbIT6uEMjBOlffkRjKPrZgd4sA8xkUoyZdw1/AlvJ+H2VquVGmEZQqY8U1M8f6l2lwhTIEfp1
hvEhCx7O0D93s7HML26aFQPRI2DlinLyRN1XbCZF0YVxp2HKn/NZv4XyPM9k5YbfrGGY62syUGbB
hk3LdWCuOZKzi8nk3Am52F4Tp+RBVJG4c8TEkCbQK7UIlntwrirAnha6dLNP2sqPVk8OHcN5YyGq
1eyUXtEuXww8treZuguCejHa199V4RSTLdXzKKG2vmjWVdctAiuttk1XHdqmHP9KF4vPGEVMOOhd
yP6/m/OVRHL6f8kJpgDaf1kb4zx4S7HN4DnDwex8w7vguvhF2USDjZFnJMyuehpcd1B3Ur3rT1+a
SSpW42HB9tfFjrJHxZWTUcASoYm90CJKdjy3NRnubB9G9sKfzQkMZEP47ow/dNdAF8ESx3pht6t5
TiFq27huTGavfOtNMfBzQkgKLkDcJr4IrDoXmk67PoTFlY+HPudjYw45eScHYmeBcGAqWoY59iE7
qVanRn2AP6pW3bE2cikOLPzv+in90zbRJCc0plA7wELonjMZ46ngIBhsy1ggPrI/ve4hYgH5vcZA
2VehV00gZYvfDwdvoLokXD0jPEXuWUlMEPuwLhAJFBqof+mWs/rTzxeERLdd1YoTVth0m9kqUNgR
50lqGE3yKGIHYSXXOGy2qbVMxeRaudhC2LsKp6l4w5bWII28t2s7mc6ZeNfKLbCWgEVMnpzawL/p
dStyLvKZY1AjM2dYvOb5Gy+mVF+RvPfhEABObeeN5yKO4dL73Nz6h9jMk6L8wwm9HVDcZJok+YNh
vUAQP6PiR6GL8cx2xH/0zP7lLC3h8wAlTC+jaxQrQOntHvwmow5jMFC3LgDMBhjweJ/D4LFmHYDp
F9cU1ygMmubtRcUkwtRrjRR7XeHHWXvXCBC1+BVGIjm5Sgw3wsc3lN1X246WCpfYQ/EzifIAA2Gx
MN5towkGsRFYEobMyuncH+wzueld+YEenUmXHOlVcWM13TtnQsq5uHjrLlG1VeswoCQzbg6XgIWo
xn2Xc6SwjUj4BppAIpRMVSJr6hTkNM5Ip985VrdJqBZ1nQGqtzLHls1hY3PlL2+TWOSyKYIeWWpo
hzUKoJUYEXqHN8lskc9/gPV0pcuPjXHQvZfvYto2vi93da97SzxuscmOzcNzboi2hNI85Ms/6Aoz
fsaJrt1DLSvJiJbMhGX78ngpA2ku9Rda68tl8cVqRNVFp/4/09/qqUXOY7vZHVmUJvP2SwZdQMxN
Dat7gtFTiX+qV3Ar4U9DLlo3FZYEjxIjBW2vc8YgmhoTNZzdGQBFuLPR5yrLJkrnJCAFpH02c9cs
Br8E/HpA0j6c6Q2JiyIVZvyW0gqhn8kUgRu2FnRsarkOIU3bIcO+jYIgqGgk7DDjS9yEYivYwPk3
f0P06K+ooH4uRgzgXQ9vu/BQ3ktccgOTroN7L4edkgjwLQd4cIMs/prcH++txatzwJUPgWe70AOH
r3ZDXuUwZqruXQarU8UbdQRw0jvX5S+N9+fioh8W1AM9rz+1vKYYRWdqke/yJPCEcK8HLf6vxHYm
7SETbNFiOT3l6C7esKoUjXxZHvOcrcW+eqYRawMYDcug+VtnOY+fm2ELxmoK+C9GzWOLuRQDO+lT
rZLnQdvqljwhLCrcyR7rTTJnjNNcXqTFx0rlfi6MC2FadIb5Mdb10QPRoyNID9l0aYn2PpqQGzVc
YcJaON3J4PvhkxMuOcSu3wJgfglElA1iEqm9Ke9RfFL+HWVFBvC8cb3ybjD0pHmf31BtaRymmtuF
jfzNMbyBdXZNQmsLZth6yj9dSpY3TWolRndlZlyUCQMv9x5FNVkozadVwHTxpe51DetgyMR4pUAJ
YBiWe4oLelKUYNPojMh+Qcx8JaHZLHpTPBCE2pbweoDblmBXS7MBuN9sTJjk/15dA0CFVOUfXXeU
qzf+1ns1Q1Fye7OIuscOqUezK8vy8o5dTS31pCTxpNskxNqMnSwgyxGE5H3Yu1c7DXd9Mpq+gNYc
5NSyEuE2/pcTrSbjyG+xwUPIli/KKcLvOX2iF2GzaHkDXhKp4QaWmgqq2FzFrb/SF8ZIaOmZtBRm
Y7T9zyKGV0/qMv3AC4pS9mY//0hlI6vvPnNXKJ/OcMtX02DWAH6Rv9rw2Zyx6cR0+ohqeW+Xd2d2
T3w593BkYR5gqvK51xJKhIbhVRDOvVDM5P+QWAGtWF1wkTuGywV5MSkEcUD739SXbYgFPgVWy9vt
guehQAHj8qPu9QThEjedkdi0BNVH03t+9oKiVutodPO2A1uQH2yO8ISQmp+rTWXugAuCEavi/fxa
ryAjK386/idjVT5/ZeWswcMgA8E3LKN0cRUJp2KwSNmdHNDEjVYvCYFajEyTNoFXNDYDviAMp6H2
fzKzyG8DqOF1n1Y2lujUGj/Ut9UOzfNKgrCeab5lynpatIoKZfpkVyQnUB3pAf584URGf2XBWzvR
Uwo/eiutyktxgW/rOc7EVyDHQLyj4qxquVNcLAtdXXG+QR/JIa7iUGek5cOp4ClOrtKkMAwp7t+X
1Wk3ct4dC9GMiQOIuNBkPEFiGO8w0vdREx7D/Ah1Gr5Kp5AJNRQXM8Wog+WOvtvG0c1XCcNkfn80
B8xNW+7eL0B9g2rHEmdcK93bRiBgaSLWWpXCI2NCrBY9/zOTlVe8Cag+vghbPu+hyOH3+mqZIMco
bw5c4LLuH6JDmcV8wQF+0CKk0mHXiayIWrvwRGs7l4lcM57BxFz15YJE25pY1dBo51NzyNQc+qIV
wbCOK37GeaLKrTmmAxkSIFCb/6Q2SO77PvhpJR+DaDerGXUmtNj2U5XeQSnSR1tyKicAWuPJUNH/
w0o/NcWaWUnVeZAM3+lwqruvzWWodnn64kqYdeJfTz31E1B++LpyLQuPeKDJlqpTFx04jiq8BCm1
/qJlWrU2OyER8zMUV0P5IgafrUy/hubimmFaKJ6kGl4YWoSkXMMWPV4AphEyn5h4XiGeCbmpLjkD
crho0HwEtwX9iWmtAce9zcDjN/B6HLjSYiX9ilE1w3DPBZ7sezabP8/djJnHUuie/2JGTYZz7YSJ
4w0mfmruV0QMMJOdgQHHSCbkzGiyQ2gIIW22C/buwnpgsP0oMzJqx0QFVXRF3g+0WmfWa/MCRJ6/
GOV69EBCZvWmjywG8Gnd9dbeVJr1C97UWumVt9J8q21psVSwBpoBpCdPwEpsh9b/ybarYShCXXVf
o26rnnh5cb3KjTyxBXgHbmdANTkNtARYQnGlqCQoG8E01Njd29dksIvhAmA0JIRNcoCQOJiLBSfJ
UBSFCx7zkEDwBCXsVxpXA9JBRtK1sedOS6hFGCCVUIOoLrcTSbTKwk3WcnOT/MIh2ahFIizKd5xx
a9BO9xvVIoUYXKftgkrXS2vA+1DJh1yEUGHQKjJ5JOKTGz4FS2Uy/H5/DlapkP75Ui7eepN90NyC
NCT+HLyhssPX8E72Mtgvu6wKJgaXYKp/7wf4ZC4DMKRhI8exS5zTSOxGIGFD5t7cAR3/ZhHtnagZ
HiVGa1hmGf9tcNyjeM9ZN10cEo8aaN4QdZOgiUiJFcYm8wGLCKhNB3/o/XVyZ0Qd0ihknzzODm0q
ioKH0DqpH2dlLbgBc6/kutHlET/NxYt4l8DT9Uhkg4AoDV7+WerhVyWQdQ8Ag0AM7elZEok6F8oG
ugstm/plVeAEwVN5boBoRWhM9nqIauEnywBU2Af0xrEtjgKb15ZQFeSFa1oJjtcFHDO6Q1ZpYwnx
3ijDi8qynBFVVIzvVGtYETr3XGMMxYPAca+Q0pcVox3sHj0olm6vW1WQmL1XS4s+DriSZ4VGA/RC
GNXu19U78s0xaOtSUzr6T5Xtn+lJVayjtBRMye6K9LMKcz2EllqwnyQSnd7n2j039bn/ZSqF4oQB
Ch848LXW/26hW7Ff635mbVYOgL8zeCeszis3gBT8tM+Ck1xawPC8GoijYp172BZj9B7pQsMa9NCb
0zHyyBhB9JyilSS5oOkMPtvgNnRLlYEYBg2CnqfXxje8hU2Eb114lgWKO23EdM7lhLDne9wsWz8Z
TZUE5YB/d606c2HP1L25AWIjWfDtyzdWV5D6EFYUFTVoaWzGJZLgG1oGzN5ypwjjzKSfE5ZlXZqY
O4dwCBxnU5/GsUKrnJt3Orex0YjAoA8mJZj9Y5fRlV0hNUxiagd/bQPOcgNUedtSfEA0aawsfVm5
diPXBdwc7EQ+oxayxBFCh0VL0/zJIwg8A0i6T/luFHuVueazMCgxkOcX6e/14p0vWndkSG2IZoU/
27y3ztXzKVUtCQzOQ4tUMOrjxx8+BdgykDvLOA3N/9jckX2ZXwR7PbdE926K+TfJ6N9c3FHNJh56
NpHRUVeWtLlUPGuPiYKZujEpQf7+zHOSXYCzXtAB/1BUFfPRY7nyWVIftyIgCl5eL4gUc4Edvpm8
g1e+8LyiL+d3LVbEiOxzZsB2UsccEwb/02//yDnH4B6CEIYXKc7B77LW5hoXiponJVAm0CsB1qCv
AaJLRV0+A7dDGWm34CsOcusmGqAmOST0cC4rQsvdGMO0ICEfv5024ZQd3hTxSkf8j1vdbyq1cb24
AGS9kYXMUG/VCvMbtyY8ZGiM2cjyiHjOpk07ekmVO3F4e62rRQ/p4OFmTRepv6eW17CqIMgR5dPi
kVYZmMXLtiyYmDkETafEPspfMvLD5KI4XsGvOU25C+bc1MZHWaiY50ANgSHMmDWsfAcgn3u3zSn1
K6X7pbD+UDAKB4+qQrhYZPYx5cAGAVnEeiitUEkJsUR1XUFDICujJ3xpDj9NlPKw6CcHb0CKTra1
gqgjPPcL0VzEQB4S//KyP2uHhGV69dR8ZPywQM2xiqpPA0rwKXCweMlLYUJKOsioEQvJd/lJM/ES
W+uTzlRlBD+1ZTdCFj7DTWfdUrMMlyt1B854hJSL5QdML1m+kYZaonxe4h+g4PUf9VhK/L0BM1Qt
JtZPv3KSuJRP+7R/BCL8EMNTCFrf4zOR7xYdYf91V8eI5eY/o/9tM51l7oxQtHSMMOWyYkQRST/2
+d/OMRVQrZBDVSPD+oUKaA23NUSIizPXcxKGmCMwYrCuG6cZ3hm3floqHt8VIpBjC1os0s/2Q2Jo
hD35q/4zT6XCzDzYGY8b49XRmGIVc3IgqSkeKJnRFdlg1zt3Ua6yGcif9iKCDc5lBui3XmrpJdNp
UxFurMbtK3V64DoASZrvjoLtzzmK6RP1sja8wtwIGidu+FDTLHGuZ76nyOXJLs5homRSv6pj8WCd
zsjWctVZm1I8Xv3doiBCnebVPpyhmD8+VFfaHclo0XCky9Qg/JTXLJrlnbieEn8AHmsm7AbT6FIo
SMvdHKfYZd71fHDsRcjmu4lW+iLblmTiCReFZdZrnFjnUb63Tt5Ydrx5SSFuwutU7Q/HpCCXDCnj
jqYh7hsTrbvOWX6FdOyHUITey1+crBAwBUX5ML9Scua1wVmVx0QrgGwMv9/VazVFa8xFPid7n6Pg
WZo5Y0P5Fxc9uXW5dGG9WICsTpO6TJdH7WX9Q01nNBlF13McmHV8cAkcf3mPt/+OkhVS1x7gFA58
0okJXGLJOicNwcccVHGjRkGpxLI26YfCPfh46Zp5mLP2WV0OVz7kFepYaWqne99cvU7LCntVIT2v
vw7eh689NRrQxagCh8HronoTNMrpJZ7oSCoFV7BOck3iH4W8WPZo1YcShQFLTWPWif0g4HsC+npN
qiiwkIv1MkIeWLEBxNevJVO/TiKanN/Thpcv5s1DeAK55ujw6QH8WiO2v/rUtUvuF+Q08Mtr4fUH
6OBAaXxv+XhbxFazVTmzL44B86yrcqefmj2CzfLZWHDBcnvjJB9AXszUraloP8RIOEQQTlP+w89Y
ClZnfRMHfZ23oq1UxGAEsUwUh36Jbzq8fp3Rsul3QdC2MdzWtZEK69q0lsqCxJClR1edaR2uDMkX
FDj3UF7ykTSTjnQzzP9WQSEUAns458TDuFTtOvXd/CAaIEz3Xdgl1Sbh6mA5MRSmN4A0+GtSu1tq
OEBsDGkdiB5u2JhgGlro4b35YYkzxwtsEiWrIWNGQnuFKkwfJzVs/7X5MpFgOd4sgCawl0imKNgx
B6UV7atO4SJu8jpf3EZ3idmn9OzY2iKj8EZOrOTUK+6S26Es35N504CmiYogk/Al8l5oEO0sL+yI
WNbpWlKnCy49zCqwQS5/qaoSCrvaUMtTr8ZqIKYgRm6guVPqwP3wLQbnI16k+nHE6d6Y4UegoIYr
NGn7bKaeWxEEv8FFfRjK2BzYnb437R6Msd1p4Yv/LI+ARCulQCrCg13lOCKC8I6++7y8eqd8hVd6
86Y4Oykt+ZIj7d6tY/TOwUR0S6JpxJMyZPXz8DGQaGwsTRrANGGBKbYMQhTY8Orfbixd9GPrWyad
MbSaj9El4btdktIKa77glbKQeELj/s/Zo1pa4oq/9hoKElh388lnnibDYfDZXZOUSFahtCau2yty
6eS8PFtxneWgDWtI20EXzkBN3DPGt7ufSyqpwTCMsTmPO8fARy+2sKV6FSCkTZdoEuaJQH38LPst
PagfwXCnD1izfL+/agV4YZVZgTd16m1jJ79+RbrxBt5JkbBPyQzzVMw3BPaJKN3/SQylNB+Pjz/s
qg/U+YNAT/YrOCT2zLyOM+dysrNYvegGjZX1OxHszvwzxKR/Bb3AuzZjiyALOKr8+uFAYLkpNOF+
u5QCLWZGP1hvfjoU/SFWpSlF7Ka0h1efhAypvQ6GVvjVpSTY6mItTx0hdUeT5HcAJrWFr5YDYwD3
/jqvTKh1EEjakhBfSeDkMHmUwOZFJ3VSFQRXyhz95L5ExBfEAe6amXaAfh4k0OMr1Q3958lZCyPd
Qbf3IeGqy1d4NTpiXHky6jyoW0LUQYUGb07lG2FrxDGcMRKdY3Ykmi2BWMSi4kOpybxcLKalUx8F
eepuBTnXrgLbuCh9iweeirq3LnM//d2eLnlQciau7iCVF+xqBMEDTuFn5qAuAI5LZGCB9xxRt1BU
vtwktlpRmUJAgYH9qrcWUVTQAyLk+eGTkGskiJzztTKOj3jCXMZUmbk3NEd5mXenKLy1bN9WOm7z
CmTq0t0/dNXnWIErDDOLRfl7d9ryvhOGaDe6RRznBpprPiG2qWN11UJ0kt52tqDRBGC+R8GfeVr5
X/VCNYVWt9+aRHYUbpvWihfNdf2gwPVf9/LrU9mHmwA2iULtZQCJGcr6IqhDw4MKXJ0DwvA1jFmv
+kWBwzerfE2db5v4e6tQ6KqVJ2mjqcD5fWeZLUwxGjiqZVSsUGM5Tow9udsCCyQoMHXGQIxb8GRa
45HV0P0rlUarsiDz6EqYWlUC30kXYO5UQceMDoSnfDjImH0P8c2N5rfUH0uqGEXCRMalmF8njLgQ
ctp9KTWK7aKhOEEttJipQ0hdz9FWCZr+CoYWolNoWf6XT/Lme/yy0ivoTlJhIzovHXSx5WLWmL8F
LhGeASx0jkwsoqz7+FPQ4abnM8xNPo73XcH4t3mxTADS8Z8+ZCrf92dbPsen6atfxBfxV/KMu+2a
8PWQlJJ/zkTJcBAcOX2nufotsiTXGDOI9OoHPatYtDN3c6Sx/Y+twdkQgtDmxzghbXLXDwxN4OJV
vdffQmdyAHhGO/oO5pMcJ4FKK8kZ9CFhPJ3zn7EGY9TNYf1YhsKQ2TSYUkmSvLPVyvX7QfdK+Th0
JEes1la9SnMrRZQwZd50+3I8Tp5fIPpcllo3xp+NLKGv/Awxmo+eqDcdTDII4fSLlvMdyEoZt3sP
Jnf/j66yAGLpepC1SZO9WPbapuLbZdop/Q0DPYZVASOA0oGj5CluUCEjRXo66pV8tgq5V1N1+rvL
ASG3zPeZsHUCSB42R4ElVvojoj2+q+B2sLGmNuccDDTBm43ns2r8Ryku/20suS6e9nU0VA1LWYX5
/bHsmmtHpOJo12+1nmWK+agolXiPXcfsYY2/u7y8We0+GEFL24gDkc7UhOag+x/EckRYsBZHF3O+
d4bnUFOjrOM2ZC3n2RjKtiQCrUfoH+xp+/9bDka0jZ9ppAS+D2ETpGVdUwFxbw02YYv50dWhVcF8
E9MBELmFSx+EJ4Kd/JU2H/lpgNV/EPtzvrAifDUzHDnWw9VFvy9S8LHaMBntgD8lrukazalI88JR
STQaeHG8yrL3cHJy8vGVrBuMhLz1WDuAahMunncYr6OIFmGcBd+fJ+VpAEX5iSoqggLZKc6IwyFw
Nx4eOW7u4NQe5Ikv2o7UqjD9of/DMHSGx1hASCEL4ZP/6LcnMONjjK/xLTRyj9R9XsTcm05eqQ4e
hf1VR6boz9HYHT8P7nqMex9PJi/uNCpnzSfvEWVDvymIpqW3YjDO2Z1dTA1x4yb9c5EjE2UquNAs
RH9257eFQcIOizHrqwtoLxkyJspfm1h6D+KEi54MPrjndfIkNfLtzG5Vf3/TIDAl+4eX5hdk0rqs
6lWuvT4qn04D/FnEeZF91KHJc68OUZovxyJA6yrSEW4o8tW4aZo01madhbvy8gFqM923E0Hlzyt+
rp18SDKXNbjxtlzUk6pK0isW261KNrIHEjN6bBeF6jlRWjUAscY5MZKXjrB3K2lIrP+53/sDG4+l
k+6LA4aEcwR+w4XcyevR05g0dNoDrV6jr7K7E4+VPFBSOYqc49lJYEBbf7j2tZ1JDWzE9tiPqbDL
7OD3oB7eY5XU9ZXpnTdYEuatyoMh/m5p0t+EGqOKgfac32KLc5kda9ng2/mTweInt8AAnNR5hdUu
dSK9FXUKig8laKWknS/sod6TF5786eKe40GXRCuH4zROr/qns2aGsHkCxdwtkDP7jvQIh4iGUX0D
2Mh2ns6sZ4pcrxO8LxzfbOanB3FK7VXeZETcKakKLYvaYGX/TEyeGrIy90WFOiHa/J9jQ2JTncX4
fE/QBNGKViXUh/2wGH9fKGSd1isXwr0HfGT1/MpigkISGneeKsaWSopR+2rgdON9Y2CGXhYB3FJ/
7Dl8DXaWpYIOmLkZYB6Wzx4L61YaGpjyHf/3BoIqpLHsqTj7fQe0n/ww1Z0qWFCHKzJe5TAvWLvp
4OGM+v50vax2xIvipXBgYqG2V1dvZtRVGQ6XY9jWk3b+MV1nDshOUFlMudXcmAr2C5glsCvCXjjl
INj9Nkjoez5/XGCRrwP7r2gtLJYmGFwXbRFPMH3Cy1bOzmrSfmIZ4zCpHS8W3HV9t6VYNq4ZM6DO
MfP2U0pXZMZLstVUhZ2o/XQnuoc+/MRGcDKomPURgWroNM4nCNCk1REACYfOKGbh3Nhh1s/5uVLu
B69H6jt6zaF1yXF6RmGwyLcKVMRx867Syak6iobdc+5JRx/E3CpjxmuzFnV6AmzShWu3Dm4UBKDP
NYsxu0JYulpUKqJZlOjRcHOpjQzIWPaDgh0XcsFmUxtD9IHyjyWRezQO1kSGhLKv9ljUcIGeSFpB
uqY5ufMMAol0b+C4FfLZqC0gmcdM/bTdGQDXyxr3c2E2jvTn/KQhfgS+dDih7uiKqYcpV3i27biZ
SELs0j+3Nlyr9w2SBWeC2gT7grPwQ6OLbhIn10K/RLEvGbjsIP0js6kiCveHS3wgAWmQIgB7qaGv
SbZHsvFo9yCTDjH0CFnT1Fv78rY3rjeY2fxGSsedu8p8keLfPl2Lp8k6fYOfS7owJGnAC2AWaaT4
zFoC7SdLeI6EACJTsV+DwCz+axxwPYUXBHxASKyckLWyJGVYnmuR5C7TafHzYoGUnEpTh2uI7S2b
dMbWWN3h6BCkiB+cjLyOpmDJp8BFbmobD4Wrx1sU7Ru7vp+HObrab470RIF9zODEi41fRywg9vZx
FcMLhWmCxK/DeQt2wGw0U2AoHmAOdmug1TOGeItLhGM3htkp2vTRdt3A3DC/vfaH/4JH2OzPK0hJ
+D3kakHhDZiJQRzFHNI3MxIad5x0zqspMSMZhneIGcN9wI7j2QFbGbf9HAiuIoWdrMV7aMR53XcR
EFABFTUFA5HHrb/2NpfxMbozXmZXhL8hs/l3q3uMnDgc8LIAASXVDpEugy1kABSb3isT8CI/vfHm
Zg8xLTrFN2+q6MxrmPAZXSgV8Kv//LMqtL+Q2BDP+YjlGjUuPhT5GXxVQJ0wvnEyht0+oR7123U2
3xtOXHiwr5wmMnclGxtMlS9akYncgYZ2NRViVLp+3NkrR2HtnCTA/j8cQYjQZ82Aw5c1aRsEi4fu
aYa/+/M/r+zGiupYitKlOUEo/W2lWdRbZQ1/4yXQIv4yCl+guUFcqATJaGL4eyOZSx99BrlcDd52
Un/0IyHcoNBLP85f5TW4c+uUQe97/dchQ6S2tO/V3OztJAVRr5l0ts3E8Q1yrcZqVDpizLxgsIQa
K44SoQSGTDdnBbZVJbNIE/3pV7yyYXKWmlQCvAUzV5qcdZrF0pt6UDZ1TTD3zsxsf0pQ67k2mHUw
RRXP6Wscc2orBbYT/Wi6rWENB0cq5UaA5uwwAmDgIyuU9qHHCTnmIEul+ZP2TURQOU0tbi1ucHAZ
PgYiVN1FgicREWe6Sj6E5nqiVEubKtUW2nRwsRi2BWIbQwym9r4qJ713tGZfXBD06Lssje15SlA7
B3pGzE8YqHbrIaJIWNmEfEcftWauYMFwHdCil6YkX8bi2C6/bEdbWAwiLv1AhP+v+G7/kOKMB5yi
shuMgIZJI82NTyMr6GzMCDBEwTsLLd5fBBlBJF12RhW+mJLENNAOy+Zf1Wa6j/cPhuFupAVlPgag
Rk7598h6p7qMRsn0S0jwx0Cr9tO2Dpo8eubUA9akbF/nVusmhV9oJ9aD4B/hHtjCIKoBkFaYWcDa
D38bZJPy/JHkcQmDQS3IbT3GW0xYNn48zrp7qZN8G+jCy5lS60sUQyEQB5l1igF37fJfTtf94R9F
bZd+YFkT79vRv+RkSUKfGJ4+ceoppB8d2HyOIYHA6RfJ169rAGGRXdirH3xM0N1pOQa77fmQClnN
rjoJlbPkFl0Re+OeEgKWJdM6uBJx8z+9MmhCKQV2S79aCXznQEMJBT2L6onJ1rYzpam56Uss7KbM
L6+i64c3lYkrNG65KLjgYa6QkjExMjnsJxZ/FQs689IP3chGW7T26NvUJFsBbhazQFawOls1jqnZ
kntVgwVig/6obgp+50HyA0DEyHG4vjhwMbwI3yDbX8UruTKYP7uTY+X/u/whC42vJtOSqYcDmWhC
Sdy9Wih04gN5gRWwccyBJ7ao94fOhRJbOmlX5NPaFjjfJhGJy6S4BXyFPSSgO9orPeoFwTY7SBTr
aa8ML9q8CEOBAiaToYcBxQb3xAKPoymyMbJ5nhEZ0DWWFW8esv94mLEnDnAAgq0cwZELtEZLJf6V
JuO4uKRfsTo56SVgz2Hz0AHlW0/CEt3p/kjBb7V2g6mqhHxWq2VdpOQsX4sSGvhzvEvbOGP3P40r
lcFymHgYOqw8l7pc6RuyhJq0OJMmYZWt/YL2B5qCnz5Z8fByliR8qTYsxuXQt30KlKus5yLSY4bo
J5f5e9pEmxhHa+YO44GTcs+NpGVqp5ARvPaYaoGo2rndNsWXNaxICJ2+PgX9qEAg26rfqQDX0eht
/At+dUw+aulfJTaDhNcNmOzD94qUcrzS+W8SnelzuHGYZXOOGlpI5FpRRg/avbJNM32T/lx5e5nE
tGfw3e5eLRW5Sw5/v0YYIC62h0YM7R2sG0wUy2zY9y+RnEjf+A7ukMvsbe72XStoGPxmjJcPBuF9
fncbyktI6Hz+ypB5fO8Lsj2z6ly4YByK32Bg053h17LO5xRK6fwsxscVfK4Z0H+/7NqtKjMhx5G/
/LLH1xCGcM72OKHVJmSm6wthmCiEHCK3U+xuPy94N5U6XK4qoAcq61wHU5YCyo8XAPVROFtuM8Tg
x5+BzylMOWrKmV5r7uUEZR37oKsGhdGkPsm0mOcOd3/hA3qQz08/cL4cHheBbiu93kmXP3holjWK
yduW5vuEzkqmLSp6dJaFmCmspHHW2UrKzBC9wQTImk5qOFb0okKIH+yTuvETLYWmhQxdHjey2I93
aGAFUQSQ2gj+S/UgxbvL+ZiOGpEjXiT2HE4YNhifvEwHYkyiteXh+4y13WNhVRRSaWX1kWjUF4Vo
IVdD07Al0rvvKn5i1jQsfEp/M6bCeIHlgQeGNUixZLdfaYQDK2NdvnEe8ImnFxpjtyuh5gB+tvtw
qHUERpx00M3wbGPCPKdM2j8lZL8IdmFcyxFMJHbb/kot8+lOA6lLEo+WbZSKGifYwxqFf3cq6ZSS
NDMir+LVeOqjQfV+a91b/qhVqQOKaGSL4qQfLZmaUBdcosHEXaDfA4aHiVQa+QPoCHbetuvLXheJ
gZ3aCG5T5NScL1uyzLFSL54UBs7KDmpe5h9Oi6ITWlCRSNtkKGQNdvTtuayKzsdJkK44GU/XCPgL
UxKu+y1cxFOIaG7/WhAXMtqU50gtE5HEidgU1oan378Plmuz/K4C92BAnWlKb4HE6aUPFstJla6B
ICvTKbwTn/hUfn0E54un+ZLXjquzncTfrBnrYBKhMlOgHUs/XjLkWcyXZ0H+aVg/AWQNpkt7OepS
1B1S5ID2Qkxf0+RlwVSn/5kU4LymgKSnqYmABrS5uQ8SmrsiYkYcU47ec9V1aD/Vgqalxf5vOBoT
cVcSXlqqs3xNocX7j+1sSUim6MDFllXmv0CQabWh/ssW0gIWuIAfyEmKZfmgIb/9iAYFUHM60Psn
HH37z1DDpjzXgqB5/23jRx+RcGxkgNXIeM6XHyG2r/R1ZH8lpzKnOv6wT8mIeIu36GZD6qNwtvA+
82OxZnbrTsiNS7YXtXt18+HBBdJ4O+y2LARqQxlxEnvBHqp0mNZdkaxsujSd7C39I7Jc3lceWRuv
7EPv1Pu8nJbqgsarITYPFlUTauRrvj2wsTiQL9DaNTW27Nq4IHARHAdmxf05k4DyV4kOMo+L8X1A
WP9qh75MviaBH7CXS0lXmCiuaVrVpLmKZ2AWSOfky3BmeimYdbgYe7EjkrGnIt9S7LL7mBNgrrif
1HOVDxHPsU0TPpAMvFolfUmULo170e0Wy2l0QSUk8Q4m8p6BA2XuYaUsWkZA1IuWkw66vneLMC2v
lPh5rArAOs7TiAplxdCXYIZXXT8tVtVxudlrZRqEvGAEPf3DCa5XBtAhNnboAnyop0x2JxoXwmv+
v17+Jre+I+3Be73Fjs1SfyV0FGy5SwHlzoidaPRgttAvuYCFjHHjMZZl/zzVGTnpe+TaI6viK6NB
pxF20qyphfIdnP6M3Z9toGfEtGibNklTxKTKzK+MgDjMJGJV67uxFXyUe7gfVTOg1kZO8QAWbt61
3EQvD5ZpySBbaM+boH1FGIFBDNuftWCMJFE4OACRAHF0Lilf91d0ycx2kvcQxOdzQkT1GaED4hTw
niZDI1dfkQ77e+erZ0FOdEj5L3yRdXwBcmEDIlAKSF+Kxp0pDFoQfJReuEa4w7FCbnKtvJ50xK6O
J4mnzCBUApdM1ZIkGEnWs2VnpWeUfvK5iP/a0f833huHs2oUyEaWpGh80ezd0/25jlXqFXcC+xyV
pyqScAfLXY9skDC8F5G4lodHWdfBCSv9EySBH+kzH/T8BY5+hXnkgAR3HNGzOYlOj2ApLh3W2xn+
C6z31MNYA3LL86t0oE3ts80c8WEmUUuqJ+yZJh2qNNDR3udPhmG2l287o5cRmAOfVA4NnWZF5cXZ
Va5aIeuOcmzbF8l/wwBuHYXsd/4q/WKPW0X1Zme3vMrOQDX19woQYSS6ngVeXHiKYJSKXx8gpdYp
tD2b2OmIvN5ES7AWRokFZwyNPemt+HH5xEIDBd++IMSRV6eVdd1yLik4c892hMGb5mgLNbqYgyTt
CerzcGKxikLJbKWg69O0pmwDnEFZNJl32uWX60aJ5/AopmErrSaGt2CGjJ++ARaOPuVTwsb0XPTD
MIH0zZ3ongKn5MaOD2wDZnkabr8ABIe1UM/8DGZIvFJKNsfsXCLE6qDcSRO5Bmm7qWm2S0Q2Ahzv
1l+xZZk0YbpJpQ5ikHPFI8ydzJnR/mspcJTR3OyqstAUMFu5QuMZt3PsE99ltzl/9WASmy7j21D0
KOTz7sjgDTrse/RsZ3zsM470EVmw9R23iPbZtwFTdl2WCy4r4lGQAC+pqamxKE5bfN7BbCSfV2Hs
iHBvd8J8Yr2nIQWcKFJhu6BcwHowDCtxU911HeVA1MbWkEr1C+lGR6zwtAEYrItuQYYQVM8sPP9p
utw+3i59ECsCKcAWK1Wn59T1Wy7mtKvuS7GrbzJii4EBB/H8sW4ztOgMPo6RFHI40IlPLNU6z0V4
xITSYWWIlUaoc/syslm6QahrpV4CABPqRky2/xL2GTOkZTbqK3AYDqXTfiREnM5Bo0cfqM7rS6Ob
eSTeB4R6RnxI5O4pgfGjuYZbTs+xW+uFtif0SyLUkmMGqcf7yV7KRuQtgmgxqBUE+dzLHjyC02SY
ee6XkZIJNXlj1kqVYpG8oanj2w2zGno4G4+t3/vkXn1Bxv1bU8ixJ6buFBspil0FmxKXK9e2XhSJ
G6Cy71mHQvEPQ96jDMm0ASXlxWQF6e3EPMZDjhG0+9t0WYyhYu4nfZ6ICsw2khUrEy7q3FdjUP6h
jIue36F31E9mRc2os5KJpmgCJ/JZu6tO9r/6R6Z80+4kpay5pmEkyl69yhGtk2hfAR3FptCjUDXK
REj/rvgDkVbrQDayiDA2P4+auMcvT+rYvgMYInHReIqJgtzgcdddlJNHZBxX2N6WdhWJqMXSgduY
p8YL2w4BqaYr1xgSPn9mhaLtoQznfehakweuuidqNNFNqv/87pDFbPrdAN+QvL2ex6yilWYBHuIs
PJ/v9bVn4U2hb6OflbNnfo2FgSgEdlB4uulLbJkK7AU68lkFUooqsoU5Y4IA9UNmW7rAYSNOZPzA
/3AhQWP/HtFxvk5rsnf8Ug/EWzbeJ6q+Dym0QuXW+77x4JAq5/heoQf88q9YOq/1EJHpdHgUda8y
9e7UkK9h860021qJQlzZeCR1wnvWessDZxLX9BftWAwd6xFodvVS++vEOzunYc7fgZK+mm07BmBW
TrYPop5aX4yjjoeu155U9tnNH6S+ztqRqGpwl1wt+/Im3wuF93RVImLZ1uEe3aDn2DSQR8rYccVa
A8NmYQ5V1eCKtfSY+6N++fVzu+uc4eY/fYuiIBwHyj6Z1dIuUUhPFAwRqWs9VrEVyueZ+sf7aknD
JrowzI2S+TwFre34fvUwW1jooD0NgtmU0oYWrbYPQoYDTFA3P2FXj83dbKPHXoPsU10T1aX+CQmo
GnOCiYFhV3KrvMZCSMrZMQdeIXuW2JXNoyF1/prVAeVYhCE7IkIwMnserZBbIef07jUNBWyBOAH4
JuGUNh8YWFcPftUMLubeH+TSTl5U9Q59d4aWhWX6yGAngsZuiifgjrafb0ULs32V/SpW607uDw80
oLgahDzLnZFIg/JidaE7NDBdzeexGjnwezp9L1W0iOAxJvV0BiNcuebad/Ieb+u6UUa+DcnNwpha
9Gy/DAfDE51Fqxw5YbKF4AQodzu+rHFjB8Hw1fE0gL4L0jpw611x2xZu8TTYJZWaLhWCzHwPsfWm
YVGUJmw211/RNfye1i2yRVUP74M8KEFHrdcjCiv8nY25sFlpQqz/NXKeXQI6oJHCruUJDhnZmuuj
ontpJJGKUvq+YI79Nszkdq2tu8IB9EX4pwOVGAuDZQYG/+I5JOe2xi7kZ/7SOxDkgDc4v/+YWxxH
fv0XM3qLut11FrCaZ99FoS0c/W58QdwlWOzpySTxPiEBVC6kBnIvrd4sJlF+pyo/TqZHD7bdSR3e
W1uUigv3bMzNFDLvXtQxVbw+3BOxGCcNTWJ7KgTIsmmebf/jcEQ2ETcbTCRJEvEruAzH6QXuapJf
TNEpelhyL1OyJFkJduyBSwiAHgJYaOFFW/FdoTCM2dpGqv26SpOpiVnz3z79a2Fiaz2hvfzoK3Kp
ldbRbvyzri7Yf2GuKoUXASAkMhOFdUowPTpTtqXcCt7GvNz5aDQDYDXl9K8Pa2OyD8lJOpdPlOFg
SA0cGoplF1ESYF318P5brJ3toDYQ7twMyAILjeWVPo4wq4Cek2MfayxVQ2sL1ivua8ROCAHAfa0q
10MPQgSQnkNbYmoM9qh939PxBEaUzVbWFUvbUTiQL5/DrP60OXOinOtYdiGn6LCnNws+GJuVXrZ3
x/77xCa6dVxjn7SU7SuZHAK20e+DcUHh0twwUH25iY3Nlht0txR7BXSJP3y991syaEXuNGqbK1Ke
6DAYcuw417DEQCg8YxGkd9pebpggmenfZkjDGGzDwiwM2Epn0bJpnB/gN+wcpZzPSyOClEu3zPMR
5aCSO6hr17cJu+uRG+OQMkV0b5ebMitFSG+qWYgR2uLkj5XtD5hlkRI+7z9wgPV0ELOJqsM9Ep7b
I/vvr4W2UXspR8Pxo68hLyhplT1leYFBKpHBRnOw/xdi3AFLBun/eNTjgKzHCqFUtaPLmS0lfnFe
Y8jsNOpPDHkRS5tZfjN4OCvAdR0CHCo6xLAFqdHxz3b8Uebt7jnRXxQwvZ588QxHNc4hDrya9FQT
JLmN+YJQxYz8m+NT/zkZcaGgVKXtc9pEb0kztRydxfBnB17G8FSpIYIYzYHSx1zxrm6lR0/L5FDr
q/UHa1Eftd2uCy918taieBEAztvcZcN4SxuP8vZT6faEswjIAGpO/4BUr06yobFw1xrA9LB8176J
zILfI0MJ5+YSnbhMRNZcJU90KZc/pIsJA0IDI6ZFJtSkcrzN78uEUFs1gMMVlPdEJHfhVorXr9wZ
uLoYli+Wtl688MTFuiKsM5gGrYm7oMawBapg7Q5XNhADqJkOi5bvJ8n979RmmtxyFfdIK57XjdMH
AYwTN7PjfheRUGwsOWEpqBRwULqrJBBZLLse/B7noQX7izyYumhyRr6Wq/lNaizXfTX5ZqKi3um0
gBOpjJ8+2zOqEGbCY/DT6xdf5iV94hETU2yBM5Q5/7z/nCjWfOBgHxbTJGd+kULzBemE0XB/xBF+
DbAFTzzaLAylByN9suwyqRAD/IE2QX9Cu8SOFniV/b7jx15OeSZZhcu1xc0ol1W84dkpAY24MSBJ
Wf0K8MN5zJdEL+yUadmF+fmUJtX6vCwpcWa5nkcMvSHR9/4rFJzNnuABLTCnjYrpuyyUu0QHWsc9
0SP3KlzflWbB78+gC1y6nYdvs4a6VeUERE2TIYxNc73ibytykTbW5MPZ280X60FExwvPFU1X0dC7
l68UHgc5qKi1qFMoD1GFCsgr6ivdME+zkYrVQFQf3EG2QKWwjmDrJnAOGnVPmY2b8qe1X7qchRgq
hyL754AY9rUbpWW9jiYnvcM0qUDy/G8/Yxdhi2eis1PUqV9LPHsdQqGn2X0pvRiSrB6FQ4Rgcw6R
0xY995AJ2TJ5KH/wepLUshzCs7nWG5Pttd5gcs/NqHBrcIZeB1QhdyoiIfVQuJpzxJGlmp4FfgQq
gmu0xk0bLcxJTJ/VYS5c9raHq3keoFTt4ERiRAA+KBRGNMn7VoT9njImaIWzBUmzq900MPZ9nH0C
pGdzTG2bnKCyI3y/TvuZgml4MWqzj4qPy7l7IMOBkuNdsoMviiqejX6XvRx7+Z1Ay5ynXJ8B8vQm
y/UciybYn23lOpyLvRFbhqVOml0FgyP6WDb5EkizDxa6u1UMAQuxrHTUwZWI2aCUpiuFVpk8mvIf
6ZyU/jl4eng8AvIjY2iHwVR/a7T76Nht3Bo9JGFKNqV0jdot00GTtbJ2zYad1Gg+oxm3iWICLK20
uWfZUwyPpXySvr+YEsTyTXcOjykp/HJMkqRGgqRVTo+QXB9d44ShvFceH4PGND3p1SyPgpd8k8M5
ju7tjRNaEhkoSVuBb09oUtwpt/QTJrh6lF4nFMlPkX0vH9hebccj1jHtGllow7P7OjmBr10TUz+u
ha343pSWCnWrW4QWEcVXv+V3JEWj+mC7WNYzHnd5mtgHMT6TyY19QLTvne0Iz6ryrMFgO1IteYJX
VdP3ZhGernipMNwjiZC4Wlu1WFtkCRzwK15J2MN4Gdwef6CDHabRBY2f6nNqK08Q+KuYsrZgYwXo
mgLmBA1VDRGgjjErPfeL9CJ6vpbTAToEmZjaRq3wSAc/Jk5Kzo+5ylDywGsEaShYqXUuEUVFet+U
WXCWLZvKHQVFJ1bSnVLb2zJ5swxalb4bRHxEe8tzCkg5ln2j5j2iS6jjjSLgqR7hh5yZl7dLI30c
6Twx8jA/TBZGuX+XXDSTSyooP4xDUiy8jidslYAj5hnx6Kxo7yRz39ac1hC8/xlnq9AwKy9wZShW
ARyE7TkMTttLhZsquF2hV+gQA6/DV8Gy8t8fsGJY0bHoHtjRAj2VVqw65rN/ACx/lngHhQhbYz3U
o4x4SYEr5ItORh8Q9qNfFh5nsU52DQWL9adRLIQNRYywhDR1bK5jE5oNc/pNr1qUF9MoyUfdjeZu
FkOBF3CENMy0lt8qyyOvJNVEJXIT50RR6QsldJnwJNT6luLLLlTMyzXc0WEcKsgHFl3l1XyIOo3H
Rh739xXPvCxkFjYyMgTgivdnhShLAOidor0iFw0eAi/7qyJGnPHm+S0+nt8eb9YyIAfRj+JH0IvY
Z4X6XrVlf7sGxJgsmuRypw5gYZCGJwj46buIlx/bnTs4VCTBWXa7Ly8emmAaCHSzGsZx7ttH6lwF
n0TE6x5z81CKba+KDZsxfPDsO03AX01KkmgDSNV2LOPMxemCGSJLsruINrm5g4l55v5xJqk07BdX
Jqe5SQ8Y0L3gm9DAMjdNpG8R7tcs3cyYif3ZuZJJoxrCkZRfQEtoWYgqdyW9H48nkAvfdx7jqfV/
hfDvOi0JRyqH7n96jtOOGyaDjrJ46Juk837WZ/jKMR0mKc6ojdvyd+2XxxfJ9KjbhqJYgkr/zc9Y
Yt/WpvYB4VJpHrJucQEGhiTQ1xeFE5Hms69aQffCzJdvqmDDN1lQlVgxK50jc+YZJbQkSTsdoy99
c+fkT9788Ti2Mj3LamLtQVdeNXojlN7dyC0yBSft0Deue/i9a/1mO1SsJWI+2pRWUYMTWsYUqj1y
dTcaCs+TzpUcZo57sx0WHTSZtoYgsYLkxFbacSPdamEg430Gh3bdi2DDpW2pPI6CjLGBtgtOL74b
XIeXy139NY5zrqPXUWYbyHOaAFSpK9pJ/a25+MHFM5DYjTOdfiGT+Y/mQ0yifsg2I1fUMiUnL2ji
Kr8AADOwjavgZmlbJyaVwVHehZsbuacKFACG6ohLCAz+qYLjYQDvOM+l7QcgDViqF6oC2sNJhoP8
i1L+S5rxxvu7c/wyn/NzarnmXp7jUBLxQwIrAdDBsLvDVr02DLbBSwyF+wEB6WixzO4A1uLAzDNl
PanN0cQvEFBhhDc+GpzaJ81DL5P1VtcPVihI615D38gMoOeLtlsytQ63biAnIRMhtew/ByCUlBGl
eu/X3/fG7Un8NggrSyVMW/iXUEskBbcRJgDj4iueFeGMP5xlvYyN6tGTDFGpulmKE9OUxjzSjc7G
AyYH+rwXIWVBBZuj/IB75gaGhb/qwatYwLd9HFnbSvCxYRbaSSN5kO/En46JL6y6hUxeF9Pq3tfO
JM5Ibvtkly+Je0EQblN0zIPqsHX3NNQ979rTwsGwzclwfKcTSrpKpxeT+F2dAjUcrZ0tC8KayVa4
5l81E+B+zLsrxx9FNOttN8JY+RSlQFtyN/IZE7dw9ds3IlCRoyqtX0s2tNZOsSxT35SUiJZKWyiF
CZTY7FM4A5AAkmzyylF+84BVqJvQAKO3S2OeWpl3cKtsJLUvlV4NxqKNqUyAZLBEmttSrK7DGLx3
p0c4ZaRGHVBlOkaghFhG/1/r8BTgBYewzx1cYPWmiwj5Op+RtxIuXuNdk7oAPBtyINX91WsuTVKC
1C12HifQVYzNkQTdXoUS1hmqPHK/fH+yvdg1IV00YlKB8d5lGiCSQPGuKpOpTsezEfIPjuBlx6wq
sivU99AUdcjJPM6DS7Z0fKMpi3cm8AHPPTgeAYWtakX6P6dMYaLRKQ/wJJedpT3Z/XzT1X2JLieD
v7SZcFvQnkSzhSzKGky48g1gT7pIMokTiw3OEX23GBy8F9DlpuBoFcU0jrc+1YIAeMf+IT4/pW3f
2oXcWaJsmFjNnNYuGmrhwAzNE0UxY1QroHYp0arImZqFBP8cznd6PqjfvwIXB2xmnV1jMExccxkc
kyOhsYfllbTTHr30KnLqFkZQTlrgI2r9NpqzOrMjmgjI7awDJr6+uoc0682OQ5rqh73TMlfD9G4F
3eAsgt8UMLhrLIAHiuU6Os7RIk22KIwDjld3YLO9osusgAYd0InUQANJsXF0lXnHg8dAfm5PnApv
J+jP3dZm/a5Htfgu0VGuTJb9sFux4YzSRZltndoLOms5wFVCXNeph57Rgj6WtZQqQ2y0RNpMpRS1
Lpblfy56Sl7FUcrreaDlNQnf/GD97o83v4aL1v/ZqEH2d0mHh1sh++VT1DfmTym7S9SaS+sgC8w5
f30tDEPOfOhuxJQUPVDn+Q3mKVEW322Ao/26RHU6CrvtZWGsjkSS0PmcIlpN64LhDb08gjEI8gKQ
7/MJ7je9VEu+CAyzXM/B5Wi1p9mAU7m6cBD645MV2vZkXshc7hB4Dkbt1zhUHudbZXOXU3OKYko7
h2NSw+gW8PCRgXbKnTSxGELCjms+BvwYxxolhCUMsH1qmSt2c2FqS083RZ9Qy6Td7d/WE8ud3ZeV
iNv7h8EOlpadcCAcKsqyUu9t+Wd4Hez4p3KpTcIq194ynNBGAU+aH9YblEyIJB6hL7e2M2crRndD
4rjtXrwNOxsTK47PFey6yhrZxGAED/QOgJnVsgXz4Iad/GzS6qu8fyWbRMOmOdzNkLYrQTb682XS
HvdnprkCIx8Uxjz8AicwK1JqR8Iu5RU1nAHYURD1XFljWisGbXa9YppJgZv0NeTdMHw8q9QRGnKV
eBQTApIC/NPR++A1jPuXAy5DvVUPKcZ2aYfA8O2mGmzw55TKKbTTxif0A3zAnYKI0Ijobw8kE25P
4BtCyn6/Qhf967VRgtjiNk4/Sg7W4wRXp1sUbxTs0aYJXa7YVm0ohXLp7KCYIJQg1NkeMJig5gq9
JDA+CtVSM4jG6YMAqSaxBBknTQuFgZC8stzv5hflW71PvxJ8FHXRtFXCMxmvu2XuwOsfGfVXa+lO
xvwxYCVs+ccl0X7kfFJCTT0cFuoniHQZMwGObr3SGTZW6f/Ukzh1A2dkV9KWcCfvBjFVpiu0QxJP
FCYGXQD5gdVrvZk27H5otMZ4QIS/q9DIsv8pqoIN5VQK1zrFiRGPgIu8EAlSX+eoI2ZqpqArJdfY
Z0gaP3Il03W2uyLOH76rT82fdv0EVFAn2m+QGj2xmjDW0xCLyIzxltDz/NnBV8RhVPkqzyz6cQCr
imb4X4tgdvGU40HLy33e2VZx80l/uobSzPQP9bDcBjbe3Qql9ihp4Jim3PUcVRKOKRwVgyx7VNjW
r9+SGITMh8fc2kumZ31ENcVYUlrfyRYU+QDhzkGZE90JqlNSF7wTi8so26NllJm0PNy+4fmW2ol3
DQb2QGR+q2AGKD+RpXOawhvxI9t04Y64E24L5lOPspQXVoYpqaG+ilWTrkiczqWF81BCcAGk3EjE
O933bBvTuEsz0at4LN9XW2KS+RgHuBFpzLBypBBZ0DnFuRQGH3qtdqSznzScCy/qpbbfi7pW2+qt
EdVFqOsXawoN59vBHZOtydq8hWyycOujiDf6iJp6QSEE8JxNCYgrm18/86CAYJEPnZDzBoCDC50K
IQb0e7XqyDvqTXV9R04Qp1gBtiKyE0ecq/XM4JXIRmawJ5j40snf69PNqV8LPkRNxflC3kxao1oN
RB7dZpArVxaKZbrlR4TpEeSOGipQRIljTQAqQT2uZCHYT894OvBVQzQ50yjy2PYvMmB3QGXGdGrL
jXFVgYuIjExBWMNqmPmiBahqr4Fzn7KhmHupuuXxvsbQMNJEEPEBxaGBzBWOc+MK6Pt0QmbIK/mB
VWHSsZVgQmqdElhjZqLpSwmF4eFkiY80QjIf4PQ2imzzjK5T8xcgRbQshA7DEW6OdDNZkonOa1qq
JIFIzsOddmnT5lIgSr2ZG01c3DlfO+5J3Q4ZhkbUxcAJFlLJF3JaQp7YJMlSw7CnF0z6WfL1qyru
12foa+Ind8pNW54UnkpMtw0i/IQk4Ah1CuDnu8cg+XxMRHW07xG2YMKiz38ZIjNJJ7eFHUbtNYlI
o629CK/XkDZk1aN5qSvrHEWkKFNgEjrCdDy8fA47ibG2upr3yxhuHDiHJ1jgfVAXEusD4cy0bkCB
lk+d+bUimaczb/U1Zpfaz2CwJWBaJmFh4/APTZHWL0I/X3RfgAk1kHhl7uSfWPtcIrI7b60tGUJk
XQTPe+L5t7iS99nO78Z8gta7p2ObolM6MbpD6QCiKiOWrKjhO6ZJM8Arpd2PxLUH3YwGiKaIwajQ
tOzVQSAtEw1+uyDuRc6lef6RAYdhNxq6Ix8S4V4+MDk6aV10FshAAbXrnDVMJXdax3d3Ygnrz10B
RIw3OSZLDjvv+NnVMPFn15rLg2r+faDD+giEPJMZMXKQtZW7FFx1UF12drEfGqN+tmbavycuaY4K
NenZJJ9DBQ3QnqDwiFw2hlq9aXJqjTLZhXfRxRFAM6c20R4nNom9MzWpSa18huEoCfrvM+kMG3rb
ORi3Tnpyd00NHm0bhyKO1LgX95NwHwsIkTjhr/CpeqTcyephT7xGrjPOikhETDd/30mwJeEhBuK+
a5/Q2ablhKtK0D9wRnoSJqP1Ix210YBzgvHkO6nQ3Ir97c94fVqR6IQKj5V/pY8JTKfBwm7nMQzM
Zbn1IwCfxGRDQiLsBtHMwxd2LmH5r2EznKeXgD2AJGGbweA2dgV5Rn+r1MCzieUHK3NUgBwXGhZu
VoLtgcLb7Enar1Hlv3jPkACrUFHEtPPZHZ0m30ApgETfihuQdrfoGBF3mtczFpShveGDT14xt1GF
6rMkFJHeG2E+U1eMlQxCj/ANkNFW4j27Y0gGtAzbZEJ1ObC/ut7PNYsONDZtNEpHFZVttrL1oXn4
1tQK6fw0mMyO/1am+XUUzlE9kNtRKCTMCKAQa+92c7PhyTkKf+Yvnw9x6ajXFg8qMUEfRRpnJkWj
ogDpJN3Qj/Wj7nhITXBi6R/fv/YvAGdy13Jas/n4fYIUAyCsBxFSMPzErvKe/Etiz0tXF/Fy51kU
26Nso5wYy01yVDfQx048uBiRHkiyKIxSLXRtgTxwbx2OtS7o3bqF+6ggjUthkqGTUoVTiU5u+jsG
ooFOJIwo0nPBZ6Kz3FLXs7ub0GiC5UXA3eoUOYWKR+YjHEaqDo2V8gUR5Bz4B/hSsI9TPA4dyECq
CDhqPV2PjlaL1XNRGLOG5A9XUQN0EKsKsKER2NNCNIVmaT7DsI9/kKM/Zf0hcpTGuggnEw5BlB0N
9M1OPTuH+ha4qSpPP5Il0xtjCtdAVcqemV2ab3PpWSEQyGRAXyCI+5DiKAYttfpCUaw/MLyZpgQG
yOvaaSd7qO7ccUmZny63DXBLeqItEkegAg9ChCxleEGx9wLttJ4VXR7C3bXeLsLCRUS8w7iVmUDN
dg+rGOo4BTFkdxDe5cwG8pOTiXYDRlrFv2LRjZ7IfkrENDGaawzQCk1gpAOq1LYg1mJwa/1XHR9y
ar7i4+7ApVRTIMf5xbLAAqySW9OgYODC8bA5snXmPQy+qs0aNzag3MPC2YOiQLCDKMbM/HOxZBv6
ZiNjE8tMZCx6GthUGJLMliH1+kw+zd37iQbro0AlIothN27DOUFVKPfdpyIGdczN/wHrPdjiczBZ
pT8J64CV6/gvMsf6zhfIhGy8o4gZOIuJxzNbEmFJwAiPDWm32VSjCpVFxHu85KbZnD+OZm2ZtGva
O8t/Ig0lDvvyMNt3Rd7V/7s70wNFGGxAFCitDTa3FRQNJM5tEC4DzhOl5clJaNQGZUEOUg0xi4qQ
6VJfXZbk4rpuLYSzFahmzqi18fzaWyFJGy0T8MOXa92151lA/QoufTedK4eGTnwU/7rf8kWrKLhV
wylGsc7tKRR0xxkpu0HWe5kOJYqvmhwMcpyTr5IX6/5gMzIKMOS1YdlGcsGKeElpjXtgPntYrp29
m4wc9IzJCOcgTmjihrBfwV2bwGagVzE10K3TEWUVCnwWN3VUjeJR+Uei8rNF18tQA/OR8UimNjZ6
SWk+nqdPTerDkn52iWMkWe6ASGB8QqRTE+8ufdDlT54Gje21d4uTjUnMfANiAndMNuX/ESYsDQQp
Y0GBTdfONsr9LxGstoEs+vm1Oh8Wz/fyjKmo7Hr+MGCsdHoGcFfcZKO11umpewZLCQNXHOoYO3kr
TJdb5SG4ulYZlysalwc4UbwXDwE5ywP3Al6JrK5Mwi+UxMpTiP9bDnge2G54DxGfN1cECZZoH59p
T59DEaaTUARMGZkTfCmnQFGQ/J2szAYdhwqoJGIHCwk7vGiegV/3tl0V+F9bNTw12MykX8quV97d
uf6X1pJe758xMWjD6mr531If6F1s53sa0jlBCIqohnkRcIqsa7yF/qZqpj0cVG1tJqe3BdpoJZwI
mwwEoy0+bfsRZLjhA7x00i8/dO46wFZjncuVqXGFkdjzgkzWV9fNTY3jl2QyE+h6sRtbmEo0/AgN
aNLCB52/VG/JrSh2wrXG4ZE6qAVdOKE0I14d6GNyQJoR4z6CnKVPwLzSiNlli6rtwr7MrDhBwAlb
zNN9ugcjWZBF5GPik8s/BSiDrSBtwzb1+c551DOAQoZCJmR16m0an5ap9C1FEhQITf41PRl2w6+2
dP1XvSDOL7Lbi9C4+rFmsAoHwmcNz1OD2c52q/L8sULbbbCJ1or9Wj/zCWXOTY8koSdlpn7yJMn4
LVnpsoFy8Hq3Q0rbMwS3hzEvmeDyDPRZumeC3aqPn4R9K7vmN5az2WXkqO40UqnwpeMg/T9hiCx4
Nl4G81HbKl4xBUqQRFpJPxcF5fqolFfa2AOAWInJRBExG1yPYnXu2KmDgM045ogRZbnwKtI21tR7
blfqNMeSZ9tZnsVBH7gqr4URPg1w+HxL/ZG0mKflCwNIQlrIqVxNoVlP0ew+7LH7xkgbZ9yrflV4
KoZ0b0YDFZzUeEpIzZYO9lml5lBZ2LyoPwO9FpetciCQoGDJrXbMbuPeaMTDXCEWPiNT4u03hBiL
Vy075S8aI0Mtvzijx9zGBAJqLxx+eAUNFLWvU+zrxQvDOK+YphGXmwzNqr48r/Xy6EWJZtHlCLi7
EYMPtCdBDfkULcSoxfu3ezO8LbrokxprIE/JD9qgAgImNVWy1zcuzGtiGBF45SN/EMkjbyiAz8Wf
hg5tIkDt2YdMfJVOQw44RzqC7UonXzxJsRxv82qF4Q/fcS6cbM1GBJk0xVW4ReluJkV9dwdnAicj
x8+91sJU/2PjqnOpIsuX3l1r9OMsL5kuUM67OTbJjpqrSIpBAAnYbSEx1A8E5NLyyY5dvAjbxbGJ
IEiAx+nr8vowIDiKXhwWh1MtmEeghoskzR0p8ipw/+gQJwYUyK1mIp+RNWsDRd3jGcg52S+V1mxF
jWsBd/RV03IXVgOJEfkBUZJGD2vtay9NHwchM12APX/mvtpKjoYvDd6J5KMlxP2lfNGnVHKhgCuW
nW1EISFD0+FdxOsOmCSTss4+7fqz0I0ZaBD3+6T2MGzRzkIGj9H8+ilTOMdaqFulmSUpC2TZ6Zev
9kCG/ikEcOBs0ZUXGYBwz2MgAVnkP3TcuYUgBqeID4hIov9Z5CmVbNsgz77BO1LfFRetF/8Jem/V
RpZClfFU/STtsRuCmKSdA8Yc1cIb8mBo3/w4kGEAo33mPUmk6pNHdmW2rTRyGKjGeLzp7f/mepBK
wF75xYri0N7XD2zs6GknOFAg63FtP4rhNnYLvhAmb+WTfXZpUWu1A6ucB/JRO2L4tbknab/WrFBp
HILdZK0bBoBDbyjjf69LpURWPkWUQpqz7WK0dKnSnsX2HxtIAy7KJFTxSXU/JCORQuMzRqD5/GCR
wubgbRsahrewwyFDAuYSQ68IoIwCyfNjoIb4IFaHPvjto2Nk4BaJ570f+eLx6VMt7d2Md49EJwVw
n7c8YlHdZ6j8EqF+Rtj2qdTmmNyI8c3uwAnrGW7Pdk6l7mCd9DA5xPCQf0ea4gCVX3AhTsSa39hL
iMnc23ydOctucvjrcdpTIMoHbzgdxni82hctDudoGlL/YJI/AfWQKu0XVpOb1HzakhNodJWsmh23
+vfREC1cvue1PT4N946NNgbXbEwGUMHawjUYcty9JuTC7gcU/E2isITKjXyK19+olNc0d3j9k/QP
j3ps4o+PiiU+/hGEj78HC/t3OG8vY/pbOU40JtRUZZ9VV8asHuc4DxEISWiazITr1yFN++GrlXUd
ELjLpTPnN66xZbykvvVWiRpktbSfaKjne9kVq3V2KZu0hxXZv53y/F3bVKzm+OH54vZZpoMEofAE
vyaas+K2H0h5Z9HDirRAoHogMGeFLaGLF0KyX4+4NLQaSLY8vfe6Blu/BK7E7N/esxOHQEVZZ1aY
zKaBQaQfB+3WZRVLZ76JhWHStP6g7EZ49Yb9PElrQUKm8Az3AOzY36rEhibgoiZ1kDMHfRmfBQWL
/Tu9jKoO4I+Fg2yd+YR3awa5l98Bx7xkQCGQz7qm+aTe6Q+ZZ1LfpIzURt2hCtnciGAUEfG5euPo
5jk2S0WHsVuJqOBeqdlZO4W4oqslz9/AwbqKYBzzJc6zSBeOTnFtPqnJvJwPZgbV8iy7nPbbqmhB
Jlmqgch00lE8N2Lpu2zSmLXfxdLxmpp870SjNEvjchs6OOZzf0A5okDbH9b93PwZy5v94qd8PQN+
aWTh+2j7secsZOdj5JFFy5I2F84LBb6kMEUTcluLypLPWsxAj3z9MT1tS7+/+dylQCDzpHUhpTFV
nOG1uhQjcJ+sGtxTu4n+yd83FFihmOossncz7ryxZW2dm6K28m6hhLY/v2M8MXC0azppURQcc2O2
th5fIZRSAM6dFtGw9QOtHBg4gS3g/rizhnxB69RAnaDI/KBRhN/ELhW027d9+h3bn3J9NF5jdl+d
JT9RL+ta2uWYMl8rsBY9IyB0miRBu0O+auzQy87st3cViI6QLeSelT8b+4BNkqTpftrL27/OoCgt
2PDAYxZWWN2cIpa1cxdBiUkFr2xru2a6x0UMEvYn+I6L9Qvy0uFvtf3qs09h6C2RxFc23OsaSrVd
0E2SRL/lLABYpKj55ohui/Nk94mVgLwETAYCqAVIF/iew+IzsSKb8g5CH7fOGmIuJqGIWUkbJvVy
yZPNw6IDLgg8IeOx2/TILcshZuQVJel7vqucNVva4ZQ8/4jFIzai7Y5yUmK2nnANITWI9JNgKt3V
JKqCKzdIjgG/a4OuloTgHIG/KvmqkjBp3iNgcbmW1I8sR8KDX5yeDbPF0MkMw2KEoSNPTpQRdCBg
mPRMNAnbkuBnC3o1SspDLxXoq34zvgez7Fa1p5m04iuahtioQbGUUdEf3te3zTiIJvX1HqILcdWj
hYnqzpTNR01WcCq+V4UdLCsFQ7OjDULX53wanDuBzlGvHyTNvndptNXPZH80EuPXVkNtcPalmkxQ
EGnJzvA+DIRYvlfFFD55iSmOKrMZl1MhY0wfdSBILwQpJ7pNsUCLWPGioe/hVd6rnv7iHurFugDz
rEbhPxDXde6un1Hwp0Yhk3QB52CpvjUIOdoz8083gIaat5/YRiAaLyySaJj/FdVrVN1MvJF/tbnT
aKFsQwsrMEw6S0AUnejzMSvWsAJ6dSOLuZRZuAQXQv8jrR5Vevx1OPRGlvEeUABckA9rh4NZi4OH
7b75r/4Aa6YUfRC/Vy1eaqawuWYYJmZ8wcNuldq1Nocx5z51gsXmBSALjpe3U32yUj2f1V4uLrfF
hIe2oZSDO8+t0I1zhHRjowXcqKAZeJZrXretw30iV/cfPLjNG+3JmBcgkxejZvjzPZvyio+6WGkl
8SIqssoaLQkdzDNq/wA8uLmNRdCU+5qhfIQgXtU9t0Q2KuPIG8d8Hg5CdtZ5QPqovqJSelDWLgod
RrBveOVi0efaLMN/EdARcwzSG1hZf1S+N0upDuO6Rk422wJq52UiUrWQbhKlJ/la0WJphX+FarSl
9FctUCACIesV0H2u1Fi4rLRkOI7fGEOf/eZlFSNoybR39HWQ7kf0GeASdNxaE6aTdT34KLJD483v
2dZ3K4KzG8loNO0nMC7jwdOPFt03eHPdd/unq9xQVL8rqDtXAvjqEMTUY05HNlWbC8L+lWaJmVvn
Vm4eScrqr4OJeBOBSiekZCSuH753ZD6d76COafO2SIqbSkUbD1snBDm0ZmlMWEI5Rgxu6KE51X4U
jlrP6wMDzt6Wl3hJvgyIMqVZWauAw9LPK/mFlbRrToueJ/J1XuUmKdu8vlgNh6+JOZF6TBiITsIr
da+FBg1nl1OsoFWM24/axFpAhZiG7WWxw73INpXmjeeBhMD4By/bCqzLyXW2ZPzv70XvOy1VZR+m
qKxk5oMKdqRlXWz58vUeMvKkYks8Sq4mcn6CSFe+52w/NFwU9Mv5OXEMfp1VgHnK1UxtOw6yM9l3
L24DlCBQW7gw9clJaD3NbPNVaY06+sT5EwRzqm9NYs2exuBeVbrT8mFDGlRCxsdwb8fzLAn0SAm1
SJpVgXWwLt6F9eUKk/jpCGb5uOAOANEPtImh8ziuOkekTCkHzxcnaRIgIW2hAWu1o6s3VDdgw2fd
65WcAIKQfjLtYhOTAX9ZRZXr/hxLJBgtbDdXhVHalHoMiHFJhyfRtNShw3KM72eXsDGGjB0d8t9N
yBQpCxeD0aX+LuND7mXrDR7g06znbO1Y0NQLNLB44Y4LM6eThGVnqHQEvy2clNAv4o+kPEwQqq3y
QcHu4RlWfMcQZvvUkKmuNNoFMPZtql3NURS/WPsLIDKb1ROWppHYv4WTttycy26Hd/GQqgn2gr3C
QWhNmHSthYEvN3UqHfFWMz8GNxlnJQLeY2gi0t71aHB8cPwuRfTi3qqhYC75IkZ7Ji31PW5QFs+W
y3F16FkF6TN6bSkdvcfVP1ewhosa3xcGbWnSCc9Sry0RVdIpJ2sMcvnMXNoN1KdtQSfRR0qYnxym
LjHSeGYkZK+FCO52SwNAmajevDT13cghBVAlF9dyUqhHOG6YSDRfEpHsmOhrHmrp/oWeBlR+EyU+
BJnbfykq7dJmybrsffW4D2C2IT9Pfgr1Wh2ksyW1roNIv5on2D7K5aecMDU7a7Ma2C90F8b8FaM8
MFPQsAXDWgb9vAwZDslVcjPfExx7NhPTovf12DItVt4TAzfk70CF/LEFAJ16CTJ3fCtvTT2vHUiw
Am+p/+UGOBipHlkYG9HrKK7vfjBbNVvy8mzsKU0EbLgSNHGkO7NNn7M1iEjk4Jw9weP+a1cLrALA
luysIb1kPJWdGNaRzDRQcfdO5cPNU6VOx4a9ulXWAjJYQAQhtrceiJQ1GsvqIW1bv6lb9ZK5Uw2J
7qRTZo8pOz0yrtVq7zG6+6m3kfocucjm3PNNHiHOwWeuaGjRqWK0E/logmvGvE5xbEzaWTFWwiLG
o2cqUXUDdYNupHWw4PlGVcyZfdw1KJpCQ711AMbqpxfhKjGK9PRDuvDJDuSHsuKH+6y1xvs8sbMI
G+K8acDu4NdMKfCMntjF0eckuG30Rq874YPuzASYISIIxDhI+mKL8IPIWHBt4J2JdXC5g5Xi+L+p
yuWux4sVujpVCBKZJXQrVwawP/w+vupJKHIy1PNFKvDXvg7P5e0b950ZiF6uB0419WEd4/I+TU6a
LDyOmMz+4VYTsCjeCNEM5eHnZaU0NjFUPQ8HSZYqPpUmRhMe3ECWI0NRboDj1+upAui2rdMSRIWM
ecuxwpjQ42B1X/35KnWwGsYFyvdTJsuxyaMhJuyhrYbl/T+/Khasdto7g+EZSR0K2TzVjT01Kvg3
7PRi3jFhz58nIdqbFhhwOfY5ci3k+OxsbeXJzCaGX/qBluNsgu3KNs+wuBwi+r8rI/OKbB36pfXD
iopTuWr6wksZn8YKlm55V2iKtFAQKSj+cGU113Hb2qt0BmQuiC/++g4kaNdTPpNWvWF+4fTCqSKf
s1T06qK8aBbm55GiIp69nlp6ywkWab44hixGY847cP7jvzDsoDgSO1VKg+puqb6YwrK5PpbKpqZ3
nCPyqJePx52Hw3ZPaubYjhgOHhs4gdVfdQZKttgzB64UQBiMpZtgSyh874vaEV9dfb7cAIaHqrm8
y+ot1kfplluM6mVbs2a/vJPRSjg/rbp7ImgybeD2REPN8vWwyFbjuOuOKRwstkocqhVDjKHo8YxG
X+1nvO8TFFoFlYJjmpMc2Fe6m9VYw1KRmCjNJqA4jXdY2cg86fptEdHuOeXaaphqUUc53k+gaGmp
zcCv3xf8MD/xbopMDpD82H8Lehc/Hcxs1E0vIGdwQj4vMZsEz89bm+gLQi9r2fEUD1DtpvgAP65N
lKBB3sHnkuc0QWfWqwyqhAxf+cjfryL02hRC+KC96iFbYhHTScugJ+g3SVIKqb+jrfdb6bp09vyU
ieiNp8xKahc6WxC++/uC1OrCDTksXAOwt3CIhaWvc0bBLTpPz6kr5dzPBZ4vXPAPcsSlzrJgx8GY
yRTOE/qiVdY9euIVNQAPjco7Y9vYnWJThgvhLiLORl8yG2mRC21RJNQFZfbTm6+0SHtmNiZiXbbH
Vs8ENc/qFteMXvb32L2QNPdHSUbUokcAWjNeSzDyG0UBVcnXTz1Sx52bnboHauYF/nyo83fEmBqP
g0zTRrjieL+Y369x4YQiniYhCH79/vBsglDdn4h2dIf+fca1WdCxs2ixrrKTPygEmurFGVOPaaJq
q6V6qpqsCus8z/CZ5cxECy5+HOciAeYDAc4ROxK3h6iO89/EpH3fUCHrzwIsQroJmiYl0ZgDulot
RhmKorn8WoC1almG0g4VMpu4Z3PO3Uu4L1lYMcqbqqTjZZIBSG1wICr9ti/HBrZQw2xMu2kJaF/v
qBOaZZQ3SvrGH/yUO6IG5X5zsH5C2fecauao7OW7EFrOjUxRD9zEgO9yl88pweBFR5CCVom38syy
8tm335d8dJ86D4HAELfGpIRk3iDm3vsVD7i9tH2a2X7CDL1aOUOvgjT67ty0rlSRDzXRi5bWaiCY
ijKlhqMRiEeJYF8sIKABryk1uQzj9Wiudjwqtb4vIMgvlaAgQD9TvLyeXw9jjkc/PmtWACcHVTUU
Cal9/PL80ke7kS1rbJZf9hiUwdGDerWBdphA8sXX5nUEgR7q1qIzxwoKtYYxQQB6+39Fb5/Ev07+
eYmTurrSb5YNzOa20BWNM5RRvO8M1/ufBMCF8Gfz7Hps4Mfmc4oX8LVGfQApXgwLxswinR8sOLzX
a5qO7WOoL8EmW9tXcRwW07vLeMr4zowAi/th/qr6DCq0SX0LCgLVcpHPQTSAoxXjwKSSbJh6BvBf
uK7vae7WyASw9tnsHP5vO9umIIzzUzF9EZmVCJj0UO+7DSi86aqONLCPPgJP2X0u2KPP2A49BSvM
hdSQVoHgQfFkI7GyBqoqlQ+XSAQKHff8IdjIa6bUgCdvCr7gf19hntmH6QGRso9XPK97sYoBWQ52
3ZEbb1lHSDVHxoqq4fQ0o45lDyaOB5vSHqHFUtH+z07N3E9McUecxNIx9V9w1whNLLEt6Os6tr3M
uE3u4c9sV7J3+G/F+GuIcBmDtvQWeWvn79omU7rxxMu+t0kHWRch2iLTrA06Nefu2sJJPyNG4ySM
mBBmVhs7kyy2agZB7037rlTgH4PreZMnhOPC2kQVeTGxLkrgX5byRojIAwKOL+/BY0pl/Pw7DNN0
/z9OwojqhWWMvvnuUvz7xax9d2U3J/KiSI0LTrrFSM/1wP3uCuoCMky/p40Xfr9jAZyYiUVwQGou
2OpniqKgZ6XyB2sUkQG9XMHB9X48ssrUX1v6hdhehJ15GhW4rxDhQn7PX7g6Phz9hRAIX7CX12bx
SQWjd7tcrjg+t4qMGfc7/UsGor9k8tuahyCZzyKiii6fqzNkum3eg9maPG9U9T5ZlLxh+aPext8C
H6uTsfJUZh4xNvhxQK8yS/xOrPBTZXPcUlmF8tuDniDGhNuWR9ckRN/3L1RCVYnybJ36dzeFT4Ia
iR38ccgfd/3f0+fEBNWNogmHB3CjJF4B4Obt2r+jiVNBv45Xg3iDUit2nw+kCfQynJ5ezW5GW0CZ
8CTTW0I3nIvA803X1aTs/DAslI27fk7vY/XXEx4Z8+NAVrnSOwJjbts5/hOWUfScCdmdGejmm+sy
CK6N+4xJEJ49gTP/EWTnPOTvoBmhpT5JZgADQzNrYO2m/9rTH3hmbACarjO3ir1cqjRgwymKREGq
XCf0NSbntm5cyqsRJJSe+S4HWClzC3DCHl2OTqgD4ix8EoJBoQgHTkcUpldvTdCdPz06IPCwQr2K
bCXU5WzVqXBA83Igy9BhGqyYp/Jd6Vyx/ks8HJCGNjzKDBydbKHHAG+YpqdGByFTWLn4BXBbtdYe
FhGiZvM2KheBkjscx/m8qXdn9eyBaOUZeOxUSjlXJKjx4mdpGD+OJE2rUAY+yGcO+G9WRUpF0zeT
PK6GVkynR8VWDsEwI3QvAAhiFOY2EDWllh/iq1B0YUwLQKLUZhyhIvOGInp5pp5fqp/I74tSI3ZE
LA5eUgq6K+bP71mzwkvO1H8zlMYiqlbr3x2+S3iH8KYrIB05sLBFkdx7VonIkbIimxOwAbtxpdhm
rMhd4q6XJKVunvV44384TXZI5BLMFBytP7nc5s/t1v+22EkDdnbv7B75hEdxmjm/JfhPVVjAhFG+
GjO77HJ8xYdCotI2qBQ3P6e9uLnx6RD0fchOKoZdRlDUNYnyjqj5ny5okFj7ECXQHAy25hGhNEK4
ToMmoH0Z/RwEPBahsQmY29vUxdj7JzyG50aZl6Y1udH6+snjjLRBp6wBy9bUe2JdDek9xEkPC69e
H11yUVcgfplrSg0mKwkH1J8J0o8NvBf7PoLulZgBCt6aX2P812lf6SOzXEP7KSGiEyE8rB7ZShGE
ZzLO2q5OD01MxCsVD12ESuix4TW+2nmjrc4t24tlW6CtXaPi/ocgyvMeU+uf9FqqCLo0kZNRu5XM
OqO21J+RDsaF/SEnEtAMXDDanWHIhyu7NXwn+XY0lxHabihDkEuaA3bMtLIBGTuwVk5OP7/OEi3u
EXbo11Oq6MBLhVfIsupRUFZ0WkjOQF4nLsHREwzMDa5kcMp+u9sW46pSM3vcb30JG3zlhaIr0vhz
61Nlcu66z/uqrdvAYs8T2UNv4zSZWvvF60KpWzOOIxotLr3lsaAGWGww0qVQQxNv7HHanR2fDjZ0
ttFGZwhC65a6CMWfGszcX9SGruvnjud+renqmz3BSbgKTPtsJnGyhkKmdw5+1AcJKdrEeJt91V8k
bWyNCgSQrQFncH87NaP8EU11Ig2qosHgMwst2jPlkYnXA3BzO0ltINE6zpCZ5Mk14Ew0GW6gj0cH
6ub1HAvqMBZfb9MMSJ6jtQ7OnTqylMS9Euhm1nq6dAPiSc3WotdVSF7zX+iTN88R6uvXMvOAkhD7
84clwf3MwfOSH0YB5wm0x0eAIe9D5HtUAEiUtnpwskB+0Hz626RgyQ62YTVAYxzaAMJc/EMTtttg
vd1oXzASvRQytQ/v2z7n0rMLIrHsnLWAGxqppvcKgy1DiaKuoEFlrY6PZrNnPz4V+zukLoJIa8XF
7uAxxoXLjZpnpNIgb4nWkh5/xWTmbN+nbt7w9kvgSjW64aw1MhL3EfiRNDQKWnLegGehVmGy3Mao
uaaw4lX48dnMXr0Y1Q1zbyCRIwavbn1G6hEdQuk6l8ow00fVhTDfFkpDyvSa8VHjFwGCdDhwWRMQ
76rDsfXQya4yw0FQ/7OM3pszKdHM3G2tYTeJNBIIBf3JXGZFMTo/zI/wOEO1kA6K2AZAN7bB6ZCy
0z3nj4BPuykNXA3Fs+EHeQ5JgLVZpf70WPA8aVn/1625K8ntga7wdKEN7bOhd+wmuP8tUZPf7Jgf
yLBQTenoaF+/v4LankJ/pYnXqy4vau3vAWOn9lCcP5VyyOoI0Led9iMgyH55LX8Pou/FvV3kMN17
kzD0gsiA2wd0ZZ/zmUDj0Ey2HYFh+CqeO8N3C9WGW28HhKMgQuXfbJMi9CNnS3B65bUB6PzLTTut
Bt0uuZYb8U+NvKhif0pB/fIc1Lck4U7f14kQ0AylUalyk4y+/jemqf+o9dZ/kLSdWSAiJ/vEBd5m
Kgf/YRw5vSVVQEAFayIYG2xFTlibJzAWgsMbMa0krv0ylA7MoDkm6Lyn6npm6PoxV9or7v00txcf
JuqmF105b1tqFDW7KEN9IoxeYlxqNUqdDUw/hNwN9E11v3ngBd5qvUHibdRQSAkJeMZgbCF/T7+/
R1pnYiYBrwSIzTwalQLEigP8HMmiEOGW2/A80KzWeKqGW/BGQgVxnx6MHzyko4qKpmTd97zaqQ3a
lFW/FWHLeILMNi2VsOidP0iKqFOJ+fq2kbC4z4T76OZqYfq0Y1wmjxqzSwCTcXckEPYOi/nBocf5
3r7jPrNdQGPrbjVamKBMmuhPHgnFDqlnnMUt2+blYqQO/xw9FyBrs/OKlP8hWORhr2PXVtvYxJKF
S3mpub35fhgzd3c8VryeXBeSdu1g8Z/nIrwjWO0XFfYsmsH+TiV/eOJuwyWOcs4Wd9vGzslgmnb8
u1fzSlD+Y9LlPYH8U5xlSiQ6CtWmkP/LjwH2XDpeeWZBJAeeJphML+98yqYTxFTfQ2tFfGAlVxOT
u+sZiUdt81uMxGu5AhfdsU3ys7HoYmd0E2yqSGdgud+RmCBDOQnn2fhup2YyBZTKAebjoL1zMg/e
5QSwVNflCHCwELRdE6GkMxrbU0WewbrT5F23z2t/+L/OqWEStzuttXL++wN/ZxddNVjwx34Xz7l2
3SM6VqnHbz+dUKtP+Qirq6ybZ1Y7sZcdYi1uo6+Ot866nZHJFVYqPjX1M7UoBUgUT2sBp6y8fYNJ
4eShFCBMLq0wH4u/LXK2+5LoO0Otg9AMjdqiFPRS/9Sj7Btatn2HDSCbNsVBtWdCoGz1xgnG4z32
418dM105EQt/cOC5QtZGJ73Hc/BJcGzfjUhWEgQGhWlaNy/5HnbaiUuVB0LuGre9a2lvUSMMv7ZD
dJuN7bV76MPlzyS1FvMXEBE+4NOWtdOhhn9ypZQhS/0ktv9zg82wXKU85f7rmmkYcF9ubF4296bC
PNTUZe+ejoKJOYHFbEUru6KCyAey7E97NrbAIx2I0z+eBjM1fpI4CKIJC9h23x/wzskU9VUwXXxF
YR1aq7+OJXMAf77dm+x5E3BLSxtKGXhUmk7AclkCyziST89qmXEX1K5PoKvFDIN9EJJVAVlSWDlE
j/34hrSPXmI48NIFdEtQjAOShzsF/LdU67Eo9FxBc/NpPw1c9tWx25aKwltt8gY7SRlxhVdKyexV
hv3XKeV7LCZ3l2VpvT8qjWGW3sJAKbwb3G4mk9FuGrQA0HQXYh/Kfnjb9fTUeS7yMNaVTzEahQZn
NLeWOXRS5eRmeczqM97IyENcfxrixDeUUv9HNy61Z4KmVkSUIypSTuzDgut/8ONM3WI6X+nJJ+/f
HntS0Nv09UWvSJgm78Z0SCArD3lXB/XoIyK6DhLx9JvwKEDz7LqpPuTyE9jtJmMth2PYd3bHvPAE
Hwt95MPp02CbmYhFM5qtkf7ddW/V0e4sbxtnvbUOponIKDwDMtJriOcDAc3LPUzrYIdTPu9Af7iM
W5gHOu8XTrdqJ+8V0xLPou28gT8FilDYbbqOf73IwEaDkU5hsy+2Z6V0fTMLJN6zl5hAXCjt+zoS
cJEEj6Ad3UcRAjzbXPonFVsW3ViCBKWokxfXCGt3MtAGvdWRa9u3UldD4MfbZFC7k8Zc50iW58ko
l9hHKQUvuOvmIn51ZCtH61qK20xbQNd5AdNXud/XF7UBAgkU7l8aXqR+362c7ColT3K2U4rjKmkA
jT59sKc9qDxHRBRkp1dbb2f71hXHHlTyBu0y8pP9N++78RyckvqLiiD6oi8hKoYU/C7SUpON8N6w
GJ2QG6eIe/GwT7I8bjN45MZ0WYVv54dsPx0B0VhROTvsck2NoPECRX9cfxrpO44gF6H8pUimYCpW
F6D190jNF23+SDgtY1dUbW5OpKXTsDbymkR8WhDvO63bneCT/RrFtSWK/nxbq87Hfy3Q8sAwshOD
5fZrZligfy9I2qP+3mBbrrgedrWjj7y6/91jCSiCmfoTDO9X0J1LEK2Qpk15vwDuvJ93AV+2hDch
Xf/mtbiheNDOUHW+lqPW0KlV9PQNpS5f3zDM8aJL2agAgS1VUtPcUGzu+y5+V597CuWn9F1CSagp
J2t59Tv9O5VXt6rJ6dgrS8vaLAUPYOYpOVd9fwQmA4K4N0tUm15VGp5YDrNBDDAFYlA+IZvLP2km
0sEUQr0VCVXDkchAbRv4s4Fpu/vy9Kx8ycOz+zJWt9FR63pVDlQDOT8jpHpWn3OVRCmLVbNTu4M1
mVbAYVNmMPe7K7GITzaZLxcEBzVnh4EsHSeKKG1kRCuPHtVsO3jIUsEG4zImsVuhSoVHadGYMfIp
pr54vP1XLtyWqXHHMU6FE3EseHdOQM9OkOH3B//00xJdrjCWzp1gau2O9uDkoi/UVNlPVQEfPDBU
KK7j8bxsUKdd6Pdyt5WkovQJhwWV+Nq8Qbkv2zVasXIzUA8L6iaHPejrDTHI35L3z6/06FS8X1xj
5Ixe2b7HIZCRoGSbVp7E37cbPGoywIuL5xiLqAD4zJjgp4bXprqaSfgE2JqaH7XQFLBArbsc7k1i
YJvemgAgLE5WhV8SmpWYviuCH3JEA+4/LCRVSIQnrhi6hVQPQyEN8FdJ80DTBW0/2KFQ7VKdy16j
0RyZxJQmfhwv09r5+2L6F4ByL5thgfniT+RBE2XlIwbC/Q/x9tMjymn1nH3HurpIzZX5DXmqeUf+
29s2XGVOa56/fHG7oaRyTKcJeaQcbN4vet1rzXVAfVONAZ9S4TUqg68gN0w/skTrkW75+zQ8gHti
mNXzfyrPG77CFNmUeT3tJV6alW+A+7YVT4pdiZ4hgTQepG+sSxDee0Zdiv6SARrcP82MDp97+abF
2T5fjTK8qjNijmKUUbK/3BBxjMeXzVVJ3sImF8ZFBpldzgdmiR9YgjDverwkY4bzi2759nEZAYmD
R4sA7hdMfXrbOkRng6UoCDZc8TG7zgJSGOpTkC77eJn/Hjz0zLkCrq4g4NypwQTjaPKFKZUCuqC2
HmqqYbj47kviy9jwFm7yXMqi2ysr1TkXivWWgrgW/FaFL/ym4R0I6wETn0bfHmjORMXha1UYF/qH
7WnzHAqZ5mjUdoQE2Yw3XT4LXAnG/6i0lJhjSHAaB09w72pNzNthgZeMeZvBWzXtDXMCO6aZCQNY
tPG0jkeVETmyiiAGjbx7uQPYJ8Ag5qobW/tjxnnYVJDLyZB2IDMibgEYi9XMgfLutzOXyMivI7ml
0XiFzN7rDxUtucSN89xjUuuAzawrURy65/qQjorUO+31IjQuTBuGBr+TV4+E4LCaiUGIPvvRWIcD
FYiHvxT4sFRrrQaCXz7OQBUCpz0z0FSI7Qt7K4cdEh1h4Mf99DYIE16sBvZmfK9iBSsF/MBNZies
95bqOVbBdck/3NbNL7bZ3mOYdb3/wdQ3rBtspuTTw4ZC64ugYR68bc+Sa3WIwzar/HrWJD3MdseZ
H/wzTiRre994juWUEsNTQLjBK1fglHMuQnljEhGPEEaWYsusMqNylClzyoCoZKICT694VLXtuw07
292goNgxlk7oo/seejNasq+Yl+0+VgDSU14AqvShbZP9FjZZSbViVOrUdgndjrJgCCgja/oM4lA+
6qnwugq6pElOpJ0VkndO4VmsrgziyT2ooPjZ+qtgm4h/xCm5AUiSBysC0yIb2Z7gQBL48fw2J5OE
pv+xCxKcPRm+PhnToKB7ptcpz+7PQI33A7XqQD/JxtFZqm60hAYX0KnGag8UB0u2cjdKD9CN0gS1
yLii+ESVmyg/du0vzCJUt2nUmFC+9RXLnPKe4vc3QyoYXLe9Cqa2FeLtTgc98bNXHmyw6YjS/CrV
YjAsh05izn1d0jkJ1Nj1UalD/VGzBlhFsq0Iow3h8kPkcgzMaD8NyGN43gR+WdjtJaglZT/evpvl
AoR0lsNF/wHZbyA9XRAdAzzd8aejpSa1yX/eqkqWXqem2rmDPIsNmYI0FyUWaONjjWwoxTgoACj+
yRXAvdaGs6DUt+b3OQ6Fgg1ELNx7JKgfvqH8ahcOpg/8hPMbUhGCIdbMoDuZZeGBDRV5l8VRArll
xHlvuVwhAS6Jg9fIu6nJaAz9kJV6hu11jeCV/3+jIcBco+u9TIfD7CuRCU56P8YBAQidS7rLyrfv
VRTegyuPdQ7hi6tM1E5VWL1GgmNulei9vh7vxhRSZNFw0NZ/R/cGneLPUXTbU0c8yVadJufqebNY
54VFOjfM/2ZY1S9r17PqmxMLxA3msPDQrTltC1DgsHwXjPgx9tVyiVndo0wccUiPeMXAmeBQdca3
Lv8HeRFtkZElur0HOG6NZwn0wM6q8vyHuymF+FGrR/g2Xhh59x1neTh8iISx52tvnfYN8bW+Goj6
5mkbIvvzp9FL139QTgSWBuj4DjbKJVOdSVaToDBBH5f34MwEw6KCkK9FIZUjfMdzwwuwDS0t4OzG
R90nAPu+moPt/K+DUwYI/thoolgB9Gh63rjyu6B4/Im3KR5ERFQpOxdE4BNR9h+Hi5+kUtxIn4w6
h7VZfXMMCqcyEayw161IikrjH1N0/2X8sRgQFAvyn8Nyp9e/sm8Vr19nyAAbEEQxoEzN2wtNTnwM
YkZNjc4YZq/qJqfaKaCPHv/tYkA4PiVI0cna3xrpOpixD2Qzk+5+eH0jzQktKagp4eSQYE/SCY6L
cghwP/KYONLRhOK6xGrQs35jhZVH0DjF6EpswZ8RTuwLkgqu9U3NO3F9p5hySL323qxv4sCCG4FQ
ZOl9pEsY8BgfBSEAkBwINoBxztYSG789JIapxmjKzka6KvOpdyqeJCy7HlDU1zu4rz9CpTLf82Ns
EUmNhjIs0rS6y1VMLeSbiQQj+iKk9RQUD+IyjG8WPcFIZXsIOrYAJ7a5oXUJV7fjb27FfSuC4kkI
RLNoT9GfuiIFdnaaCfgnb+tUDzNQsHITkSnY8/hFpWBeX8wHeQLxsDVW60N5qEEt+1BLPqdthVeX
wdav0f+ZgPmFYPXZ8wMArEaXLoXH0sI3G5DD2LbRVwMRiEFHuNgDixP4Y1UwY8xRFCyUD0ACdb3q
TciYq48BOTYXZaR3VBMRN0blP9nVGQJQlb+h1yqtbC2eeEIzsLNGQxeyzHWV139Cc4YO7YRi2v0Y
cf5Ky6v0VGDQyZe15aN4wq8vTb8S6Y9jGZCiu6a/UDnnVBizpb7kd2BhR3u8fVi053I69123KYtY
WriQUWAoNeL9X53bHlSzCJHqzbhNpVjP1/Rf+1HP+vR8phC2XWJxrRg/1ZU6wChJWUIl6pJ5fuYV
/j4dQlO2tf53LbeN7iWP1Q0r6UHjZEMD07L0NVblKj8+ZpfO80ed7linwW2sWeqn72ylo9u5GS9b
THDcVxXkaYDRbZMy3AHxyyTFi3CGhApyvaUOdXJHi2hazpnDjhuSRVDFGUTzv1KSdR4NjxZkgXRb
iOoMUAfIhpn1LjiwFWXSOG/9U8bWnITb6P7QuHgQ88sWM/6naX2Pfrns0u7BKWb9PhF6j/YYcmMR
6nK0HXoP0blmJq/p8S2pYPaYlEx0cjfrlT2lKAnWoOS2MP7Kt0xG8l5wHVCSPpO7w2nkU/zQrLrX
+yneneXJ0WNM7/5iwPowfjfQRwkQpJhtswGnuFTmws2tVWrm/tGzqRkiSW6cRTIWhXg6U+Km1njn
NbdYpAbStSj9ILyqmC9U18+HGDrdgbriw/fK0LndFb6InVu8KYbEYpP+S39Fh/i0t1ty+zOH3LJg
nwo3F73ZNwvkCuDwdkLsI5/pPg6NvWbaFFp/bvkmcvbWj7CLVT9tX0LTik5X4kn2aptNEjnGfc2z
lUTK2DzmqFkSqcYVVyf0su7TuVdEEvgdwdQZ+n5BaLzgZtc4vI+B+NRc8Q6puECEIHoK9hjFuI/F
O9MAb7khzJHuC9LwPTqSfuXXN/i8tgOuNAip8skpBiRrJ5opDcvUgdK5/J/NNupgONsFMsbGw4bz
YVIPSNw908YuaLzlhqUmxsiFDFh2b4zeF6simzdhxdZOcG6nIUw97IEa1wwqNS+u0wgcZrioczca
eO2mVaILOdsMZniybGO7qJ2yLMx20V+zCFtNjqwi/Kern1CY7oLZS90UEf95OMOpblTR2qRNCbFA
qQ4WSY3A7LVlacdocSHEtfde7Qd1t+KxgCDH6GWDHEP5JnEBLLVJvGP60PRWuiBtyQjfog0PT7Wx
eAQawVHn9RVRMIsIYn/eCFOuX6q+LalzwY5yELUnATV6/ZeEBcFrJzdGmpawFd2mjZlE5HTG71sV
CGbvQTnHaIEaIjS0svSY53xfvxsk+06B2QpU7KOYQ6sMMpudjVQsA7u2zL4hfbcMItam/3QCtmvO
ZLyVT/YCWezWd9AZvkOf1jFAgmRGHSd6vtFDVjdZXc9EpU5c6zfnUpdflvQJr1E/YZnkxkwHujbb
oGj95enbiVPH8c2FFOaOCpkqfpHNEi56Kyg+Trm9ousToJm6t6KRicgzSfV/Tn1UVDy3uyLWTuFC
xXK+HiTHGv+SprCi9PgG+Jw/mJ4q1RwljFIgHsArxy1ZqPAYC9dqGcojKuA5RToDfgUGyOINGm6O
EMueFGf6vPXxZEaMJRingQTPYdG1JzyTau50VCI1KRMt0/gdbYzO7BQyNsaJG/X9Gu3Fea0Rfyj8
FfgPoi1WHJS5olrYvLwnCVaM4YMGJzMZB5vMMl39XXz4+2ABr5YOPHbFiLUPOTLnfQXeSBbe8T/D
zaXafAMG9AxEBaaEmie78SkWDW2RkozPQEy3PnJShZ7owBOa5vz/8RfV9XwIKTLSuK6qINXCDazl
u5KGCIXJSUXnJ4PcoGCa08uCJThvkwui7zlDo6BxvNSoknOpIlvrjLX7LZ7tRIq1GJu8J3RXj4wk
Gl2H83guFdDPFzlP6WChp83K71cdCfnDYIlatpz/zWhDdSBurLoF9ggFuDPGy/8mLrLVIvhU98zQ
LiHMSY0PzJVdFwQPdkyBujZ9mwwKtCtX6mZqh7BnP8Ds/1FmN1jrNPt+dyBIXUqdYWzvtZQmBh5J
2J+ZpD7DS3WihG7ZaSV2WevOqh5yrMzJBX9o/G9y3lwRd8hk86IrvuVpxkyQXrC8B2KpmOrBx1us
R0c6cTAVzdP+M9JSb9jnt8mRAAZ79f9joH7NoqErqs1PzzXM7vz5EygpjuaQKngtUeq6u3UCW5Ne
AQWmGkaJ5ej9QVua7hHzMe3rAMhWWkC9TUiiAKpJs4W/rWS/Ul2FwovwsdXFrPz1JZoOuplA2Lu2
0UTv0vZZo2cYq8FvBPWCO/ObNJZ3gGCNZ5Wy4VwbGrSqjri7TxTAoNdcBl5P7/x6fars7bDnN9qx
UZcLyfLRBe9pUnh1zkEh4TqfPAJSpQJ8t2AFQoyCMiFHTF9RYlCwsf1lQHtkKXeIASlqF8UebMeA
0NAej+Vo5TekYmoAL5qTPPvWMYTDWuPLfah8eXnkdc9kVk+1rfjswwLbOROD4CQLTo3DaCypE6I3
6vjfXBzWdf2UKkHxSR2hAJPJJjWtZMy4/CkR9GWplZpSiztq2atlZgQk7EvjZOBpDr69w8x38OkT
+Pob7qZF856QE1KBG8dsFoQYLZhwhBeFzZ1k7sqLeREcb3vt/mcOo09HWc9WtToJkXqanVONcwzd
b+JjQamNB926++TA3+WnJ8yA+Hzh8S8QFwScMTE/L0HIU6M4k62D96+1gL/y+gK9St6WNGXDaRQI
OzMtB2cEiO+FcY+R0xsBAT0veesVTmA7s3Dj11k84m9xnrVjULhIY7rAEPg0ztdQ8bs16pGB1X6j
ASXKxjbY05yheK0X6bPfSelNOH3NVoQXH39i+83HEpAX0u0dcASmBvYNX5qWMqc/jh6tRVLiBgN9
WdfvKWcpHuamOEE23vHXD1wI1NZ4FjPNXboSOROLTmdGl4HTVkw2pIBG33ujj1EzpTYZ2MuulTxi
b3cQ3aag8xxkNO1o007Ur15VUkvxcMIDH3NsUbs5rC6L8L5muKp/LQ9N+lal26TtoyQGHXNY3NVW
4d3m7rFX49fxAUwenXY50j5R9T1oWSsCS7Tn0L4bS+Pk62c+JH0uQyEwI/33d4fPOANwI5mye19+
jxVY4uiVCFclbBdFjzDbLHuJenN8CQU68It+rL8T8WaA5Z2eotlE6h0hMtO3O2+gIHDkJ+3ZKlxn
k8NmUqxvTEnm9Ep99WLWvUdWxaN/NI54oKhLwIYSnOqqikkwo+SsErrhE9GyMF7mX3R5MSj5lt6V
mW1v3MK6MVj/CAu9tvy506N3X//FXFCQwMB2LsgVhfgr5xgR7FGXsJIAr0PK0mnmE75Qn3wXeLpL
LtH6OhswTRipKS8a7ATh0bfRwLyquJtUFfayut7adjms/fcN0UbgaBfoPP8PAWvimr6/YHNr7wWr
v2zectD4GJmlvgf0xedTUDu1iNcmuRUdtJ1RcIPbBzhxUiKXdPrW6VsGKc5JkGiYlms8p1aicBIF
hyNAXYsDSpq94iltGHyyQ1296g0/uSxsaQE8kjF6EsDwJw6dWZUWKaNTy8CahafHJlKVUXI7fSY3
/HsyHQlXhdmW8rTY9p+QZPX9UJRutYSdMx5+1eZ+mfhE5QsaX0nFLmeq9K+6nHKoXux+hMaQPVzt
yp4n7VYfFUkpeRY00cYObI/1ntVu2cqVpquvSgc+lOuOqjrvG/f4qL/RADpUL+6w0JMbmNoz9n0m
VPGBRNgU5BnMBWaNvqA+hpbV4TO9Cjy0LVA5BUCvHXyAIzAZu3lmPgu8AEDrcvtLJajbm8PjGwbc
/39agRIlUpOd0bcZFfEgVDf4m1Yxox+qnYcgdyT0cE+ZxnbVviCIx+zxfmnoDhtM3ZeewC5oFldZ
FUSgO0pA5BVjbWVO/7KfRiPL08eTUBycNDWOhOtnEIzIBiDnwlQGrXit23j16EOKLCRTpmPyb9U8
I7sKR+PcAeumqEI/6RGF8zf8CWBom/ddv3leIdap7H0X/6ATdiImAeIQckHs4ZzU+04Q4Iq3Qor+
gszKWrx6r+E3SBVGlu2seIUWvwjc9aVh6c9lCmSf8tdmZi4WccK7U9g4W9q/oj8RQ1tmmGGN5bHI
QV9zrTvsWz+z3NnoFLE24nFaBHpo/b0uBeOtcY88FHpRhLutPSexhGjyK6fJMFjiwrzBqpoMeZhC
soIxK4wiHcg8xkdzXqNTz3LNO7aOtXKKQdCjvkVcZbvQAKKuZ145tPwANhPQvhVjogvclsC5pqus
0r8hwDAJc31VIGieg8XjZ9O3Q87MM1KvT/2vVEoaT9iqFdpNWF/xbK9wSsEwc7ElJnWZoT6WpM0G
DdN2EZGCgk+5OFBOJmA4GbdPBMWS+X4yQfpIMXjfhGAzoeXrR2Va3sa9xRr/7uFV9KR/ezX13I8b
8mubzswYAqSPLTbQKxDNH46174iVfT8TK6Z25yO1Wax0+Buds5jWX606UuY9CFgeXE/g3W+dCX8d
2pjLurIZdnTpD0A3+h3LA0mwWvLqN7z+3wv9FnXRjtHWhBDfsWA9vUSgie0UPu4tlRx9jqCRzE3V
tOzoJphJXT0eFYBLaorp3P70fl/mzbK02J6crBhs8qfEoMgB66cb9U/+QJ0lZlyPgpumlR5YkK46
3OhnfiPQIDmjBddZDQxGEQmajhHOunON6y/qxpwR0RFpDK9IvtmK/97ZkH2TfdnPxMW2y+zgX2MK
Ub7aKBU8LReOWntvkkQxm5ywM3Rs7318tnFyLoJ/9PZtVRAmEaiH4dxEpvvC2oIFZB2ocdXbtEGM
HwWmxVk/cxpYRQYhGjHy0DpEBVS8gNevysQO31EFvWg5GiKGCWWfU6vnCdu9nOQg0V99FtICq1Nh
j7QeK1yJm3nAeQ5pwgu+PQv4EDCP0bwJbh7FKwPnlz7gaNmCzSJgpOhXGzuo58zJKCKbERs4mK8y
EU04+8nQ4U/BW21gNjwkVW3NNwk4hoPTxW///P++UwyJb5ZQNJk7P+6UiCYL0zZ9BtLrbZqbyZR8
fPEdsAKDEld/STNdHuevmY3lJKSiFzmc/AgMZ7dmU7Z3fhIarT6eD4xV+3uQxti3LvT5X9jHv2VD
NPq5JACYoENSscb+Akpi0S6Kr98qpgxv+cYiWGS6M1HRC8oOlkb6mKtPM4sk5F+2waBaUrcAYU/u
Ckx8pizW0z6XncV9yIQoRTgdRprs2Q2raWev5Vu/tyKEPrLtPB4qp4xgcxdrwoDdGPlP97FbCsKX
o3ofYNU/YwxDDYQ0gOjvVPOI0iTTSYwpmHbxfcPgASKbnQMNaL3VMur4tSJN4FpevT6UgFuANYbU
uK8zhNnILLQyt0z/1Vxs0Uk64XL3YQO96Gn+M4rxT98nFjW2iL1h2+drtQQJ7hbNisU+HbRqrkdd
o6S/X1UtDdQGJ6tU3rqD/e+cNDNAYrn7Oq+F6cRxvCF6q8SQYDGitqqm6TuFz6Yr99uy0K9MEno3
jPklkQr6p35ABKHm7phO4p+2F7VskdgV03nK2EdMv4TEqBFLDVm0f1k+KN8sWD2mRS+y0N1QWvn0
tN35sZ/Cbw5SYx8QGVy5GWTsK5x+6HgYJYdrDaAm976fZY/pmPABJlG+61J/hu+hNos3hNydC+q3
NPJInObGeGefJ1UBWfC8fnAwCyZGHU0vcYTsT32mxComtb4MeR8gKkGPenEjwtTjNYGmv/5zitwy
LuhwH8gGI5/twneos9LQyHDRJ7RvpsIIz2kr4Ngfs1pgkUIJV7I3fleQos5H5/8xxvAATzpbfxsC
WZ+11kqY7YG/7CdX4zEH2J3McTvwoWrn0qlBji1Voq/Dt9jXV6YCs4zLNEVCtbkNCGfi2Qq6U26F
ts4U3nuDkq4fyOHrMprXKI+Jf3ZtM2Og1xQJMHRoq/G9tc+GmSAGPRQaGxV/b4Y6liX5d92je7PH
d4TR3hHSV6kaVafbdAEiLKto4gH3W4NI5mZ3wcOkdq23wPzxzFwDrS2DPJAB+0SeFKh+ExLRF8SS
l7Y3wOhoeBLCf+pRUZCN6pPZDrG1iNNmSs1Z69v8uIfX+7fhRORQF4eh1OmaKBo+aGgynrVY3M3f
8y68p6P3Mqo7nS03rXspQhww4MHC0ASKNyd80eql/vrGyh1qeqe6tdqzeO9UjvV95PvnMFnlv2Lv
/VcNKQypPncoE/LobjUbLmJWyn0R88VqoFRdZTs68r8u5sVDeV7h3yp2b8sMfZjoL5kYVTPxgA+U
dFibioEu6Ch/uEciJtjXU3yqbut1J6ysveHgHjmEhLetM3X143K2NStnhDv5Sw3Xv95gtYxrsDIS
+8smMllYvnWtdhSsPQFjQI1U6vwZBoGrgn9eE8z2gS+tyUjBDfeoe0TO4yN6IMmvXC8yiW/LkkBC
Q21XIviKksC9zlb0PWj0Noo+EuCc6Ca+WH7pPrbiPd588sNyRIo/E+lZfaAJoZTbiyCmj3rqoHBV
UCr0O9sHPwuQ1ZsU9UhAx4qOWxDq9Qk2ixLDjhf3H+b6KXVwAotHYyX/bDYVeC6HdQi4IGkhWARi
a2lVTUdDCg14jnu5V8znwzbguKKmxbueX7+7v7R0N6X626Iy3G2Wgn5eBi88FfGA/0UdkPXuyhrw
OxrhYdo4K8FBwZ0a8FBbm8L/UI+Uyjn8ngbjYbHKJ8/Ak168rz9+w27yadqdEP/GL+c7S2+f/Kae
tz9Qpe06BFcbu1GTV5t2tl2gIENih60RX8lUoWKxXBbjdupdPw24/BfNBiF9xmIMSxW33+oc0uFy
6rpMFtnN/ujTw9D2KEMgXF3xQqKWRB06+MeCwR97DNt5sP4NQ5pp5Mg9IJWbLARNDW4qqjrjYv4q
g97sXt5zW9fJuu4/0cFWWEo1OSJ3GaWw0t2V1mhX1fu/Q9etjA5aiT5lepC12cgkYEqNBpWE6fxZ
EGFOvpKktF4qkFd8n7iCeX72uLY2tFjeNfPyoyCaVFyc3V5jV548Ru0Z8z7JOar6kYMI/sBk0pI1
qVNkK+ONYYWSK1TpfkvCL/gKLX5Qe0BjGc/m7cAHSjnZLbU+Hoovvx79exbWeJVzfpqEtlvQHVph
WnDrpk29I2Z/qHKBswLAbSBmK9kHSVdgP/S//EpDZORXWf6DiAEvsZ1WIyneOkS0BcRzmzXhBzZl
HvN8KfusJZHbwcl346ssGyL/PCyDSfPXPF7ncv27v9KJZqUBNgbFp9w3/ESDRlByvspt066omeUB
bnie4p9axUbeheHe2Dq0yjggzUL+5jUd26BmmMxBg8ZcEuHKwMDtOFQiw0U/CN2eK+isTjiUJOH3
6uRHOoUFvpBX/q7jjne5lqRwBTIHWCuw5ajsBxs3yKcNX18DOSLHTpx+R1Z+3FgTM4e0mKH9q2fY
V73+/nKz80YN2A28CZwil0DxT9nMX26pV6B5SG+cUIdSmWDcuHzzRRHc6zUslduwQypWtX+uxiNr
EJV8ne8HpQnrtZsgYN6cNEg6DBbPqaAZrFCGn4uLflJef+mwfNvvSvsg0QtEz5DGjyPeGLKdwfp9
mQtp6K/6QIuybmKVe5G0G1+97cU03ncpzaxlreKwBGhvVItzYO4n6TWWA+bO69BDrfKCppI8AVpA
73f7DmkE9w2L6/HbBoMVvwYRDyNfy4zepCNyWl2jCg4TpOcnroBbYwvat/5/idfrgwkqrzHVC6zO
f/f0TRhz6RiV7kUCOGLxPhHiGvEuORwx12qwrYcpEwDs1L5L4YfQaiwqyAH0DLTQJ6kGKQlwTOUJ
fDUxVV69saJMRt0zhovqoGBcUeUeQchyW6W43fwP6FupWakCoVUYf0ujbZnwumTQK+y+ZURocpS8
y7Eul2VNNfayCW04w4l8MRYJ/5L+oqrtr9S2TFC+HpGtBaXZarR3dAcNQTxHlTv2POnOvF2fiyVl
SJjI4Apb7ygTyD/3h3RKHQHE5COxvhaFLMoeempzsvFY/+TJF8Yu9nLZXVcuanCjHDDI6LdM71pj
HX3IgIXxqd9XJvH9PFgy8c4tuwhdaowr+CRn01FtvcqVWvK/6IvAH3aYiLHaM7NB+HweXDtKXQqA
cc6ToWrrnxEhaRlbgpMl89cP6U0AOdDY+Ooua9+ij947JKa5qYBVGviEfEBSY2o6yijwRTKwpHtJ
U2q+jpJgmo5Coy0bHG79/gpF37zheB4RQSFIRQhxlqkvTvGOCCaADV8JAsyDrFvsvS1VeNtmTuPp
txlcUF6WeC1bTPfUvefHQC7obNPAZjxrj+nXTTqHkKsunLPNz9qr1aEXnnKf5aVPT2Spe1DAIDSc
Lusd56wj5oVbZTt/og7vvMyRPezrXo7vPsfn17FArkMr8jNYXtW7CxGbS8CrIPIdiv1dfKAqWrhS
22VDciC7dpJwGrxI6jOViKn5iTYomSihmHeWratTv6ckNj1bx21EsMii8LJ5NWhlRciZ+vtiZglR
IWRjpT+MfruypPm0PHn63Q1+kwEZw6uNczbdrZkRO74Vq7epGzxGlGY9Nvbj9FAQu8rebzZ/DRO9
gtd20D6B5Uw2VYCCGa8qhBBoGtIh6f3xymui9XWbgP8lolGZcCyedFiq9IYoY2mjQ0xXJx6BKZRg
CXgBLE3Hr0clRanch350u0+KjoC8gl/fFgIXoeIGWDLqXR+U+NFk9b+gNEV3ZvFxO9iL0BNAzLFh
Rj+9zLZretWw0yzRdlbAvLvGMvY1UT4iVNprwfo3nR1J1/jGJQ94FThK8s4Nb+Uy2tEbfYHlF7AK
q3UvM9xExAqGwfPiqAiwwclg7Tjc4DfCazJKLYx50/7WFZlmneBCo4PXPGnm3EwL49uZO9PrFukw
oD636tIC8ZYDhpzMBm88idXSL6JpmSSAT/3GF752uKZIs6dnuCjdHTHhEqY828jVoDLPgHWZGw6R
6q2qRgUYSfUvWA46f8T5Czjtnh15GKfXpkTapmEWB3RJo5JVRCxMNl8D6SFfbOyIQRig8O50jrQu
oN4o88It3hFbp5c0AsrYG+Na6mTFBlJMqkKCUF+ZbKPa0CIK1n9ZNeIWzF16GBpiMv5399naC474
I5y8hrDfTb7eYNTfa6POBj2CqCRnT4N6nNuWUSwc35dI0N6upAdT9wjPelj6Ka1KXmpapE6udyjl
33AkoG0Ai9H6YosGA8uUwtGqGA63RK4Scq8KRseZ/8Xn8IdNy1+Izr0+8gWmqmOE6Qk14nmJ1mPl
iQNOQTrbIbJTS5qtg3TC14hbOjep7pJLMSp4obaZd+BrlILiPZ6dF+XZLbfwLCaS+3/thu61vMEy
fKwimxOCKMjK4GvlmhRs1AjX7VvWcOM6mq1RJmLrxt9VNy2hMkct/BUI0zsXL3+yETPsfOINEtAU
pID85EgUoeCTL9JaQelu3xMpol7WRqVW0//EoOwIwGYHzvPuaLO7tv6W+fgv2jjbrHoma4bKM61v
ylyJVxGMqHJzr6kZFtVEukAN3Hspr17CSSGmIFE3pawpnyGD8VCpDvs854917lEHoY4miR7+A/wZ
VRi1Q9ziPEABZ4ls95CXcmHkM7MjjXwuumL+AGq2r0giQ1/GhcjEk4IDrtYXPWP6q6lbO753M5TK
ONuEoAIm8cbaUkIeIXVBdkGOY86N1umlcGJVSx5YQpvvPl2vchYcdRbtdVK6vlWrLBD6PLbbgLRW
Qz/JTTMPVhpjJUm5p4QFbmnIV3CZ7H/UBIyRdrh4IpiZoMxi3KdmDn5Tz0/ecmC5UFbH51c/5QpD
WLmF4i/Ql2ucXH8P0dnoBPEZmnNipNXPfMGyu2hKb/X8cTOkMQUrjyjyeVILt0VXdFRzaMbMk81s
iwRXlHRphYKCYm/76vPYAH9GeJr2d4ZqiT1Vjj59qXIDuaS1I0m72X/nZ7aUIRoGsUzB63eNgY3B
yPUQ2M08yOejhpfrrh7yKYIgaUG4Xzy5x55avawa0REAW15g94JUIQySX7zgDtIbjy/10DTfdv4Z
8DzEGSp5Y9OrQRA4Y+KtNJVFCqGkB1hc56xCYlZSn8TK7VNWvgF6sYebRUVZhih8SEbZsYfqyLHi
sxenicZ2xgu2hvPPkGmkG643vultvnpOWyLB5FHV/N1TF+/PBod7dTfN7pLOX7GgJhWXZQtSwwjM
jNPDZFrY8rgqLYNGcnGnAYwWo2wvlq6+9Y5Vp2ocCYDOzx+KlefNxE7wcSoFUOi6cUFc0Bd7+/vL
ABnMESi7WdbE3f/UNrNOkI3uIbQSqDXdyGW5tmB83SvNTSFapuHaItPepC9kN+Vej4I4+IX8NHCh
ZVDdRZh5smr/FETJEy9d9hnBS5cS58b6fGuT2VdbQQUSV8f9HT2Gv48Ntfe4peNrFea3QuYI/aWl
OwkKyLCyF7UrTb7XGrHTB/LRxLw+uUQN5hffjAF8Q/Zc4iB5EAbvCSVqWSaQfADUEL5ucWddXlWN
e3KBPJ0rNyLw0dUs3J7UiBJICkYe5OYrZCC+RxQXZHsuPQEqgpWD8+4fzzJo/570KY82vk+/qgZ6
un47rCavcuS14sm5jA2SNbPn3dy+BbE5TScFcV6SSS45ib4xbEgqies1VptcYlDefC75ErjND92X
od3aPz4cFWhd4EDktFZdxUuZrg0EeDLLz49x91cW/UZpADHcCI9VccWnNUVLenbICYIS7vhrILuy
i1M2MJ+zHZvI5auHBUFVTqNIhN1UBf2ALYZTXr90oZwaOfrhu+6mi48gudsbP6ymEc8OI69VUnW2
M2YKkPcO3FB4X8TnTePTN+tMf/Vz0j/vdAm9KFjvMexFDCfFhK+ytbFWlrD05lisBbo9t3kPbPg0
vSAOJOWccBnQCF6NvjIGZ4pHBnAyyekrboDqBQrdTlAk4ZjGpF/292dz3ryUmhHZ8iSidmrGdmXQ
9+w8R+LMBY4QyPCkd76xrcuh2WIZmpHFdDhiWiSqR8sdWA2SSF6UPItFLv/rT4/3rHWbJnkOcUVS
9V5Hm4t+XMn4jmrNghLj1aJEf4Qjn7Su86wEh9kymKJTtzo9fEp42Ri2ikdtWPDhYLtFFbWK/mjt
zxIVrjBvzwbcS5Xo6faewMU0KoqTwdfEeUYbyAL89214axv5PwHXSadGup8l9NBx2xTREP8uAJv1
OAgrDc5cpId+unJaMD+L4gUDK6N6ufPnId6emHIhTm4Gnu0YfFEc4mwsqgxEyD+MwwqIPj2YS1t9
tY792SwDeUEor5gebzTFj54Qbqib3OVsrIdhX58wH1p9LoremMAZDFSMu9BG3hOgFCC4TfHYbbcd
2JjKSWetltvIF5Ojf0WbvpqypRsEqu+CY2Qs1Tsu+LuwPvLWxGeJ3g3cMPyP0YB/a19UjM6psAmV
xtfsOMcjGh/emBptc5jYGxsvKLVDcrmJ1ttWTu955oFVGoKcIHTwnmfWj8FatA0l7qUHrYqk8LrQ
sne9CQOFR3pNGy1Cg31XiK+YyGXB/0OeFYip+RsTeV5Xz9QwBnbvKZOLhmhEQZeCcQHhqbU+PT8s
nnd+t/J08XCb/4WXTr6eV2FpL9tktksBEN58X1TU4IUH7DEylPpHUK+GQa5JQiFIM+Y1O9v5O/Is
lweQ5ZXw00mUoF23X0eOGUmwJ0IbC/sFT8C1ec6sfatdgz+AosuZ9TBNAPM06y1ofVgCevml0Jpe
jSKM9eU1UdIGZqNuEr/30ziFNatQbDYSR3zqnpMqMdpsaJ+o6LGp5bSisbvJZVuMJxxMDzMyvON5
hLlP0S9GsKqDV85CEoziBnGJvUdB5ebclp17HG6IqaVFsqSlkhzsUp856yBKp5bdb9hh0nYzTBQi
I3UMSL3ZM7sLOCy+BlVoxjSm2medl0B5XpD6IZ48745NHYkSXtNBh632sPu8pGy4DT3jMZpVTxlo
7OQnZUQhWfpABW+4NWAeeuRM1p8KcF9WvyzEPZs42DGmHwba9tzLSQ8yYxOntkj23nkU9E47pMA5
uRn4gDWDoHWqbtvKgT9SoZNg0SdnBViQ9Vwl9abZfwDABlJ9tdbVbDpcRKeZmTEWXQyO1Q1NxQJ3
DCFlzxPoBnxI5KsIiDsImSrX7pbu/iZtpZSKEpbavQkWm1iEwSvV2gSqxn6flCMEDySeRUdJDA8P
M3tNbcj1E8iU5tcIINl9of2d4rzvzUa+kxxTmrN6tgsW5Xioh7o90GS/U08S4KHXsZTrCCR+bCYr
J9Erz6ZKH9L55gU9FKfXNFEuPJ1uYDbLtfnrx9pP8QAsTmES9DG57Pc/wMKr+MH6xpyy/Y1fTlWp
oXOzeG44K0vow/27ik6VDlFJqnZXIHaTu2i7S4bfJH4uOzuHg1gZI31pxh9O5SkDFrPuZhEfgzyR
23wZS42mH2+NiBKljlPtSuMJ1ZCLv4unetVa/Zmlxxnngy7rjzzhJtiu1JJrr7RkCZMgHOrSfIup
GIFtwNxF7N/JF6clAS3G5I9l8YV5KJQTEkHtIlZrP9tiR4sGeQYZ4hVS7VBlzWB5VzIvXduDC5qn
cle7ybT6EpnGs1mNF2tNLoX14nIFDFj6keuZFGM3bIUDkd8AKOKXA4qiIL0/a+VOap0XnJFDEMRJ
lulv4s6dJ3xKQQXrjNs8BIO1Ogy/DJVBxVx8YDV69TaIw1Uqs114bCaV0eVOE2ZN6tlXVCxuV02z
vu2SFrRy8kmFMHHXt4b5a/wdOd3rcIH8+KOStRlTSpSq5YQvcCHfAYMslQRKPZQtFC0YAACLE1Rs
7C9gIXEJWbJ7q2gwn+HgdQlbWEqWWLBglvBRu5/shsFRWWLM4jnlfH6aTR5OL0Jq0NjtqqQXHydg
M0BV+bK0F3Scboe8aiFLVpD+ejjdL05Abl8WXQ1SumvwC06Ke1bAyCEgUxnNVW2jBkZhOJWNuHcB
X5PmI12y90XX6cftFk5Qyrs6R3LbjaCinRhAf38nbp8vGdNQ5zJPQYOFhJjrU4raVKM3iNs9G7G2
qnOSRtmgcEGqogMvhn2M7aL8944x7wnCy/RXc4iUv+f15hKXS0OxfuaFHrcyAvSTbLx5qrj3TrBT
HQBykwfIzaX2N8ZgBeadEQ0h5Whbu5wtNhF3P+WyeMS5g7yNsPQoDU9zHGVJZIMQKYU+vhR/1r2K
OGsKHM70FDNoA5iZD2nfrpiEtz9CMlO75n7dbC9dCxjdI30fVN4SSgHN9gqHC4LCfI3rgI6Dqz27
d6tPoMkWr2d7bp6wF0KZTbaaPbrbA2I0FiQtYqAbWGLz3lxBNPEHRhww6CydRhdW9bd69SDDs0JG
75NeMVFkLgf+GzWuAbpevMj0GzRrYpeOam+HA3EK7EDBqbDAzC2D11FIwaIm0ofw9+HHMKsJ9iHI
MtRO4dQ2HxPAZIQLsWmnbvY5Y/n2gLJGLUWhaGt0LMQ0rckey9Pp7+MokMBZ3kKZGNE777x4MyGk
KtD//me7O5eLbso5SZ7IwbPJwSziLUtjHyXjM5Dr4C4W7itF7mtcIeOvcXPZ1uc5aw+agmKzGtIh
IpK6VjSCrjUOdRa+pA5REO2Ilzh9vNO5tY3NgkbQDnGuu+EUuiFza2ERuMzmBtgHdszzjtk9l0wc
iFBMRhF1y5E/S7mgCnxUDQRbXOMtOyheoje9Em3wBPleAsH0Uh3TT6BCiL2C0sj+iU0TyQGlNRL2
SK9MWm25miOz0/6qAlHhmmyDB7oXH+ZcvYmSEnpgHm6RN8Dwi2Owfl7cTj84DoDqjXxpD5oaM63h
o7kM0kLhZXMHr2T9W2sE19b2CWrqyLc1SkGJkmEo2pS9F6nJHShomqir2gh0a0V8DPyWzMGkXpRH
8LGYTdBUEG22ckuxzntKOeLVl9X6UQF+Z8LOUB+HLhKNTpt6Rntrl0jLCf7h8YBASy4pJcWUpduY
4aG89AxPrD7BvnPcJa4yLxqK5mRbbpbKK5vrRuu2LEwLsPWmia72t6G+GwIJDhJXHCJmUBS0ErXs
L49uyUCytrqnNgGl7VYqRZNgOjmwVLjsYKkBaMfxrhVjv0zroCp8g88rGuWj0me7c3C9GAKbA9hh
8WDyBZwQ8189vj/M7MIaEwHv8iasv9YvbEmk2CjeCq5oszQ9MWu63XCXvYaEoP1O0YRXfWzeOL36
SaBFLASsKNCxuEwHkTyjGQMENofZa/1k6JkJodi7BJm8Yu6SLBfhYPQdINmwJAK6bfUxB0I7pKn7
wVV+XqypJFfTL2wESdgqqBIsyZFwB8EzMjFmTE7V3Lnzz/dx0q/8jYuOVsxhV/411M+2KAzKxR6F
N30uKAMSjXgwaYCpqfKj5bPFl9Gi1ZXfk3vsN0C+QHEfa6r3fgH30dx3tOhbKe0y9pJAEV6VpoVw
We1w26g5vAgu8xTbAcHP5/udbG+IJhz8AbLwvYTLC+FvgAjJQASebv5Xknmyy82fMM3yPBKSrwSe
fvhx4lWOJX5lKMtUY9l/WpAsydUcRuyNsHDTnJxfXHsOBWM+WTSAyIlGNbfJ/75LP5GTIUqE0q9y
Ku/QNRGH8ccW66m3Vm3C5ysqpk+BPfH/83rFsI7ThGno5qxcaj/4OruopHSDu4l7AtzMcsYJsLXv
PQ3sMeOvQM4ZwSHP5Dws12vmizTz0dimFgKddT4F0EFJqel61khWr5xNIqnVqySMD/Wix9NFELXP
JbmJCI5CssGrjMnW4B8PtnnV5oZTt7qGSZFLfzea/m5/4HUt3Y4ejrnfcnys+IQTde8uScw7kSds
UcZ054Dcyajs55Udt0KGHQb3D8GEKB90yV75YKa4QmstT1gPGGgr1IRKxmjrekED9RtiuaKmCIO9
AMf0TMio7xdLr+qZCFnOGKwG0TXVemqcAXTegQBX55h8DUwbkKzCSGZ6Y4Gh4wNbvPB56pkU/vQe
BXtcm5w/HWbowRb4C9dnejU3hnz2+DSh1daaNVfr8CZ3tdlVVCqrNF72IWBTdIWdXkuTV/0a1EWE
17O9JqPxGKm9J/gmKNvwnSr7rsl47w4LazCFwIq1aZq9pNZ6nZJabeEZD7VRaD+Uh1l3bvucQAwP
rqDHgCN+4rp8y+sUerqkb5VEjPKfhTrpa00WTXiZhyDM5+xPcG7UvfaxZQgeC1iOqALW165ADXjZ
aN1PNRzNDIgWg4B6ZYpABq1jlB6K8e579ZLlnLgObfMQK3RqQXlewXEozckhqJKR4Wz7fWIkRJuG
S9wYJolietxLEy6n6qvEzKYpsD6r9lJngot1FM5i8A0iOdF/Aw9R8vFtR4I0045BJ+1+cU3UXVJ3
5VQ6/qbJ0lNJwxen/fAqLQxF6l+JVfffTzPzvjd1OARyCNn5dmWyfnMS8RJDhHlifKzNZEnVF1M8
P96xbNaYhk7rQoCErQd4c2rbw4V2GXYx6ExUO/DHT7swYOP4+RYyCZ42x4FKwOrw3gfoFJJc580n
p7Wm6UaY+MBrmO4N3fS1rZ6zilt+2M5lB4YzeGGeB4jVNvvVr58X97jJAVXdQpQKWx/nanu06BTR
pwrUZYx0/cAqlN5PXwZo0VEFMCkTuuIDMlwwwKAiWNOj+4kDCdFn1Kv48JwC2wQHqs+FeAN09Qy9
o8x4AICqNKNFzG8AOx43JflhSbe9pKtGoNVtyFsavwwImcu4HSBDZZWMdElblKVshsy5oOQFb5j9
QkeXXuK8At/fpSp2Wz0pQEKPhHDljUXjxdlAkvHBr4l3tg5vQf+8N0FctDH9XsoD7lDpo5Y9GXn1
agZTdBfXnf3xJmXn/YdoogpTmWwairQ3ZTtNTe/+vScfNobk+PbyupdbRDVTGmNyp41Zs81ktRiV
QLJWCOI6SZkcvDQf+A9a6pl3RcAQ2h0gYmmB1jUwVR9zam6qbopzjLmxmc3TUZ8hTxTy0shzCC32
BrLlMARJv+U4vtJi5G0B+uDGYsKDjbvaeTJywHz3ZUVtSBSzvsHSC4JwLcsv4VJEJenE9bUesDGy
gG++sWsDoTRGMeOvsNaHy+dTauWCJURQJYCWHXwbEtTv4BmkpUTa/hFT7C2TIVOEZfJyM970ArN7
9qk8ojyRoR19P9EJNXIdb7bjaZt39bC8nKTYPiutGVVGa/uMzAPrcM8u/OBVdfmotXHZlfpvH86j
uyVktGPp+NS7JDNC8QiCI+uQDLK7wf4JzcP5TUVAXNMGHD/3WyXbuDxxwUWjlOq3YUgdibZBdhYU
8UnJ4tgwpWKoKizSxDGFOMDwINtruZPQvpe8dq4Iyb1DCwARF0pLgrCeKw7EujTjSnLXMmPCmhZ1
PzIiq8wi6ANIAoR6FasD6BMtWQOOYOYVuuiC8S1zN/cbSCaQMO1N++X2w2/1BOuGWReBAtL4q6v3
1WoACl+jV0jCnFivZmQkecYdgzvLzo5AOpHrIEBzVhWB8lMtw9yW+aNHeZmng34MTtuu7eTPnumb
2aHNrBpPxJ9D+y0x/ctKhbPBJApRUKPUvSsoKtFKtnmmXVkRK4qTADKphmUoWeiQiuQdF3WuBhRU
5iTzcmaeRc9qi1ikEkSxSaeZUEbaxqXUp37yRl217jxN90PSx0lc9unwRA1D4GlfTsPymfQpcD0K
1AB4Af0/+xRcTNioFWdxgxorKkqDMjjzLCP0FxIaNuXi9iBd/h7xVSw2AmGTTGaPpoxN1uq1n2uT
raQG5kugDVR9Jpa4OoO0lhjE51xyY6D63s0Zts75qx/VOgxQFznLsGxR1BvBOXhiJJ3AM4eDqj2s
0BEYQovzFQRldVmBVR3msfCvkkxGFcupuaz0tf0PO7fJRmEEUCTn2ClLyb7aHKGsXhBCXlA9Kf8w
loCSApLd/DdAkh6ELQ4VXQEoyGU5IAPDdIM9R8r6Prb7Dg5WVql15LqwcS/FyLT+Nnr2NUukR/x4
g1COSRaAh/rme0WITXwEBlUlFTEO8j1Qh+QS35GYrFEa/63uh+aHACclEGqw4lm0te8fBI6TIZ84
T7jzKPztrvDhBjzDh3XNa7cTRIj4MN8fQzPoncA1hw86rzGLi4pT6sRiblnkCmmAnUd2fl8SWcGp
citcbWda7OrtDGSCd87+sJDGLoSHGK3l5J8FvSzt3WgupiemlsV7NYTdYvQnGTeIno/StsFXcDI/
5fasN65SM0yJRq0MknsR5wpEdQVNu6aodCS5zb1AxsQ6oeZ6AZrxCKnX38HO/tNoPzqCBxnM9LSb
SacA6MzaNkwdxmmbyY6gDbq3VEclIpJP0U2kbcdoWCBNTWI0Xv2xEhOCZWA47PZY+rBh/SegWOCh
3N9aI5ks4FKBDHMgGX9ToqWTsbSSvaFvGViYRlcar5fMGLmPG08yT1wbwJwdCUp0hZg5S0Jp16/F
3Tf1mPFeiAU0TgH8sXsXyQonCOGJLMbHuDHDGHfWqkIGuOxmk8sL/3dHBSe3iZpYchlmvY/cSiXo
4OBW1eQ35nPtvTeVbHQmkXUvSXoA0IVg5UeBRVl7FV4PL/vJEZ84vbX0lziaUdsMwR3q5Cc3iywr
RQrWZh5U7cB5EcJ1TvsG1yNpImyLL2f1siXcO7zYlRufInJMtpYEdVv7WJE5rhaNSiLsO2Ih1i6E
gJ5nihSQbNxkY1Id4XbrFw4klz0ito+hnFAagtjJaweXOW6tGRhfAjKQIuJY6XP5oadBBI618zQ9
6fxvCcDdG/VZb4g2kVU+S39d1TtW5n2dNaHdqGL/3D71BTsyzebwxiZaMC+naeaTdX4gv3gRnIZW
4R6+JIs3nZ20KQg47eMbwub5iLcllxbf0OjdYRoVhgB6OK4+7H1SZlbBH/hTOSf0I8HXh8YzHydv
8se1xIS31I4fT2Oo6mNkfPPOh5Ee9TcNmTrj2+DYYHPqELfNVdixlSw5jxAO8WfspCsTSWfVyBpv
r+z/i9DBLMqOnrVhNkcSAsQstF/i470xtfHRif03tKhsFaNbVsgXNVHBvFfy09VHrwVcke6cHyOA
7n5Hb9VJoiywvneUuengWSfGvOrbrybnfJB30gUoXmkPGIL7nLh4Dkrz3sEmEd/IkZ7ZNpC56tjU
nQKlAkgkEc1/Uz5Wd5vMgEwv88VFRCwkvZAkDyCkqbHw0iWgaEzZrCWPPFW2GtVF1wVqgaxBxPv6
Tvf3qZCOW7Y4v/j/ZoWekoysTrGOayNqs6Ewwj7lWIqCbsGMbW85VFTUdtkOBjAyWNGTHX0TrY1V
DhypETKSryghZ2Ivn9GZkNenJpa1xk9rGEKeMkAi/7/aFc1ZIAVrg/G25nQi47qJEFKBGlLf5hJy
vITMsIFF1OVg+Gy9gyCWTzr72cWDxT82bKjiTU3hw4gesWsDx9IoSQuM69jMoqBOXswJAnCEFs/2
7dxBvGlNAnLLEWhkRSlN9L080NV0pE9SZ7quanQimt6u7RcGM68vAmSiwI8oKrHO4MECCcmuP51C
96esLdilTf7ghu7zSXY6Vvl0Pfdu4mo6/B7ccARFMuJO3jdvP7UBbN7J3/y30bmv4tuoCRDzljcQ
FUn3VYxcTzVAvT5/f+J5G/ApLGKNzuIZ2gEe7ClsJ5HJuSmQeWo0WwQ55rNHvbIk/4KI1WJ1yO76
cwryO2EWH3MC3fFEqqr1Qfzbqtrrn/0e0ZiflkfR1RjZlPibC8ePvrizZ32AB6fUY1cBVGtrUnPP
UxHGSPLzPp5CJlc7STcIMscbYRb3sNyn2DMgbOeQHcpohdSdhcUSZTZj7389gUzCrV1nl2Jt5t4r
B2wbg/yoyr/TCWSf6PD8oVjldKnWTH5Pb58mVsm6DBjWxjJHJUFctVzR4vGktDrpdjZ53tHJLEr6
5D6s1OJxof/kC/9DPbo2ZVqMlxto9u7BS2JlwbWTwKLIULzdXRI0jJf/YsihrnyTBEY0baMMGHrA
4o6NHd8P75ORoqR4Shz4IefHR3HdFZT7VWdU11V9mtCcuN5I7gINpmHusXkANUGV/VyDSDN3o7uC
rQfNsFKpfl1qlYPSmaBbgTEzYHQPxpG2T+O+IJyxPPYbUi7Ts7wPbtvR6RxpHCSI5SIlQyzCbVnZ
rUEdU/O56gsXW+CznVI9JLF6GFTIYLXtwBYldhPVFVlQXTtfoBgsoq/E6qnropMPCd79J4Uiuzpx
dMTRhXZchcgLUoS3SU/xTrYtpmtUglvsVl+2eqwvAhXs9LkBONNywQDmQtbX66xl+m6mIK6AClb3
dqBjePUj49N7oeC3qgGpZalsA0lZ5cQ8rDwv5jcNkWbDGjO8WvsSFCLkm7qnTz/AhwQS3ygNhye/
JOF+Ysd6wM9zajDLRty9hAlivQazIijeGNlOtHkfmXUwiJyhsHz2Na2AKhq7O2NjkJR7bnTdxer6
/vJR4eL6P1guf0UDQortQ8qSPgBYG/Cs61pSyNo3AGRmZggs+fMHimtnAr5Vw34F0JkqTtrHjoo+
Y6ofH+4z3YrJAXSeRFFx2hBtBpbxu76XXvty/ceUb9Ib1GGh3t6AbM6jdlGl0gCXml+RihYdPo1h
/ZVV1qvTdD7SeAMYKo3znRfgc2ICOI2H6N7t5baWlyUDf7dHYSvPrBdq0JLApGa5HV9ndZCUDiO3
HIgWo/qxDJYpz2aELIN25B/rPC7s3Nk5INF8yoZWc2JQjF9+gWm4A/MKxD8lBrXG7PzPzlbGLua0
1TUE4LH62C/9Ngy4oy5/FYqGzOIxMhDCah5rgoMNXdez9P6rQLGRWqYHTxSMd3wcf5ibgaJ9sWWH
4KDZ9T+9MiEHBCd6cKNfKZGQ6Cc5FBwTQ/tqPWhfTuL+TJpcDvRA/CSSFwSEFVf2ujS5eKFdzwDz
iQ0qY2m8Vv5ZOeyPMqzZy0X1mcPA3pP8FcEIApEdG05yf+CwShqYuh9lwKjv4JEKPAmmD9JvE196
sZILH8XBcE6KOBbq1isPgvKopmLrL9ZXss/q8bupxOv7ALBM25qvzy9Xkz+MXgB0tewZLROs68+t
YyLu5mb7LwXknZ407Oo8ngtR4rUa78EEBAprQeMlFomZ5ho//6/xcQrTytgt188SAjHRzViih62Y
zQJEb8oFIIIBDgYoJBMBI9beWj62cjZZT7BPn1YLje10CMyvxT8xJRYsqGoP0CMM7A6y05ChrNBv
e1waC8CYyOMkCKEcjYuG1t15vtSOC0xQdKZxoti54dCbFpe5+9gX7srHFs9eiTFPHB3cIKxVTlaN
oWlAZlClKDHbet1Qi1sFxe8kRywbNLdYSffpAGDbBDpPtdclHf/69KoqFjG0ieahulEK431AUUy6
wGufcj/Vlj1C66QlMEaBUBe1ygit/6h/l7eeb9iX9paq8Hf+V4hXTs0VhQcFkr2qurf3gsOoYdMG
9FaasrmBhRd9Bbki3oVJuOgTcz7Z2Qe/p+q6FnIquQj9I9i1F7uzetG1yGFEgEfGXA0bvo+X2Dnf
9Rr7VB0qrbZP6PWWt2ZHitLUSmUcEQkf7SJQmUnmHr8/QrIvxUK+kYVfp350JMaQLRxvbCRoEnb0
WxOAI+ZpO7ImI4uda8S3Inv1XFZWjvyjcXkqzJkZYbYp0o/5og+jYh2QG+auqfRqHjzkaCy1FGzY
etzjl3vjjWy7nOWY94vgX3PIHbxMy62cfc2qEV8lAQIuQazBHXo9qcAoSk8t+f8X4BE4vmxhi0ge
sk+JoS0HaUZtVS2EB70GwaRSlQrksqpLo9dIB+aqvt/2PWAI8VwnL7EGGgY3P4Ud6YRtl9wifFsB
KdV7WKqqysRP8f15fszHkb/aeRK3pmQASfe/VzDBpqg5bXYBVWECfsNL3rWQF/aQHlnUaZ8D1c7Q
1qe3NY0YUG5n44Hzwxpvf0cthnh78VMuSpe6PwO4yfj9chnAL+Uu9ZVIXzzyeCuTy2BUEOY5mU/V
kDNdCoQHKIQOv6Hk17ciiw8gENS+fpNaQM3uXjv8pB4nB3DK1DEq14PRcn7ymSMdeyVA4JaaXW16
XYo7TdjZnnEJrKCt1H6+pzpFLM+DY0aUEGsznfnB4gwFzQjSzT0/dHh4OLNzCjKjIpUdnwFocoHo
SXPt0DerZfuX/gmxi9xcR8VM0QqH9ZwJYc+ozZEzHWugaLqTxr571/A/gUR+P37QyxMqn8F6iWmh
MbBSa/WwNZodaLX7EqAHvpBHHDHhhYK0T7D6ZMSfBDSujKX3JVGi4/Q+MEA7+coH/pJk5ej8A/++
Ly5tcGC2mLGSAixWBPTVYLIIawDLeFzG6L3MQ3Mn+myThr9pb+urjxiPnSOvxOwcPMdLTTqe6yQg
Fg/QTs1Kj6UxvZsR4Hvf+n9vKs9UNwEwjqzEdPQqNwK52UP8bJKdbIEODuEWHDgCnVK5ErFeOHOU
lOsJY6BS1LpV9/LEtdTK04PjusSDG13xoyueSR/OVlqeZtwGJdBGuD/TNHj/n3RSKnhYzDGnIsRW
9sjAG2n49dnvz5myr6JGKk+I+U/AF9OaJCjj/WuAiblmpfPoZbcYLMHfjZzA5k/4ZHhTZfVYBLCS
eE2NU3x04bjrC605tjka3gN76qowTbSUwVj1oJpetywb3iuts+yzHu4Lh9e+bwfUAoBwrPThUs/V
oEtx2dfLGLQQhkC6YH6dCThosNSTMEcPEDgWCGw+zjfDMqt0OsaWc6PJoRTv9KvHbT2NsyHTrKpC
yIY2L+7qBxK2wnoISOF575RudmLWez1EzfD8amdAnSz0UwlY94ezBohLKfPwinSaw+B6pUjH8OcE
H/YsLwC7tWAm/4Xo7IanI3P0AT1CWAo9A93ou9RLFybEyCEe5UCJI743qmGo+6fKA0v47uLk5l3l
QU/NSbn36Dv+NAxNvs+11pfw9KyNKHwI6Nf+y6/BHN1hTbR1XDek1gr8Cka+Cz+kCc9avtiKm2mq
/huvnpm98JGJdSUKpKxp34EuGJrG8Y2fVYRU8rigP2nLK9q/Po/eNtSE2vh3UJKx9leR5GrMg4Rq
dEwX7r9Qd6gsGdMFrmzaYjvLi+JVQjnweWEGQqTg3EPva6OzILIJd3zmfbKaeteR8Qa1xe4ksCsz
WRPPAkTak2B/lNmPqAZkaoAn4Z6YOoQlnb9ffqCSuT1FZuu2Ic/QA6zCUyQWsBwhJYda9vOMI9EG
r3nIKUXqlCZ2h7PeSR0iEFhaLZxGcEOW4EtcAjG43ludRQPWRGEsmtQQeEMpKJAB3PaJXPrbrAzs
OANQ0X+q+P1Whg/CjSAYwoCBiN9j0N12VlbjXiCreMneC1u7lmI2gAA6ioCtOp4IM7UIK5UM80l0
49/EckzFmapjpQm1Q//8hRzrfnWk+RCP0d6eIadpbJOrs0SywvGm1mRosJj66PHmq0LSIGbthKdS
vHEjIX8rJzjJwMw3qwHNeXJ9IGgbwbXqpwlE7sRj7CuVOuyIzqEiYCwj1cP8nwf7pr5ntk416KRx
Pte8+XMfCVsHUZwNpU/YHtZesMCGpTIx0HlRpYb8dICJU2yJ3g52X+dszSIKDzGvxxT/wO6VYZ8U
RoKoXHDZGMDKK6eOdn4W6KcJGmQVreyccJVwIBtKNx3VlfUyi7FOadChFvXc2kQXkCD8z7GP/X6W
1v9AA+CGF7jdOeeBFupL6ASUl8ONz9cw2irmjlgG4aUoIgGr2LU7wXRkYT8Q5ojSLG1AU4fB7wGQ
/9iGhxKvh4e7Lu1CvhXbfL4rklik0YJyU2jX08uJoTFuWcmKiC9jcsCjGLKKZhcm36pBqCDvFkN6
UGW5G7RQxYLcIbXpoXilnUu7eZ8ysi6doZfTmVoxKeuZ+uQCOfsJzs68b1PgMYCKtYpnyZGH9xKx
ncNZ8HH5+4g9mU3whI9O54CiQSAKesqHrlN4qcViq6POnTvbAI6w1OmFKhtGToyuQoUsfVJoOr0u
ibepVBFTFtO187SH+PbluvrXW1rzL6yfoxISDZHFGUiXd+40H6Jime7umkCb+SxNJ8jAAJIki6h2
qoSHLIvP6THjxTz8uF7w8Dlv3YSdbdhppTqfGQTQxkzEGjaebGyLjP4bFiDTSvqdHTRan8Iw1BWn
+b/HjDsTgHAl8RdZpC9BXbr9qzS1pDegRLWwgrLLRrSErcl9sqioVrpscLflcq4OsI3/2EabRBPz
ebxKF1uarJCkkv6Imq64FvAgthlkXAyVucEI4Q12iwms5liy4oa5gZG2vKUToCjqdnytYajbmTNP
aAhj8wJUC6aYfU0wIGDw6cB6dLoROr86dsjBPw+PbvkFBa07OciS1xa/b8FAbTCqN86VUBQQLzNM
fHrKChWBalOkteHeB8IgO68jh968SVa2IFa6q9ZO6PSzZ7t4WG+ezVyWYR/pTjmwPMC8SWWghQ0M
amoVvV2f5ZsiJg9PtDEoaiMZWDRqWTvpvRrHI3f8oHzxh+QYgGCEikp+6MkjziLEmaYDEWtSPBMc
CXPcRwjuDDSAPARLnEyoAX1fgwVOePIVnd+U+Q9wkkPj5gR/cCALNCNZTiWmN8+VtS7uE5DCs+QH
jAwFGu0SjyfG+81tWzxY7iGkBXk3IyvikmoTGSjvgHfeNtij285qFUzPAwVDZROFLqQI14K9xHOq
F+pTn4UU95QAPtCjMegrKB1KghWambjDzr2HHP24LbhlOtPPyUnMmbDTVbAghkuSrWKr3BGKiuLx
HhBnvN2CV0HtV34zEqrhZxcKHVzfVM3ER2oMzDnhUcBGcmlGe8ERFc5ZANSseOpuz3shQvm0vN+4
OYDPa+05wzgJm9g/nyka9cD1NMeMi1a8xJH3pUOW68HTdxU45QtlI6/9muyDNHevVXd9bxGioV47
w2jclQTJPXu+P/3wCLoWYil9CXWVtdOhwAgS1FcSs2wsQgF0cZn5qTdBmT0iC89+BS2sw843+V4l
KcZZNxK5m3f1CXR/AJziTwkPZjp9LPALtR/B/1Wt1MZILH1rpuEDl8T5l+vLKNzPYgkkB79Lq6u7
6OMjg1e//EIzw1chJTYDN/a31cb5mDfEKzXkno7Z4Y4xjasJjb+sGK92y+JdmB6+TYfTz0HVX0wh
gVKx0vr374dSbD5tF36XHcAUkk84ubL7x7c3BijVj8rjQ3adVU60YMMDYodUJmvUbBtFDb//zOdz
91Md5EfuqJyVjpbh1lnptaiFvl3+PIpmj7fiBiUU86+HXNXxwjDjzbwMRTdubIcNwoaJVr+y61NP
YRZ3jNt5X4wCKxcCcLtltAaYKTD+4xyntRwolnQkXwBYanjEjdSuJo/14Haq+rI/JkgLdpRLPbs7
AqrGIUjEw5wsWkOt2zWi+tFkhnvm/zy98A59oTrDz01GBwDoE81eTAr0+hbFY1HEEKAYFIi3IUtE
v+gNDLIZ8Nf5ZnIkV44xMk7/WVJdhbHhGSc6le13thoDfVM0+5R7iUq4eQt9TvITV7t21yJVT2bo
WMbiOdzNgTDjMxFCffnp2jXAIUHGv6UHheRrZzrhneIhaPkij2N8sx2YeGHMcHQW/YmnXenf7Wrs
YCHK1Pj3xpcydAN1LIjOu82RAIIxXXNSh8f20FiT/3kUwQeUaHqu205zsF/ywZK9/Wj1VfzeEu3l
HOiGAUzDtw+f/XAmwtgR66kAhc1/KEmJC2U5wa1pOnmpfNhQgPUuE2/HIyK97/Iix2h+8e3jeNJW
/JdmVmWAYZ8rpu5dqGy86A6LZKaAZ6J9YUiTniUgIwpxn9h/9lrkPaYqJogGjVAhpJ5sGUbXQG1e
OgGwwRbd1K+ZOOCM0m2gUIZ8I0oN8RIsmac7oSwJ8Cj7CTIIzgrSnYsEmVqgyiQxbMuRMM92IRPs
7UKSqezGtTY6yeJbP2jtKqbSGr67eSoje3VtzL9uOXhQn8TM+TTdYtD5SiXjVEuZwDmlDf5sM2JH
T1VbrTmEGNegWR8GIDdClzuxaZfCIwVNwm4/NHjJM2z2zya7nip7QaIymcRKLrPnSbHE+YTFmR3U
iqUR/BmCuSEWFHl9SYA8ySYA0cBNkT4/FfY7Vv4PoFIyeotga2LUZYxVEPj6ijC41bsm/UQuGRps
YJs9ck0JPfz5IAGWnpLlOFLS/wxE/TumZEi5rDS2hVxWzj5fb2rfmR/luxjR4DDwdlBh0MZ5gNqr
g6xbIKtW2yQFuwnhd2RIw4mMPOGLJo0kB76syAkB/3UY88bg8geUowETqo8aGkues6MCF6d9eszp
Zmuu4Q7PVkhz6qrvOKNNK8FcX+gt9XWares19XjQqnVp1zKLsjeDdeOq0TR2WrNiRVPSaLp9cH+D
9DB6w+TSdWlaQthRyJuI/lwdcgHxH25Hxg/wdJ4NFzcI3iDrHC/eVV3zVdfjImSWrnx/yBVEOUb2
f9ng7/i40Ot1CMeBoNtpJFW+fODMWHaNW6ldlwlGUXwI18Onv6FOCcg7oOWUEV5+AWnR6kt5P7/K
GSPibMwrD982C1puXJWrMQmcsi5gDtkDz47cM6LrVVRiWNwEzTMF8f0dSmpMxSxIUoDiGNDt48g8
L8Md6uXJJJVcMFpdXopwlmVGJffh2h+K1F7OoE81nTpW3TK1MUWLo3BCVUaj46fwZ+lJkmbE4LBU
ro1x4MO9F7lUOHM8HOZC2wjGfTBc+U5JrET8vuauPLuK4CktM68b35dUn/aPNo6rUtSWDi2thxz2
/w+oDXZAvR6MtKLUgjFx3r43bHzU7KzBudDAsxIMYIaaCFEcD5ccx3Y+oj4qYQvI6PWeQdP8ZuTD
e4LObsWM8q1vB6HU/pWNLsMxUOT1mCAPpjDEZJbdwlTbIheFEILKLs5FJmb10ZH66vVmXHE76tcz
jjBdMZSRW70Jfo8FfCRPkYYkE7I4ERVCa/UX4rcyEoYP40/qtoYRGPqpaOfSt7OGby3GnVpnbZpG
svazg5wzJ7ho7aa7rJXfspaU0jB+Ym0TJQaCGPNobf46T5kg0xf10AWomXaiHS79cQv5AUZsZGYr
4W+Bj5tDf0TLnnf6tshXPLs3Rv3oZ/5PoJxPzSOxewIRtAAqZLzDCNZAeN/rIG8aMM3rX2AQJ1qZ
Bjnbl5BRfqkXcs4jCq/q6OkCP0h85WkdrSlDw5hN6wiBmGlEDiyHb/qCZ8WxoMyral1M88C3WmBF
uuKOpqmAl1yOkN8epMTzb7nU31XfJF1Lq4IPDSbVV9+LvPpDDaoqiAaiYgdH1uAjLfiCIN+0W5i9
QdLl4hds1k/ynQudGf3pDpckrWRNjXn2Wf36bxyOcnitQjjZoP0/zEO3iTlsayCJhOLoe9opGpxT
44othYrTVRsAtg3D2QFiPawVQvT+O12MXuzEZZ2T4n8kKOgLTkGwY1ztJA6g/JdQVeHu4xuSsVXL
QVaKUAq7+LtcrnRvgy/UMsaWPnbRKOSAoBeuX+x1FbHL+5tQrgF6xwv6Ss5fhHECl3EbBp/qMMXJ
I/k5Uz1erwQVLSPKb8BtRyKD12JV5n1o+dqlxSDjEwezT+IbFCnZxHhVtr80Ieq+E9Ms1EJVc7tB
ivcAPxSXXxNsJon7bC5rPhcJ1wCowJbqQo6rYiG+IaiF60c8DyZUnY6/m/QsouaSzkb7G8kPUOqc
fSzxJ3oQ0Suv6TJqMfJFgWVqxigj3kLSQ8IEnyV20Xl2Y6kY5PKz2/iFgamJo9J70ZvWWP+Ul1Gk
pFKYYWVbN3/LkxzrJ0zkWCi1XFqZyKkDjfG4/BKFHsZZnOXQjNca5GOg7CtS1GeG3ruvc1GpQfTr
4KT/Y0EmCiNAvcvTIYlN8ghfAHnjsJIW7DH4CfQDatbm8z4KkhV6maTOd5KlgRzJkTUEUcauIguC
K5qH+NXABPcVYEOfkEJLCnRbXKq6rTGYCxTq4C9a/z5/CUx04IWyi7Xpfn22wEVyfX0ymxoPj0W0
LPw4gVxsLCcHB/ijnWVivFNHkX+LKSIvxMg96YC6kw8/raaxPHRTWjw1xt0stqlOEKFkfNuQdXH8
X5cJAx67OqD+3O1Lfnrgcp89W0KSopZ6F3TV4cB9lF8cLA8Fagz5bDmTaqt+WwlrG48aCR6x6JS2
/EPes84ytxu9c85F7g9bt64nPwG24dj1MekM/aoiuhsHtOPN8A0RhwEzPu1qnKOnP5Lf7QBCOsn1
08245CppKOgm6THjxl++napE3iiDPYLCdg0DwMceWf45jOjPfmgmNojvrXf1ir4hd84nIadcHka9
ScxWuoBMEAINOAjBxMFpLFlnyYRxRju9o1ugoG8kuT0//TrNiL0fUjyJjIt26Kk6ooFu1XyTlE6T
DH2CFiEOIg5Dz2YlLHS0Rcryj/hzJHecO4vuUg8KeEMVndOIrimqUPmyk71AEiTCsL1SJlO5sFHm
NwofrbbyFYaLc9dsWZawOOfo71aJQYvQrbWlVm+DB0ghajop9sGEfSJrab+g+2crbu73pBUbm6wW
sHuOg0k2CITwoVj8tiN1KDQiXm8xdWH9JTSzslPRF1uxGcsOFNDzEwQw1A7MVm90MPqzOHyWh1LU
MCmlZ7xqFRN9Q5liS9jergD6DWFhnYdqmT11YatJNd/D8k2T3oHa0InpralL1giB0287YYfHfYrI
acR/OJ9DWExdOfc3EU2lubhtHhYDNmGp0qeHTz/4rGwi5/vJANYAfTQx4onmHCPe1OxNSVkngfYx
72vsz2PHqM+DFg6So9sYkmtWJtTT7A3hHVLLsy+OW3Wxt6g5qYxQvvRDXcilXXOQz6zG94Fru+az
e6BP9gYDTzwHdy1h7TN1tTfP2Imlf9L6d3mNKO5K6Jz6UlGz6rsWc2QSp/oU6u68syKf0M88h8u5
o17Yojrrtipacm8hzNa+fO9KiiDnedkWdY5k33B4EB01bmgr6sVc66+8DI7mDBRrwUFraQnSoS+P
Yzht19MXJB/k7O85OCYu7Va77ok0ISiIBPp/wNHQxtcU18bDUoc1OEi6dzyjc9V5GPUPzIMKitAC
n/ewcp93VbCSETntFEE9klfdnVU5fmk01eThZ5gKtclRYS3NtcXtoSOYvSq5qZVNYb+goIdZMWsB
id+xZI8U35fza2HDvT/WrzLnV6bQynjSRPwq0mAAdsd68zCql7VciKEailXE/7mfcRpXd+MwVK5X
kR50SLh0l++SeRaPEeZlVdnWs3wHfTUd+DGBD/aqgSC7jMr4HujBFnUR/sc4SbHhROWzMDwyoN3o
8W9tPBnhHuSy/T4IjksMwfTA5+2wHlFHK7XWzibohng0BJDvJV2MwDgCP1XwuW41Okoem/N6mUK3
whDeKi3yy02MS4uAvYEBv0PZCPTam3GRoNtxgLglYZRJ3v7cvXx/ABr3+yHSvZFMY/dkeojMukSC
C53kJSJOSLQqrOWkboPywFe+YMxwriV+wi0pFZdgAQe6PpiYgTZlr/e7Rf98xOFxL9TCXtRc1J9x
Hv1eF8UbeNwHHlBMIuxKhQjaXosXZyGdtcpGCBI6EOUVB0sfQF1AO2/A/gxugd+jM0MFqlBvocOv
gMGxCYKszn2w7sapA0uua+AbVTP8RMavrEcpsnFSM3AAFQWad95m/cCSFHnoiLcIdoue3jO1ATTT
+pD87xEL2JGhg2Sq/95p71aCg7NWNA+G4lkZtp8OdR2F1ocMuuxRxBygeO6nImceO2Za7645MkXY
y3Jxmq3fUxmb3GlbWRZogltveytU/50nBxk5dzWxqQuPMZQVXLcm7TQ6od6IwG5U25UtwNDPjb/h
onrTXy40ApEFI4hxKprAzAAWACjoqWK532XDVJkPdC7D00d2mG8wuCIDq7H3oGy723QlQdVj1dNw
0CDmKz7r+TJD0/NslX2fuIc0hgPaHsPeaHDVP6FHYfBQx9Ul41iETKL6iVy0ozE5Ce9JBFA9XFps
rOu1Y+dwE90myxTUuZFGepkdDZoGcurw98AKvVPsdvL5IgqGNSN4lRWcmz4O19Wvu+4p83a00Fwl
9S6Ka7tFeB8k1BwKxJGBM+lMdlCERrNma1CfTZx8bgJ6ByHNKTDW6fybL5y0JnJU48CyB30KJPk7
ZcoVb69ryp85KPDcy5PvApdMS5fieIx9vbNJSSasV+eNzxC3j3MzGqbpstVXj8R1K1H4JLP8jvax
Jdakno8MGOhB5pvr67ZfL8R6muVodUP0hzda4ACMwnrzmOGqFZ6V6BNratOO6b3IxLXuarpQDLqG
cA7so8KY1xjEaxZFrqt4FGwLenBXb5Ycde7y36a+lBnd63z9Rt10MKLviUL65RUgGYQyqXo1Zdfv
UDg1D2YouIwF3o41sWgKopSXJSO2yF7HSngBCIxUYzYudPCJilKCO9S6UvAY3PqVDV2iK6i+xDCf
l7BR2pJE6MUEzkfYJVgBE6wj5wKfHiZdSUDfdZrEeOiD0CcP6LPj/oqK03gVLwpVfOEqEDQY87pE
K6fwJhZo1pdCz4oLxRhCsePPIQBYr1emhcBJBRhUkluvcDOX732GBzwqRNnmzbUes5eiFr72A/Yg
93mScEEeCZlrIQN6BfIT23F78nL/WalkK6GkCvUiqUNqSbbPIVAMYTMpMb4ZgK4DlnZAUZgZ+86J
FMjlL3DieLWlK0Gd1DrY0Rrdq9N5iWuhpKwRDH2RGcbRQtYviXpAX5f1zYnqtpzaqxzXUWE3avDl
ti7axenGs80Tjvfi/cYusY7Vsb5OSOycqdtL2muRDF8oHbfJR3ZMEN2Fbf44G0YGf4G0sytCpqgB
TqgiXR6gAUfzHd5iSEafxFQrAS5l37gnCAX/cjcV9lDVmDjnCgt3ZrjW5eiUZ+lOTVUXTjl6JL13
kTPkWnF4B4MLSJECqV8X0UuNn9SrOI4Cs6T5y5Tgj429R6PmibsVoa0FOqDRmuShAkDog8n9DjvS
9fk3C0wJODrpgiy/2/qWoJ0l2Ouz19yaq91sZdGeW7youX6S2g5RRQPl1LGFxaDnhGSU93xhKFj5
qDyG1Mg/k3f8MQah58YCEq3A2FzXE5bPiTMRS7whhCpR5lifdCdTEzCVE7YMvAYEcGcQ4+sNNnui
JQa4hknOKHgh4lG4m6yi3jvdP63+Ah8VLNRves1Fnbf4aW09XcQY4aFTTfy80UxWAiNhTbbgGjBZ
HRfnmEG5vsxq0dVrpf9eFSdA7kL9qo6yNaHgBhECDoHKTsxbp4y00FsYKpp6bqnSRLmqLexqBHTE
lr+aSI82mNmsbDQZ9e7RIakgYCnYKd79Nq2phvKGLv9XynsXwS4b/baml4hRjmjXqxZj4wpzGKyC
e5Hg6LKYHZnk8ps7TrCvDtNm0ijt7IvjZcQFUGc02XHtceSAsM9ePNgbZtu4YTg1YJUv97JeEa2t
bXhhRWY4XsAoL3k00fN95WMKDtfZh/zSSURD3lC0zuYCXnvr7k5JHx28J0urCKuAc7i7bglL9sUU
fEjcBciJNKBxYe9Yn7jk5Hg0eCZRCu8O4J+F3qyEC9MFqwKfFp6IIbewpajfkfs4HmbDo8Ofl6mS
cuLym1MV2qLkcZ/0L2S+0nwEzeE/VvH4RUw+PEhfCmax96cf3lgwmYUwQFO32anUtUkacyWhEREG
IREhJdMpG0Go2xygrIohsGLgLnqrtmCOK8FlmpXgyIz9ynFBeTu0T7ws24uSWN3psP1LVJqqv1qU
iHGSxhvSh0Qi8gVzVwuVnbal2tDJPbvGHGcqjsM6uhyEYj+XzxUswPQ8hvu/sisRWDY5yVqtVRmr
a/eV7lO2O4Z5ZnkmLouJgsEqaNa56BRzP/2lKJwDCw0TFZB7+h1FpkzIsYfBvHI1tWRZXMAemH4T
lkExWOsN1wzHSVkRbQlSNkbjzNKt9BM1dq1j9oTpUN0/4p03LUd/++ttOEtUmXwpLpObQUMGCdvS
tCxMPBlv3Km7yhDhzOn7jzqbA1qmmSJDuCWBODbVS0x2KmwmEFBSIH4blNt2QRkGTO5QhWzsieZ/
brPQwFaCAHqaJInH+g5v7CLsz4UNXhgf+lfUwuquTBBxnt3HQ27hxW7eJod9Mm7IAkBQyEF3HzeX
iSFssMqvzNkVRcqgSuqfjxG5Pz/UF79ehE+oBQ+gRZiMtUZdkyOyo3LL+jxlMYoKQW3+7PvdsiKA
u/Ve+wCiFGMW+rqKlnw52BKRRSYdjFqI0N/an7UDxko0H6xzqlllgn9ATCjYb97D2ylB0EY2CrLt
Fh6EKX8Ja8CbbYWLHh0A8lgUQGBBYvaTmmfgfhefwxE6R86RDw3XOZ7scoXZ0k+M64e6zwwculzS
9ZmO8ln14nT8it/8F81/c54vaVT4jSDVtTa+lapNzoyfSOqdQoMWL1ny/w0JcOrB8/89Qy78gXEJ
hNahOXTszeb6VZUOlaML9r7x4Zl6mqfd5BcccnWMSmUu1fTpmYgonmcsWLRuJ3fv2tRhHIRY+82M
da6lLiQmNCu6yFV6CB1LHJqhgfFLWXYl3RAUFKU/02I1P4hyVipr40Rnpm2M9jm83V6ap1D4KYFc
9PRT91K0KlOPOWnXRaS0B0EanbeYr9s4xKqxXNsJziyKdgnEiL63kUD+fw8AZeIR3Z/oF88hyB+g
toko4hyoFxvm2isus12i1L1un8G6PZOnj2bCTy2OxNMHRzpBFXM9GXqOV/7KsQVOqX6IXnJXDJvC
DkoaWnJGzq18SSCR5Sv7aww9vqhFmoyxlk0I4sNvl1gLiDqNBQpd51XJkmCDw2Og+M1VyvVwzJye
YsbHNu8XP0WWk3BQxGVEpJZBvrl4rBIPhwU91ucDtHuNCyobDCYihMtIc9kLScATsW85nqWaFwEg
aVwFb9Svg38o8h86BqMvyhIplmF/dIxxq8gV3ATZa458njtcrzYeIHM5ikZuHGtQf2OpvFJ3igVM
sfwSi6TohfZj5vyOWd0IC4x5dDUf6c1DZP3ysxw+dAm9qIvBsjF6KlB6L21708AjpycA69iSlpmI
iX3ZqfZ2Z90TenZLPDM0+ozEjuauJu2dmgqgF6SmxNVi32qZtR2PTwy5baFynIxClnXstxKrlhrz
muMLoY+t86cywv+2hbZld6VWiu7eMHRQF6wx0eQN07smtAMDhctasbArQJNbF+BbJWxD2dOd2Q8W
p5v+PBLuvDTufayZd9ywm3z94FPCiwhw8qAb3vLCieXxclIu9BBU8Ttbdck69OCECLvA8cA8nmyS
iSvXpKRCl/fMMyYxDv2iQWF56NBvpBHiGK+prueT4IFSlZlaS/WExPZjDJCUTi5Dv8g3G2ZKIOb0
NbXO+is+VmYTqSXEkaxnSzFzYjuRE9ZaWPuX7cfPoD81s/Gs9F77nA1hwvY/pQ/WzEHT65Rw2m1p
1wt2+v9onSGFro0V36HirF4ZIBBARsAsu35XqdsGC7dW9fGk8onszs6Ns9bvJrTXfKt8Ag9y7ID6
BZeIcP2lQq3kkNDCiimAoIpVZDauP/f/HD9m2U4kFySiHajGiM1JzmozjvEoLVa71ykX/vxvjMgg
rjyb0Yg2wgNf2ZF+2R96OyQwHoNH+eezcFaUpqR77rJsBlmSSRLi6PE3LZ3hlMkSCcv4NXvFGxdo
depLiD2eKtIGh9o7K75fNlrBQFm73q5CzfVGJVLAJ43UdMBq5FYuskhoI4zmk2gTkcdYTTRvNRIi
DCzHXC+AreBPwGr2agKS60QisDtpoC3R/KKlhrpF6HWpZzY+7jjaBhXoKKh57mR1OtVymK0TFnoY
Dz68WULma1WYVjXJxr0x3qWNqTNtqOVqbb5UabSk2avWP1JUNqOdn2xU88hneYohH4/uApvZM2I2
ZBfYeHv2msYz4gJHSK6uXeUERXInMZG6WoX+nOASnwvseTYxvvjSaUwYSJAwN+pCqd5jDKSchbHy
+ILk0uPnYK6l80xtpPeF+2HlpmQBd6aGrSVwm3m6Hc0QEoKb6Gy6pr7yH/bOALIXpLoux+Y1tidH
AVsrqOpQ6F9Kjnr3TQAOI0mOikhSiL55Tyta3JK8QRGjZ8r4KdXe7H3BB6h/pvFh9tPyXXqKw2SC
YQ1tdL3EEzMIqA9st6MKWui3VDS+6QjfPy/KhDWQXc5tUjosSscSau9Za40CEuxC4Nxs1whLpden
D4Qkqc+2zMrp11UWzKe9dI2VN0KTFCcF1fBU4ktJpVV9pxY0kB35b99t8j0vnqJHGKiwih4BEJRs
Uqyl2OeVOswEkqDAQPo2I6HqufjygpN2XHWBLOhFuz3Dxn6SpJaKjjoT28XZmOeZpBNtyXyuOnom
wK15igmV5ojeMEmPi+rpWFedKEtHdYF71gCxgKp7vxWy01OA46jqjQrG3Tj2GAwiWzEfdVUVQZs3
k85KdW2z3xoNf7NpfAAzzIH5qVZ0gzFWo1dECRRQcmIQ4pzdHpniosrm+msshsb11Bpc7tmcAWwm
ywBquyPaW7EZ1zpjhELaY50/GtjE80JR6u7QGW3R7loYEIYMMCimyT1L+dUkTHxISzBvugRPqRBU
luOSjl0X9mI9NUIVkDWgO9dHCUrTDsqJnMSie377WqdOhj82/wpyaSwtGW667+As94lb7TpKizFe
CWIhcIDTCiL7Xb8t0DPfzV6eqrLiIvHnaEGwqXOuLg+Me1TkMqNsuPVXLHxZkcbGPLuMhn6llBFW
SO0LYrEEM1hPfv8eSifAaoJ0SnLs6tQjbnrzVrnBXJccOwVo/YJS3LPMcxqfrrP3yTHxtM0Gxjsj
ouLJuOgQb9pKUDJiGzpo/Zd/pPtKn9J9DNX3nD826UIohFZzJiW+5fEI0Pp0UJ1GojESjvCxDBSy
g6QaH/1yRWiJ3Psa23oaVFQYY73IoIemd6rYCOipxHsuGANo+jEGot2VJuc55itIxoLAUJOLx3ub
CZQBF23R5JnYR5gJBK/pfq75a9bIrs4r4ZL3K9aNxgJEBH4Fu969aHssNWNVZAi+ypRdgTzzFdxe
ryV+ZwY9/iCp1/8bDhGECWiTG9IVhyLMRLTIcO9zZ1cxacXq5rJKLDTclla7CmETnuOeDes/1XWx
Nh+dVSpAtcrbLzrRauaENEIikN6+oGjSTS0nvCWzlm9UMMR4LNvdBN+ocC3SB/Ja351wylaGZ8DU
USZQPG63t7r6TgSRhA3LhpN9uDBfjKZZc98HmrnLecgI6HT8EXVmARhdwdNsmPXzYnq4P4E8IWo9
0jAeqv6jiqjN2UVk5dkYgYYHbfwT17EajbuydNKy3xmXfCfDCOzKQggqW/13a7+AGfr2vISVSISL
T+C9TtBahXzgOqObd30C4spFUapfi7A3aqNMeoGsvbd7rr6SL/SuI6jaHtgITKqoHKvTwGpTfbdO
ph0iWcWGj+6TyDgumkt5WBtS3qusrmSQuNIu0NaB1IEu0BZRRyqQ8VK4HRcumhg4VpqnP/VlSwQh
2oMavg0gYV2u4IIVc4WkR19zT3YziMHXmcAEmJv5OG7XBw+M2IUm/PONEPixG71fY47U0Qo/Zx09
taz2whLeB+NgkIsc+lpYzeWcZtF3SQZnm/UiXxc95l5nJkf2QLIrRWMF50aIcIlp7OE/0LXAPRQE
QKmyiUGy2ymHAj/jAEYDTX2PpBxPV2P5vrbcMmT5rpI54SM/h+lPbwSUEH3Y9CTtlmkvmBarBSn6
r5WFT2tgh3OisJuCeBsC4GQOBC1FuVAfGMBMY4UV6Y3QqRT/9r/qFyAyG6UUPoUzsFH7t/UOlk8O
J7ywZVkUC2LWioGHfAqfL5CTut4IEYcuXekn5o61c4dStr3yqU+Dn4itLbcc3LiLX0O3cLCczCDg
3qNEBXCOl7YcNoJe91TtfbbcbaeOk3oAi+Fnw2CfxVIY8kUFYaa6TTVbyk0EvugOztjGn4g84+qJ
RVyLFzLAb77BwGvsMUUCwB5JWERuHMzM0ZFM/3+5wyNylHyCj6vnktGGz/+y3xKAiX2uHF8B6cdr
xEZgqbdrsT+08A3F8H6nQHuqeNkDcQ0UIYGbg25ssXyU7urUOasGE7WSokqQHkLPFuvw/G9qfc2j
fFr50SaEbP5FJkm39Z7O0zz0GAp58RO7B0lsYQ2Q2ScGFrArXihoAPteD8gIpd0D9GOfcJInBSP/
jj1wnfgIDF1uPVbFOrAjD9v/EB99Kxvl4UtO8PyR6TmDOhXDn6mIvEsos6sUBtuiMZsRT1/9yI8o
vyNnMvnPUOI8Fnq95XcSZDBL8Isa+2UEejf9vNHi2QXr4tELVLR3d2kMYBtiEMv6ElR773Jrxpb5
ZHTS9y+DMHajfMNsF6gZXbPhcnyIV0YnC/k7AIm0YzIFpBTzKXCPL6Px0a9ObGm10SJwOaJNfNLa
2zKTrVYVnfHnvYEgQwTkHCw5Czel7dK3YssMedY67kNaks16D9Onl0n50Aj56213eRKxlvV83+HA
35nUeiLfPs8IihvjR+f9oevHdPwboiWZHNhw+fo4e+ep4NIUWvoyOUmmPnzYiWNcNpweweTLjssB
Nd/prTcXb/kKX9V+MVREY2KtpgLx4XDzTpWBKb6PZHccs7Pc51RvQThMeXt/iJ0bl2FDtE2XeD5U
SHI+grqXW9FNN7oQj1BZ1qdmtkTGwZKDFvn2u/Peo/uut1dPnve9KqCOmUAy2paors7zMZA0hloH
Lzp9KRjN98RzKLusBahAdomptA0S8svhqTHuzapDye9PHPv5Dlhh7o4u0lllIHazmBKAFBKJQ/vG
KkqGe3ydSD3yfVHRkQvj+JCs3LwgF6pzmcZG6AWn8OPhOewblH8jkb+qcn4U7pa7+7yvlaVILxgy
xm14SvbmUijO1uiIdyt6Tyn/YMWxmtIsT0q/S+E0XtV6n45l+yrRJ6UV3ji81RjXb6ipOxWcopwi
X80JBZJ4B9zUL8T/BEQK43T33BQLwt0B6Q+3vgpsOKpOaEuSYuSl8XCqVsoSrvsT1rz466+4Ka9J
MuFUIuHCc9kyX2JifmgOpKGEJYYrU+qGdbDJ+T2yfpZ/L2b2YIrxRu5KUJ7eAJhRESzx1blZVtxK
yXDfZnYfQgn/YSD9m3RSlIlMYpvYErCv9T5B57833P2WYrTCHCDo5TE0bE8D6K/gfLeWqTfJpif1
kOoFo374qSvwm5DmHnaLZIQCF7Uun0haQVuTmWzhE7xCmt5ZKTJ/p4M21Vdn7HiBnJTvhQFvhx++
PZzr4Rb0tR33GHmoa0l/soGXRu0mPjB5Z10zSzWBnpa88Wvve36tPx0EX8PTXQFVi8tIVc06lA69
6aFUBgPP8NtJMn81ITaBMhQMUOjSbVODMDavhLjVvLAQAHduU+YXVjIFDTXdNUuEMWj++iAUm6WH
mQow8/k1SDntR0m3JBAwdJw3WcQ8h5l8oMBOXGvXMPPgtciGLalmf87za9bf6CZFePKxKz3SgGlv
2bPJJdev/7jNgnIk3+oJUZsfpUMRUzFeP4IDjqFXOZ4/h4MMeO62L02XbkAjCXLY12ZAdYVdiKWX
oI2/sxyy2JN4HZBvkcnbw3IA1c+UzOQVoWTZ/GPCBPd3pNXjJTusVnbDrQu7iQrwqqNtsrrOwcnW
R/eDnE+faJUGFGreETvkAGCD5C8l/FDNwFPssvYnc2AQ7ZyUb/Yfk/ogYyDq2znnJ+lwtVFHvUQt
5mbfPkCBua4GAdAIZjQXS4E2Xuwa8aDXPHhUiA7okQGqjvF/U9mIIqia/l/62bfoVaRD2R68+L4A
PHj50aUT6ulfDyAdknzAPoa465smjAB5688IWNAsKPpYQ5yogmVKpKRiGpBE+03pENr//hTUhu3T
5fe2NKWqIZ8aDr+a9lLLL8cmAsfNL11UB8UNIGa2B1NQP/wdwuCYPycjmJ6y5xdn+kPxx75TxkGs
mavL3r3WHHhRK2ENi2hWLQ1vgpmPdwb5QYVFPCaEP8sv+rQ3fx+oOU92aTUeYQnJ2E4dzNiFNsKE
gFdfgFXQWOlxipUfWbEGTSdWlFB0/1oQCabF+2L998kM+Awvht+5Qxt0eYEFd84dFK70GgRt28dL
lbf0UqXUYucgS11ha35UCsjI1Lp7kKOT4tx9zkgnRhQ/lh2biMpqud+PRVCFu1BjgLTJ6PCXUXsO
/9Qa9x+7bAJL9ZoHTqoOmOGi2P0QxDTSK6nOSLEunNnar/n2YTXZi4gYGcQUQfyTKfF7te4LDrtd
qmVIqbvgI22hO6pyUosdyDwE0HKyborFKWSHyeBGJ1fKrZJN3hcYFpXlTLCf5LBENho6j7u7XTJF
6JivxTrxTjVmhObMeyTHSjQaCh16BpgXkHZ0fyRythVPooPtMEtG+NOFtzh3GgwPv/tJg5gN8dJu
y2AoTZ7ILGnyAPpGiXcUI52f/ispmpLJr3R+PUybNHO8/sRXjJfBIxwZZzEyvoJxD7xpx2eAwQIJ
k6wUjp22PYOMJ89aUN3oMT+CWVhloTjM8prE9YJdvWHMtm6iYFduZyQELYepkFRuyZGkAZ0wJwZt
LUsY0Pdke+v/jwf05DPPP8NoQ3JVJeZ0u9qTL7bVcF+xVKCxxrtPszpL0nz7ONE17qegUgg4tNhR
ic9O1Xj2Gp1tCZLqJBrZghB+yMVbhYBzKtR/BzcI0o2AZlfA2ylBiOa8m9dceXbK+pxtIHD9HrI2
USzi0Go4zrICG4ViG2FALfNz8fZwM1THO+JX0goCTfrSrX5j+18Za9cr4inBI4KK1Ns0QMCuigj7
E9t3iju0oaIePib/AKlbuV5hQ5munnn+uzdjxU0p/J2Q5Apw9L8WQuldhE0Pjj9wMoqRIN5yPF5D
GYr/R1475lz4I+il4yEeDG7rv/ciVsTnccaUQ6r0iWGSp2g7eBJZiI/1QgzclxZkKDdpsJpOgJ4Z
3mdEsv/ou4ERjeJWcUuO4Z6PoiKXaVVvYKiamBZQ4Y2LYSkJ+vTr7BXIRbYEGLLxJ9BEniQYzPZN
mTEWxkWaMpx9ZLibew2GmefPvjXbZN2dV0RNGMg16IvrXPq9ZV3zTHuCEhBvkG/ozxb7maCZXPV6
7CUOHf1X5UvlliL0TEpg/SMQFq5aLGFSMxqLld8UKNdqSC3bpxkAHScW7zWTpaSQpumHJ4SjnLny
PgvQgYju/OfM7Il3qt3/jHe6BGVdo6S4Ij19DwQQ7cf1zqzdBDM6T4kly0HPqv3W2b/knUCXi5th
PhhjHrSMx2Fx+kBD4tUbqOUm80wpVUKxE+GHDB0UdlV/dVrMyv7/9sSi/7s5w/tMODt+3PnTkOyY
iRVst0O2AYYhIEx/J5+Jy1TnXrKGmL6bHdZN83z6EXYCnKD6j0c8ylIez+Rs1UQEXF1SH+1ZfN4y
/4G56nsCO8IO7qojGzAs8fjwu2Y94rwkjLbudXNMPxt3ak4AApPZH9Q2c3/SeJX+/bLsZpj/HTjN
zLAOGM+oIQeXp5R0y/QD6LUr3ctL/IVNC03b+s8PuhtPyKAUccY4//evgr/o1DmRTTs/JJvCY83K
W4N9xNX8kyCjrqGKzKAeoRMZvJNIrJhK1LUJcPSolYKqwGHX1EF92bnpDsXBojYO3jFg4gDW650P
DMvldZmnligxRd25SgjeOuzpz0sGdtC+3ZqHDpIUdpFbBw4UYsKtSWVeKvVWl88BfekBVFAcIFaH
ByzzSiwUY+pdZ3ybmI5PyzOH8UjadvSRLlccOpHOECAVEb1N4+uPqcL1rDPQV/euaG4w+EuGgx9f
begmbA5X0y2OSDkNmA6zZkMrn0PuYRl4G6MfIm2OzKHFz1b4NhZSALnRK61MWwaRHW+9ExIj/2Vy
SeMUzfoXrdUllIaILygsBfJKV+J7guzOpBxcM1OaaedZX3VzPWrJAzbFciM0imdyGHO0anLisT+E
5nbZEV5LZtMvALo7+1chnvmQAoxT0a+c2vM0/ThjR//2ZqLjmvh/1DshyEsLX4783YJ11mfRLaFo
ocos5RaOeHqim1rhDFBv3PGT4G/FPNeqWTuF5Qfjry5mtvEZIR5mcIdAYrHpK+sOFcns36sCa5KQ
dueLjiE0Om/PSP8lbRml2R0tdG7sNhdU8BT4A9s2zuM9ipW2fQV7nv57jqQvCwtmIzccUVWqAmkz
rZgyQWTRRgH+VJ/JSZdC1MfAabAs/Fk9EYZZWnVsbJjd/sUpFqOakBhmf0g/dc64gv4OkUDMfN0d
BM0/y1ZBb0pzKSAuEmti3y6DVoDZdQPrCLfSbXHjDCbW1QHnuOrcJNeegiJgdyimRPrpAJoWqPNc
SqhFy0TdVXhaOYAkA99h7LVWufDuYI4VMLjhokBLMY9NkSOOdoth0m8bRA7WSWu3xk6P96wASQ3G
8dXgEXImNummGq5RcOEZRTkGJe+80g52Sc4BZJgA/wfIvOO/Gp/WaFVUgcfNL23ntjGFzLo4eeud
1TDGlcrwZ7927I9JrXtxhkX1V8JUf8VPF6LohYAJVW74ZZwdBSsak0VlMQZYUuZU/0cdh2ey8N9X
AR/bav2CIFtFQ0sxaNAsClaR3Cil7J0vSEcviliJsW90HOz7WiF0qXxFJbqEC2kkhArXqvAm4B2A
2y380CdxRwVXX97NXGMoYxWyr0JLWufQ8Ij5hwPsksr+B8VqQeZmJNKzE/67bTCX2FUDCQAjT/HQ
HDpoFqJviWtUg2S1eF/m1/HZnKRelHRr7UUcgJqWN2/kGwxs8Tg/X9HyCgSs5xUzcdfP9Rhc9Wvk
r+g7I7/r3bQFns91ZTo5KmxMwhGk3ZGRrvvjU7C6CafsU72GZQBtFmt/CEZftWOZL5hvr5jNbHXK
Cgil3Nm6ec0mApQNCzajtsXqZHPp3fIrNe7QGrihLsQiQJdKhVpOjy2uGuyHkrVitNcBVJaUUAS4
MB6YWvEYFn2uKRGufJnAv4vf2KEhUSqSpJPcyhMAU7Cx4QX84a4Xfvp5BqXCK3OHqXpM4CyaPROF
vVjFdwW/hOl8Huus8v/LrUkdjnlak6cvAcGUqMFbDjbQnu+lvJyz9xkExEsanqvPoRKWcHHRqt2j
UlLCXmhOvRbjPPWjCht1MY+7+UffxGBMX0/3T2GRswJU1qFcQEvhYarAys9NM2k6OLJh54NenoYB
qRP7sPYW2swIO+36wnVqfDq4Lpj1BmzukhRPY2QMm01Nue5wzx0zaxZpOTp4MMmYe9N7fFtVw1L+
I1Qrjx72xaZDx26cczzckiW3nD30u8zeYGVDL7nQHeDWuJltMJaYATHO4/Ig2ndcTOp2RkjcJOI9
fnMQdkH8j06cWOLE56cGs2eV/YbY2Cyz36kcjH1RcvwgPa13WRFwh298brcXRC1XKuSHjLFWIT8O
hyjLUebAW4mhw3syrzt+oJSjahTA0gOCfQyST/V8xkEjoxD5tceFP7CTq5BcuiTUn4VQhQK3WjEv
JE+Na1/k6X/HNcLKs0IdDq5CWgqZd0QIVoFTAFLxWsbpVkqA7xSSl32bzuf/bfvgjosJAMYbK6DZ
rTtofrv7hok6bkBTy/tAJ7AHWOMKTobCEvLRMzo7nnnSwsB8w0Cpx+MMLAyBqTeTbGpuLg+DcjuP
fNmouDswVA/30HRaAH3qP0pwyE5MFNW2LY72FXpL9E3gJ8v/4sLJdD4M9ekX+Hp2Nq/hXIvN0iJ3
Mn+RIv0ENCzaKduZvYEe7/wh4MVqZ4qCGz14+HoemxBeN6KEopmIXT1XIVMCHtEgQy+wGfnXnYgP
bBgcGBQwPrBKZeVohpd/TVNKJm0h6ST7XU9W+Y4OlgCN3BnBaoW2aAXgkRNRhfMBNv+tp28tj5wK
lZmGzbsqg7uyrGxjv9wjhxfbFh74q8A/Wj0hfPT4JqEX5ibOMR2Mefvd8EPiDTh4iGBLdbUU7yi0
pU+rCeYgXNfxMLZk0jQgwYkmUs7ycAQafy2wNWe30qNChQZ+e88vg25DUg+w2p5hO/RF54siUlMD
4PU6NSYEN/CwKjRufm/jVoSNXoFz+4w8XOpEktlGPvCMOCOlmFA54ukpPi/ElNQUVqVYaXk3MoVj
0LuS1sx1mM1GBBlh8LesyY1gBS/YeZyRCIbAaV61YaKzMxg2lYHwmnImtqXLY1k2pzRtdQT4SpLt
SxtvD9WYEzNyTb0RBN7c2RyvjPsPkVWEm/T2dOa2IQ7umeSPYI08eqsI/ONK8W0gMIbUF/p5NnXC
LTgglLABW3EdiSiexSo6+M428kimdFSPI5zDFam96VZCKEmxYnSpGoyIfVrpIiImFRlIF3p/Et4f
jS/MIkx27PvyyW14oA+EuetHnI5xgQELTvtsmgxt5RCO6M6oS3qfk3mp4i2emFo3oZvOXfRIxI2u
OpdIinFBbHIT48/GG9P0w/3OnddMxmcAujJ1DhV2g892YUemuLT1E4ayvn6KNGd60t8viZwN0bjI
tElLGBg1z851kAvTMk/pGZUyP+A1YNgMFyiJyHNEHW1xLtrRU8n3ZpOmqk/zNI5sQd8jT6yaaQo0
EkNdTCdrKRaF0Qqb9lXV7IE3ahcdiYT2CSHTxNVxfXQwce7bnOkwFglRX1MRD4i//OXbENoy5GW2
QtQr5Z6etcs2LYNJ2lCiHfQcWz73v8l/aL7rNr01nYBmZETpnJtcknPIcg7BQAg095jPvmnI5l5V
SsWNwhP8j6mbd3vrM8yIBXmFhIoKGHjDJgTiYZ54n8aAaCr+2Qu88Rezy152en5ns7KqBLU3eBiD
y40Lr56VUAhAp5OeV04VXSz1lCRk+KneRdtbhurbea8wPiRS76qzBbxjJzmuv1YHxz16dko2gGUn
9c39Mnj2bLuOugHxOe6AfyQHxE4kP8q9z7Ccr9sOPFiUQ52JJcwlKI4amsjh8bg962P4z3kwAUwx
kZ6VQLQBu+TMPZTJAOPoOqnrrxpHM3XYxCpqqbvz8tQzfqf/5+IOJANplA/GVOZHF9SmNMnYjtDQ
9h4Cto3BQeqq8xE4cMTfd+BzsBdbtZb0mcu8f7iQRpg2WOBP1MAp4G1kQNjX55uvRVnoI5Kw+vJL
cQ8ovLvB5AxoPTPGx+QwWlt+DbkOTFXm3t6h3+bW9WvyEnkE7azbn6cltyYXJpJewwCXU72+fe9b
hU+lce5JtwAeZEb129iSKYmjmRs4ioIIDLk3LKvpc3hNrGCljs1GJYs1HQKmFd8H9/0obgH3LwGB
fkztbzp8RY+wI7ISfKTEr6pL87ZnZ/TKyOWSI3K9ehOrkwfKfCY89f46pEIG9GnMgBBe2+54+dhm
mEUXJYlvqZK67BMUNLI295g2i82QJ7atZU0i0RdMAoHMm5B3n1KSQGtSc4BZdmAVOCx/zcQ/dgle
JshhKZJltJ5tFDmRNleR13snAh6y5oo+dGqlknA0Au0TLEV2LExrQIPqO4WmylzlSdui7nkkcIjI
9UsdSTlgptowWnuuj84YQEyFY289thYCYVlp5HIP14j7s03lPT7tly7b2KQhwsxEIN3R90+LFic/
opTXzf+K0XjkXK5dMnVQqd7g+vYTN8pPhNsponctTp6yq5Y/mQYgeyAofLOz0ZUd7HUW6XG3848Z
z0GhMaquRh2Hg9kYlSc732KDSue8WH85adErdxioDotLGn1Wr/rQSprkiLri4EBsyhzvG4yxj3EH
iALwLDVCEg7dSrdt5eID4iwvkyL7FLOUc/jIu8IiJJnjiaMTx49qC8J63BfrrlK8tWxDfjIg8yT1
z6uPmvJeqz0u+wUht557por74NNEuGsGOVZlgrdy//wKHfQ2ngF0wEWU+Cqcvp/TDCgqxqF2xZIB
4JLuLRdk71DrjoFU0wJfRPKnhwE1v/mH3GZwmHZh1rsOYEmQMSqOV6Js/y+/ePBoMQAk0yoo/fpK
d+8K6DgCyqzZEDzdwn1gNwpRxAbp75Q1dBjTO2KqI5rpJTEf4g6gTLX5hzxlLFZMTw5gpfZagB3D
3ykMGR6fY3iWxuAt6omeqT8gBNpIc+kKlh6JE2krx2T8iCGHFfcPHZOsc97WNyURQYGNnNrc/vwU
AbbKJCUJ/eIcYzdjpWoS0yznfwRs139ywlaegefDL5air7kLbhD1lpJhNyMsu5vvJbWeX4DfphNt
gtIhuqGKnDpQmjaND7vHy7+1FfkdlAW8KuWCCE0L9tq2dgmdRKkyBhxdCVlr6N+JY2ZZODw+r4AQ
axkBKc2RLUFtdc4/ypGK8ipnt03dMf6TCezu56En5LbbwukuMkWPirhdekw9kAl1txDPz8V0Qs3z
N0sPdwfPKB7Nt9Z1bHx30G2hc1Ws7a7+HKrIVDgYFL9t4uz8cxpwzEe2j7xSkgV4qDOd0CWpDb3W
WXPPVB5ZdwVdDBAjPCEpLQd3b0u3xMFkGTE9mfXXbNFCKeXdayMyN//RELaZ+7+9Y1t3hnGmh8sN
yANs4FkhApKYQjtKSQSZw61s+o81mheo8eGxHbctfm5oL+zhXM5KbR/S29aPCf03o+Tt5bmluNaZ
SJbUHbdqwTcSKa5eVAmEsqVeMuVVP32zwWzrd0T8lnD+yoS8UrRMCyyERsnv4Tj9Sb4/eqFft+iV
qyfyRzCuyvAgD0/EaY0TDA/pSIv1ehScyDvmrjSaV5UMC8G4s0A9u6WgMjmhrNm4lM+OqkL0rMws
rNma8blBeLgapmJ71232bekmHuV6Kl50bu7mMge473RnknjWg3ReHUBgGE0EfEs2YGxVPuzk4Iy6
pg9hPhkdiSh9lrfjxoesSrBADKRaKtrL1mres1X2h18CJxyJ0aVirEQRMaNgc8d0cdfbdJq9Tsd5
TxTDLxDHFyoSmH2/YArkX9srV8La20ZKWT1EUhs4dzZ2hNlhMtTPg8diIsKSmM0WnffIUJIuIV+x
rTlPxoB7dAyErW9tVAQigbBJOJrOqPAk5f01MOp9C+s/7HxkKdYhelbfFOCm1uJbsuw14aEIJ1EA
d5IP9x0WK/iEBZY4IRby2mCwQ6c0lf5ikauETurvzbWJOqYtJWgkxFCK2ypvNp7KQqgNvsqlepo0
1YvYXB0oPPSvpRhz2nFh6g9wBLWdX6wGlTVBgBf7waQo3xTCkRAfM2xZs3HuSeNmwuzsHiH+RJpO
VbdIJfMqHbxXh0wpqx+nUoWEokpULoFQGCdsHr+FUBj+475HpQanvHazV+GN1hJRf3rejHaKkCwW
/ZJiaxZh5BEXzEWnF0Kpt/EoWtdMNzY5g201W3wYXJrX2qeDeLYJonH5vAKkMMSmDIzesTuPtBlu
oG0siiAJ+x/A3uWQIJoDvikub+h51jzVhliv5k3TxTmkvIjyP4v+l60A+UkyNVnj8S9zLWJgGgaD
N0gitbaWok6pqdf5hugI+Eir9+wXXA+8bJZ7rw1JoIX8MTIbLqgcUMfIM/hiHMikAdUDtKlanhzI
mGzXSNjoZZVtlNWhfGa8njGSVjxYfX7vGvpCvU74ktLnCi5869HD6nsNGX+qfdL+aJ6eCn1igWdP
iN9ee/1WrEtu+hVuuXO6Q5WmBJ0e6JttqHnmnT784DUMBg2A7agNAtbTlJQfombpZidT60lvLOaF
z2GuYazi3OcQOIQocpwBv4eQ17mKXjtZRKZcX/DjP4RDBx/W5g/1nAE8cJ2+kg7ztZPBNaPWar3T
bkaoq512ZT6bc5H0+RDd8OU/4r+dn/qKaMIepINTY8T5DXrBMex2nqr29Os7G2MkN8q4jZolMGMf
ZuYZQoq4O8sH0PLapBXJn2T39yqiUxvlZyWO05wbSEWeSLOopnuFo1c8+ygQ3E6+0tpVuBD9ijNz
KQY8nVIWsMT7oiPj3G06jlNhMJCmj5RpJGxsEVDA73SIM5q48gNxMxCiSPj59NqM0HSLC7IRT54m
w2sYToT9RD9CfiM4qTk1xQAQcqFlGnbKyAfZONGxGM7uLNX/vSb9VZRfA93wF7Ps8dPGADXGb1CM
G530VqBhSyp7cOOtuHRQOyz6RzEoSnm2IxPY4xZ27UtWYPxm4IcHZ/mCLGCsDIFux6cbyW6sQGAL
4B7aYNn7l7apqqHcw1rckIVcy0RcW2Qgeu9VEfDFiBIr0izE8XthiW321Z+5/ihw+hCPDobGCfAC
G0whObWXPeK49i95mslUy5jUL4hvMOu2MFm26lgONHQC6+D6Q8RjNZjxmKGjAiw3KgGbJI5yHJ0V
DqvjeeQSAo3yTd+eXL98ORbf1gPo4y3wNsDRnNRE/H4TzWOjOtd80Xh+stimzxBuMck0ntEukgLq
azPHETxKCGyIqeZbJs3qzzEF2EwCyJpnJ5R8yvjgh35CixPqKdhwqDUrBudA2zGn2c/fpfZ2BUp5
HmJu1nNruT1p0DfDEFpyoxs9iuQUOSj3wYnkmTvJw2oyDbn06wBMkxDlYTtVaUFChP6+az3kcqZ5
YNfnhdM3AXoKRDKrD1zzsxtoxLKJrr2AsW9zMk/ihTsg51NUcVH2RxH9c2hPzHmIt3YDtos9zINW
gmKARMpFxSe7gS4vF8/1kDYvcJ0d3YsBTPgOCgXE4mF2BoLAsU+PzZTiMp8bPnta/q6xuoHN7Ej5
96QWG6inKQ9lR6H4Gaj24dxmAG+0qXyhELPFldtEf+yIyE+fgqNnUi78BrLyTwJ1p2v9gNguMWD4
FJcH7NvfFvZr9xITAOYD6JhVOLOhcXFkJ/uFwP+qJk6lJ4qPkBFEo1E7kcfsXU4tzbedq/Wsg18U
eJCVCmHToh16h5Yx4qgknmV4woPH5403CGHp3ySQyL25tCItCd9sH4Y7YU+UXLKhOA9bPY4theKu
2j3PAUr7bZ3i+e7Uvrdo2H6csHmxw78Ffc2/irhvF0YX+3u2xpiPnOAInL58ofZYDLNEDdNQB6CO
0CLFS/7mE6x4cMrn6gMI8mY6gptTK2Tohz0xBsF0wsC9QB+AvfmjD3bVNSEY8xEBv6SoYC94MHIH
5FV4iAqMvPVghQBXeo+yewn6uCoh1uZh5CaVSfd7MG7/5E1G/Qm0LxycIRysbOIh5e9kM5rRYRVR
2NuU3P7i+/6dbr5sCW2Lu+HyWtoBLDIRGhEV0rzJ7MfC3CnbdX/FsULRgOFvm/vwTofeJ3Gp3lTe
s6clPXOY6gBNSdxZB5HzAPiuHvbGgHZx98IO7828ZlJfJS9rBW+jqa84BBVuoAxN/jGV242ejkUQ
061FZQ4JY8vYuI9WwbSbkmo8ncwj05jrr31MV7uk0BK37b8DV9UfmeAbYpHto8pKiSadMvAcX6AF
3/Bc4UiwElRMgBd8u4/pvIFAcnlyMaucyQNLufMLz6NCtpRAKN3w9jnSLnAX6cNgjFQACnb4qUgs
8xGzH4c0LY9oCAmwcijvPgmyUYJ8Hab0avEDCPy+aquPZh6uDUPV98BOYUYiPJPj17FoQYObUGd3
45ZvOgeYM6FrXE2FsDnClPjfJdOm6tiSGVc08Pwyr9c21o8QVYpt15RWGbkLsU2jg70TXGepgSFB
G421zL3/MO17e16Or5LhnI7mJ25jVI4ctJdxog5/CSK5nAgoR15mkgQtkV/c5tC+aXUdRIlQq5jy
tMvwb1ipnzFBx4M7LJqnTiFXdAKmhwFEzfkIQ9x0OkptW8E5z+6cs40i7CHghXCWDj1tMcGlk023
DHl8Ev/7y/W3tuEjuU+h6+oLrhwk+6M5mYOEoeqo06842L48U9cXVAqCdNRkIxKmNfMI8I0eLPZ6
527gY7rlP+vUUdVBMwSB0NbpY6x853DPcaUm4NYEeJjOneXm/D4G6U0MLnCJhNh4gRdN2LT1yEiz
7hKC74xLGv/YfKADLiWOmw5USV6sfQ+vtjd/8zctRvpQgVm4UAadaFsBkfiHNG/BVosiQL997zYb
xXkbETtTDYY9GbENyi9v4QAbSYFM2t2yNWasVoY1dadl7uCpAOucmDVgoD2XDVZcRoodhsYnzohb
meYWOMvxfnfRfnhw/SGc4KAG6d4+tWvwx1vPAZ3CDhx5v/+ZNKiQkwQ0rjA1MbvulVusMkFN1TKo
+XRves4zB0zGsAkux5MMU2SaKhsw9PTqkqUgrlvg0UAYMTQg+SrjiYbyplF235jjS9CqF8470Oaa
mD6C/AKgZ750dD+qC0OA5e2ucO2Ai1TmIlPGf5oV6lPYVc9mG7uoO2uHwRut0jTt+TtixiL1PLFP
QNqY4iyEpayMpkUq1DhB0R4yy1EggN5ModCD5oteHM8EmOzOIp+KUhScCENYh199PMvmb7tA5Iqc
T3DE1Fslrq8v0mrrPBK63gHpLYuiTIwEDy0hZQKgCie9ETXK8bebp53GxI545sRqD6dpFAUDofZc
ZdFUPXOzfsAJNoxwq6POk9gQdEe6ngG4nEGwFs0FeEkhztyxjp1gj8K9yzI/CIUoLwd7rNLego13
JhTqs1fpNRYv6XDywHM6WDyZ70ZP3sJg93pOG2dPFc3XiPIDCYMpwilm8KsXoJyATYEPgt2TeHKj
t2sfYrW9cWNAE6fwCSgv016sfOoxY/S9Mui9GINrXz8LLdyOfgcXTWzzzG6qC8K5rswD2cZaKtNa
gKDArcCTfhu9jXfLuLmAbphzlnH/AgjYNjU4aPEIMXYkeadhWIlXFJ6qB4GKyQb5fP+gaT1KVR9r
BE5P+IBydbhj6oLvmHwWjxrHW9QM0WgqWQ//HXy7h1ibisZFJHuet3K02L7G5180VOpIGjhH6ErU
7EUI7FPITnAvhDudUueWWsygBcLETDUpaOGwXKWMiuCdAZY8h48jvJKN1LZXEYj41fYWNE/y7wUX
uusJLJ8Lxaj061EVpouC98BxT4va2SfymKA4+khZa1g0vu0YSxY7GsWc3vuOewawlXz9vZ1nLuTk
KvuQWBRMEfF5BGlZAABXkGSR2EN1u6PEUB/ZySbEf389nY5jvbVeK2/1pmNX3yZ0fiHUEp55hpaT
6FVQoUacEl64ngA85d7KU6KLE3L8sI3CKtYl4s/dsE4vM2UnrOSuEBNAoljdAUUWDZs/NJGteunE
BxEMfBBMUNwv8meIUITK54mBlEY806t9liNd9/MekRDmYASX5FOufojy6GbAgELHuHi7hSkNU/Vb
uP4/h6GwCoYqdX3lHG/nXP3gkaSJt5gbRm9uMiBKSpd7y5U561WHmIarp76CRaGvMIJIAovEgATC
0236U3QyS3zOELSa7Xq9UjrBVf8hkmYaJfoj4vfxZsxGPzAn4sAS5+cJMpNd7mG5simhaPWJfCAF
NGr+7mKhUCi56tXDdAt5IqSilkKHpfqJStTUomEV8gRaerOgOGdOR6r0JU6T0rUZhZbiAT8W0r8M
wc950CDelOcLu6BhIo3MWLftlLm1uZi/VNbFecPKc8DkGarOsoFF2wYU3NnxFEuHwu4mr5tRMCAN
fUfDK0n2XY94mw1il1sbrtF+U5UIQ8RDHC9tcKUF5SXP9E5IiZ3tEMVkuEyhCtJQl8SiQDcKEB1c
FJsbERg0MBVRXgqIg17yk1l4dqGhbaCn+2M0qnwqAR15wy39fkK8mnDEFzwb2QI2ZRzu5guMJ2c8
oZI2nZ0g9yxclbIQs0rzbiOc1w2V+hTe+LOGVNcHb8dVDBZ93nlOqO3vRy0SreN7up/0KdrVlBtV
5STD0dMPxV06gRxIaIU8noueOgAZjtxNJfWmgScyXiAfgZr85fOdrRKY4gVkZYQaF78ajfXLAD7f
8iptyauR0KfcDqjrH5NcMDdL+aoPaLyHx4Kioh750Ur1mnztvOnWxAZU+3gwitHILDyGoQbtvL3o
jLAWqtxX2XykM+XNnvbyP3wJdKPBqZYgUF+/aSLRhd1eSyoOn+EqwEKv8844pCkrN9GP1HYDQs8j
zKXmWBKrtUrxCrPlbgGyRkQW5qy8crjZV04zH1g7EFtiJf1K1MmNN99YeRHIQrbduoN1T/wrfqpa
p1c2mYZn7vvHy8tnrRhrAFB2A6zw78+kHd+m/zYEhPKIpaiZKkLWJ5gtgXubbVYhcPtJN6QcJMUD
8oAIPASLIctMd1rSms/inZleQhbr3ufzDCRMLMtZ/bYelL7BbwcRhd2iR4C2w33Ei5oCnrrBOZJ3
DtbwA91pstcroHUcX0vsefbEVoFudIej+qKK8MMrFChr0AmgTpo0PYAKKhW6Lc+D0evC+/NLTGfk
s83pZtwDT0axbzfByvwbBWXHIm16oZ9RKrANVbHNhVDQDtoN7gKesoAHn7u6cpb5Xwrq5VLne20h
vJVVg8NUYdbd7O5JC5PTjDE6ZNhWXwsp6ir2bqO894vnmpK9qSSK1//1LcbUCkQjGCjsBSOFZ1VI
ve2T/m1LY2VGTIV2bLp081bzKt8+be/mnkB6LXUb5IgULLC6VxpXqQZ8NvdK5+GceqBdfu5RdgES
o2BSIhkY5WbZa4uKhn6KnUKqzaIaR4wxK376/ZtKnV0FmtQHyh9MRXMZJZZqVvr6B8m1Y1015Tzp
p9Kr+q8eF9W5yQ5xSpmtcZHXEV0eRHLuKq0hkjKPCSlzPt5EPq0h+ARmdb52+s2SiT3SS7PnBOcJ
qtMR0v1WafKsOhihkOfio6uf73Ok9MuKWLyu1qZyV6MNM6flSlVkCY0EFA97r64cQjlDz9NHODu0
h7hvCt7hC0EFR/dP49/BfnYQzhJfG+MLztCg9w9CwpzJ0yxlWMwGZWIhOPZCiScO2ZX/crhbxSJs
Q5g70nsdkATW1GEAlokNRLAyjQHbEBudQTxqaVlHZ0TNqR+JBDh2TesbshSrTdI7gvzFQZipMzkL
8Q/s2byNAxtXZzdwuW++5cxkLCCPBpaA1o4mpGm0N27/YtQSr13MzOAHXHVJJ3Bo74iROkVE1aBw
561Ofzqqay2//F93+6ALPQ8Z3tvEnKh2kc0ta8e8XBwtvoSWdceceuIfzs7Eni4rMms36T3vniHS
AnKAgOxIjPYB+yn4Nqq6YsHXaniMytM8HGcRYN08u6rBAHKGDB4Vbjckc825KeI0yPbVVgvpQwuW
E+tVmkuQX4gZlOtW4TorlZEQXEU7BkDwEuDz8ybJjKUmmYCgNN0BPiL+Wc1XicL+RlVO8eKo2/Yr
vdPrIhYPEAHPXrPQcfEU5aasyM7kdt8+r4T/3hDugEUM2iuiJs/eSO9C/ECSyT+ofJhw/CmzqPlv
n6FbIX8r6UI0fpacTlsHAdSq+fzMedE2xEa5AQZc6Nkwbnp4951CRdCIEboeOXTFYFm0OtRASc+4
5dw03SyUlvOgvT2gcmfkiVq9nxQkWyT8WgIFS+wlYAOfN5xJL2Mc3IXZ7rpRfgznmkE5IupugWR6
auRIFzm4jhJD7LoJA3SJVhpGV/iELjGolLU5f3As0BXjS9deAq1tianMeg9GLOqjhh1vIZASdUPG
qJ1p8hi1ffZVPvQNpBLzQvo2AZqpuBIQPm0XvWJpuXWodddNfw2DITsrpz39wiVdBxdbiCwVpPux
Kcxn2E097EmqvGO+69SLg3CY2vlyFuovSJAc09wXi2PlbqrKhKzCEOX2/STTGoGrvYAHdHQ9RK6S
Oyf5gt+wXWYng4WrARAtVBF9xIUCBgt4axNDJeYbACY/shsHk+kDa3PiRScOml0EQUfPIo19Pby1
0n9DtoevMki7ExB2s+bMNSpBdHLr329D1UBKrjU+R3MXmruOC2oHbx2lmZDOqFwlqiBiqo5toZtH
izdgXpMNpdlcNU9LU25R554sJ7Zx8irrLOb/A0ETyS/9w0DRmOUNj6XLLFK4Tv+dB6B4+NZevnV+
78BmNexw91I3GAQC3ICuRBlRLAm+U+cEEAYvlWYFxk/7wVyp6Jyn3C7o/AS1fW6y3KHl9Gtc6uo6
3KDmwcvZn/zgd7fUeqrOppLnjqY6Rscs2vR3SGrt8n9BGOdyiuGjJfzQl+tL/Vc36GJ11FT11mxN
TjTe2W2sOt1dJonmf7eanFJsrhOPnYgWbRKdWzdcbFrupy0FtGfM19kSTQZhzTeaPwYETr3xBPA8
VrnU1Gsq+Y/aGWKYEGXj+JdqyUrIXnkovv9BTSrhWL5unpEo6AEWOL2k+XLRCyQdVTfA9CLqC+aH
xIs9SOtLIl4BXIu+mUmjm/Sm9vF7TbSJLZ19KqWfZMbfZ1gwqY0JsDLoumY35dqherMjxk38ZJ7V
fuNT/ecHP5mySP5ACroGP+/jomq/7SWFZtlAuPXv0rcQHfpSzdjk5TdKqPlDKWlgA1sECxiKW+p1
dgbScdIKznaOSvbMBh4qoQlCo8tN53dnv7hdOVwhGtlV0/9aHar0ms5CtTERdAjNV+ZSRiQJt0+X
Du/ye+HdvRLS3M+8CsmPz0xus0ihXVQNj7xb0q/WVFqn9dSVEiJ4TEYTBbdcnl+xz316g2IGxcsw
lDe1+LbR0xSllnnQrQJTLe0QxK/LXXuSTd8oZVEu5a2ZuPDIy8kZlY+acmLau/x5f95rV7Lq40uo
3Fjna7RYZfXxpwK5qBCjuGUdc7r0AGEefTMuhvfCjGZCED/RFYN0UHGeKzPoT7PK+6/qJujKF2lc
f5wzIMrFTOWXXAp4bNPtk1gzgeAKL6yRYw1aw4Wo05UOK+876Al/YTdxUGpRQpss4xUqxWzDBpmk
V1LAtlDjwfY+ZEI+NnLIN9GxdweiowZV2SBqD3elA+xYfDIwptFw7Qk2xSBaUbH7O+jJBgRqb7Cs
qNf7o8L75k9LTZG/rM4ffzx+mXXbnLvaq9wv109uVYSATbiGHAuW5xsIluQNERJIJxkCS+wHe24h
WDBIIL/l6foF3cOIXMDP13yCct6lttUFz5MaKSUD60UYpuZeCHZYvhZO/Sfv0P+gMXDGqEX5sj+y
pKoUzVka8yNGJcxr4AEzfrZFelA6OUK1gO1CbjzwzGSxPqPi8IBn8NeyetVrzOCQrq7IH6KPdRFj
/QdVsTa1SSuy9ZlDJE5CIFP8CBAAvd+t/tMsJ5VobXgDRlys7NOWgtMMIKXAp1sFtBOGVjW6CLVH
uIjcnyG/bu6Zg/EApo2s7v1nE1Z7u6xLk8JRmhWR49HrjP039FQd3X6kud8Vz3ZBd0+cJ5QmdUNv
buIyVA5fEiswkI9DrDtyfiuMMPrGzUejtNLuD9+NNAXm9rNiItk8EL8v56rnH1W/L1LEE6oz697D
oSDqio83RrRo7S1mxX2zPY4+6nqJGbb+Nr4+Ep7PMneEf2ZJYXnDUWoqfGfZvjsvK7us2w8K0Ew2
1HaKQG6Hq+4Gal+CCGEwNsRfhfAwymdQMbie0sf/E1Dt8M7viQLuVfLf8W7V/JjpvTpKaVBcDXOE
xIwJ4Rx0TgBkGc/gHF7JZehIHPTmfvwkjGq6oapxP6M+WLw2s+NEjdkJPL/soFr2FrOW8yqnWEP4
oSR7em9fh63uzEBwU61j8Z7w7lwdw4cB9Q1PJ46d5+EEm+jERKvW/FJ9n+DoKaS8KSgj/oiqwS8p
RSAH1bZ7AQDv69+V3BBOhurxDc03i4bBrBYFogMnFsrlVyQFJ6LPtY6kCrF1wkPO+kmgiKnpacDw
qnruJKtJQ8G1wIfenN1+6WQfvywDiXirf4dPiAUuECpJ4WGrCFrHkY3gS9xHTE2LSo+AvwX5wB+B
TkhWBDLuey7lmRxqxaCcgWcKU2VVBbPFYUZVEbwZesms9jhtG3QoSvegUh05LCKBRDAyMNDzCuvy
gL5Mv9HYrXZYHh+RuT9HdEqhW8kzRwrRqeheUhrV/umNytiIcMx+Z0cwV0atmcBIjocLHITD8OIy
r0nh+HB1mTmZmBJnptDnq5VM7NXs0ysWhYz5tUFR1jAkHC83rnIowPb/hyIPeRhzxZPsqaXQeKug
q5hFVm+V5QFjw9SxF/OL2zGtWkrElWO1vkcwhRm216K4GSCNVsC4812xMs9k4YSBU4E+YQdMQ7qK
M0DHui6iCFy+YJQBk8o0ePmqkOxVz2KCcgnYeRSHjfBHqG5ufRi7WFDgZ3uIJyd9CnZdQzqffQ2s
6PQ9QuIC0FZe02GmmycaOenNHucijGs4VsNNT/gROltWreBLL0s4p184kt70t5S54Z/Nzt3pZ0m6
Ai33En9ci5ubu2H4v23w5dPR1k7lx68M2iwzLDlAL6dEQgoH6sfHgodjGIQSnKKt07MXQlD3UABZ
tx/OP+5j43aPKfKiNq8coLDrbqGaZxQ55tImdC8RUxopm9qTqnpnCopGsdHBoQJaxIgwWtNJSFv4
T/WzEVkneNtVf4zreZ7KlTA6Lwqu5ZnyieqJWzlXzIUJq2DDdAHEe5R29QUaaM1Ug1rq1ZwhUKOs
XbJeqbAxUDNcx03ImEg6K/1svsZ3FKotPbr0Cp8tLETLVXDfbl5CSeo6oB0RmT79eljJ6/HlxqWQ
MPd2NvH1f63O5O7zXi9hKOHl77RPS4UwsEC0kxdNJblvT2s3hiLbex0gUyzVDk2zlZumoORCtjhq
gtj+ZD4oge452DWR74masnvb4UeLtUdqUF+ztbwHE9YvSe7etBoSCPbF9uSTgADf011zkSkoLbrG
qcM5AS85NDY+sWrcCjC48ntV55lwS8MByENP5FE8ZqE2saO8hcNcJP9MbxYhEAztnMjvn9wp0LiM
Aa5SVRBBBt/DKXrxQ1d07taqktoZfYahwjIXLC80KfUKP3EBC+ZgzI84ak5GrGj1GwEt9ZESa5o9
cv3F00JIl1L3RraD5e3gJq2NUIKEHpbTInrYFQeBl2LlQQ6Qnm78z799FYA4FGJ8Sn7y2B6xb3qg
ADVnGaBWZ/NilkjnNAKRPnpnBpvusn6B+u0ZUT2/1XqJ5Lc5Ae2eRpw06b2eK46cxIxb0Au+wpze
tF81r4IaO0DShuxDYuhKV84Y4pSOF2LIRhSidcm39j84xxYaN8QaEss8lPeDMdQUZF4ma85/bRH7
7kff8LGMScrsorxE81YUnFcxu34WpUYIdHngqPBkmbzkzJedu+13mdUQwBmO8oHBsCvUYO5DCCXc
X+qlteUihyy0koUCqAtxysEk+pfxhstqmHaENZk3e8jlpgtYmVUaq1xXS7q4Q5Ms38ZhEGBNzgEk
R9gFxR8/MQdC75IOqfbo1bFWAZ/ZNXdhqcksBpWFKHAuh+4TLqUd1+2+qOp/v2dUgVfxROUc8ia4
CVq7xRCKnXqraBiGQ/uA3mHeWqfMEuEGeiUATGuIW6gXBFYaJtQgZNNcakUnfIzjXngwEL+nsr/8
0KiH++wl0WyDkgND/hihi3IPJfV9DrFuKzHq5d/mV0PDyiMSWWQCW4LtwOmZ1EsPBdMcxQ8K3k5r
yFLhJCVBFP66Wu5qNPwj8mvFz5EY8T7ky4nprC+bNzT4blFHDTU+WLvKvSZaOHmjAVumBwKY8/Mm
LHlrSpfTfGn8O5SETQz6P0B6xUKn8BMgjB+E1020PP4gjE9cmKKM2Q4vrD3dzS9P0m2GzlWY4NNU
vNAdFDAAIZQ6WHpldpJgNUDACtheDeg+05ry0fTBFdrnX7rC9fQGg0rDrRkbGqsG4V3i4Ymw6EL9
AFnnaEXb0+clqv3uB/MoWcWt6RgaOsP57nNeM2Z+4WLhyOdRmXQI1q1rz1uUnMytfNMhQ20SDqul
Ma4zIa+qwSrPsP5qTTyEzQiY+vWdTUR85qIJTebGm/NhVvmsiBWzvIbhx8+2GaaMhsb2ZMDZI02X
M6EUq0UsOqYjQAd3vZFeSuo29CjRsStl1q5bZDR3sVZHgY5ri91P/dfD/+FKtWg+b6IrozpDEjtb
3nlYVU73aYpaAtSd/LDIOsfhMaRTKUl6xWBHZMyYhbI0mK5ib3Cu0fxFUl15fyMfiiIh8nFsU5k2
GEJtqTy9RPAYe0BVdF17dkyiKNa2+Zsc9Y8P/xOpYWtiWlpPDheDdzdpfqXlprjkEnSERoOnI+cy
5o4qkM8aKATv76xNNdPSk1Sn1hqGE3xgzuN+SpSBNPiLaX4/7NF+l1GTmvTotBCoIdNzE/weyeJX
PeWbqQHUKJtaucVa5bLdgQ5mVwY4pJMNBo49+yIZ0U3eJt6AWZji6oZmxUefps7YPnRX2NIlcRTX
jk4hYDauuzMQrJ36eEHmrQ1FZP/uUyJtVJmw6y5OvxR5mnSnDEUB/ZcZf2XS9v7MhfxXlQF4nQpZ
lDJ74rGHCRm1sd6SXA7mK1QHeuTDVxJn4bD6UguXQ4fy//j21rW2zs3m+Wx0tbXMTq8JSsqJx3CJ
H8BcaqB9Q4TyrMuLilFm96hkUFNA9nrY6JEoQlkt+a5nUofxDVQ/ciKwRIN+NOdC+WxPdJR+wb8m
rtsD9W2NZ/6VnErYO5pMaM/dx9Khb1RlDA6aL1nIME6NsMtDNMRPJ2lZZk4reQyYW+nU4gvFtu1G
q42RFKyH5HRKmLk4a9X4LvpHds/uLMd7cz3RPfbCm56emqbADbGOrejK7nM+8UxPu1M61p3jZpSt
oSN4hR3EFewx9XRB4Xu1+koSs3MQ48xe8XBiEce+xhArO1fNq1sIGl60c2dmPO0tUwVhltZimrwY
zbO6gLeDae4yX2cK1xVpoJDkKszXhDL6UDiftjJSd/xo2OtYHYY0PUHaH0KlOFnLjKNGni1slKRt
wYlTXmrD2vAyyyPWAk1gUQEVoGZjd0CBHrZI0KqNsQLKNxbRfFCE03RBU4/6fpSpw3zmVigF6mFS
aB7r8ZGFbg5zdIXoUpa/PreaNzEgGdNRuZh46YpCfPvNM/xy+OrzqkgcavlAqtu5HMjjIvSUuPQj
QJEULAhj5CpSfKf24f8QqihnI4ZGYZ7NLbWpn9l5YOzeZ61p778y2Ojht0PC9fVkL0idwMfMpo6l
oOh0jpCFfXlUKXUDbdjE9W+04BXC2KevvKI5yFrulbCLlhJ3LfnxF1VgQVmm8GRksSx8rF1TqXbc
xGWdKAkgibFBf3/zYme+obuT7x34FdvqTaqVK1toTuAJOdtRegoSMe/CvKBgE3cDExOaWCQPkoJp
wAAM8X8oQvspOcmSiSB2SHd7S1ysNsb2N+Xu9vwhhOKtMpaHYwcgdrvfD9Ww6nFvYyzecJueHmPP
gAjprEoxCrg9sNC7Ig/7IsP0Su9VpIZsmkcSTgaL3ONLWMsC+5NjCaw7rONDNB60U5LDE+geZcAc
RT5k3A1rgkuVSkqJDo+bSOZ44MbOG4zizXm2LfzgDqQWVEFbQKQ4dorTyiGVSmNlC0GANTinHhja
CN7eRZOpb+v5L882YjhiNDI1uGHP9r3mLZL4DYp8+NafWVnGCxqXhVjdp0a88sUtmgJVUUW/z3Fa
J9Fzj7JaB5OBRizzbndWMf2ZHGIh9EUyzzBFFWa4yJZiLbURlgwlt0iN5Exk713q7ftEeEgBaNwF
XQIyF1tQ6puJHr8mlDBGBWyOTKMIbbEGAUuPqJOnrJ3DaFfK6/YnlHdj7p/d2k2zDAXU2/rgYdK6
hwhViVBxZP02879r78uEYmLEq+YsyuFSiCdqjmGTtcFWr5y/3RRHZ9r/7X/4tomxxCwC70I4046A
1vVoVO8j2EKC9G/jvv6u1odIU47Kluz+roRNTJ+XL2D+vOjjMPNEt2JqEfLtn8RXVW17G9/K1KmZ
Q10CkYWEDGag2ulXmgbaAdwWQhoUS9b/aJoZ0F2DUZ3ZXtT6+7x+Tf9kSZ6/NYH6Hos/GLFg5AkG
TWjPalz0h+ot0rRmC73kuM5hfuBh/EdWVLtooNKV8Uqbp6MVMFdWbxrhPr0etNOYfUw2C7L7HF4I
23DxE/NJc+f4ThZL7HfSn8tLxwADvpsTH2cQjDV86AasbUEIO/MvtwApm0XBkZj5fHf7QjZZfjfB
5WaNj33bbaFp3DjF/DcLvWyHZIRVUyN2rHQgu4XsnrD37/XNV4W9Mi7wXTfPRf8yd0D1ECf90VQ0
HvhBV2Iz2n/SJGWn/SEenbW7GzG/jfcW4ICb5/7AYA36j4Pkxk1Aho5V/Ypys8FngQ+rlB4L6/Xn
1mcuqpsYx9Id9eRM48HVP3xJkYQ/m1J3GHEGO4kAL/oO88H9/PWUPbiaH5fYSLrtPKqrkiUZ3KGH
zVcIeCfTPA29xjgo0EdqUBnv01bRYiPyeD2j4onHITcFy4n1Ys5B46SssPooyqXTkhEfSqMQZ5Q3
udWSewxPlBxikyp0sc/wtMkyG5ku8B93AYQmOUh114V7asBKeXQcyd9WcoflT7nDi9BenI9Ak8sK
eS/njnfsnJ+Wq+WNxbWyJV6DsjcIgDeqPSYPHRn9YWbsQz487IleFh3yig45W1jRP0KzIUIVikr+
+h+4c3kmwE0wgmXsC1pAw0DePjSDiavPDie3ZPHx6+VB7NtUX6Zc8f0FADsK17sLKAjkKBRM/lPL
0kYm4hpa9Na1M6vQP0Rx8iFQOWwqBoXKxj6JefvNCwJYFH6G71y06Uirj534YuCUGOzEaBg+cZrG
YKwe4OlIueD/KebPIi0r9nVx44eyofhRBfWuBjNfD22O/hmJ23vLMoRUi98nzJFTyw4m98zrZxWz
6SXsOkjjel3Lui+A6DRBAbi5qJn7bNUpls/jCwu+Mq+77WzWsJbODIWYRAeoJkQdgTam/GvlBuiv
g/fkvPxvDGvULLS49tZiw2384izRXxa4hX36C2H1TsXfhXvv2nti2EEVkCs+A2epfgUdZIbCwrKY
iN6vMIM5BmpOr3ou123rBB8QFCjezc9yncB6fxCshzFL+06un+z6OmoZhBSD3tms+3mr/yl4juvk
SERx7NFAhRJp0M3JP2/KV3D/LN9SXwSPxupk+chLYNmu7XWKIPFkLDUyLi77QyW3km/v1dCDwEya
QTVM1ctvhs/mevLxgPwxbJUDHNCS3ak7qJ4SRwasABBUTuHZ0/7TH5h58u56qMNKkEpI9B6R4yaX
Kl+HZR/DDdhJA0sRDcrcWtsJKEryF8a7cDl6ZV9mfAQ89aglUPf6WyJWxDv4UD2Et6P1qYoEhFIA
2ZqT2Y17v759oGTBAfiXtHf3KjckzpewLemHGpvgcaR3cPzuVP/IGpKMHcTL5xC0cv7/aa37aDD5
0MS6WR9sWFXPskfm3OFdbaQTAstf0lB0Zr78JNZYoOOOWtgjxz7xBqMmoNnhyK5xW/BT8XafsNRb
WMWNNNtie6PnjYja+O5JHYUqyhrCL8zrqEj8YEGjo0C1H6WVcvP+Q8F4twPEnbM8S0NdVpgYgl+J
pmHp6qPCbCgrodlB0qbMHBxP8AKiPmXsKV4z469N650MsMpgFtvIBoQcXE7EaWobebYhFBq2EVnX
9JJbADWTlRliM0NTLwcZ8WEbhsz9EalaVgJ09VIdEAIFu677WaS/nkhtDCJ2evqX9dbdtHt5+7Z/
UGH6yUuKBYgotxIT7DBHvRwUMp17lBPPWMZG7Qk7KtcVt9TPUuArgOhF90NUVqO76a3D2DsyFYtq
XAa2f8OYHGy3QKnLnvsUghjRGRYKWBDVRe56oZyq46hK2Kc8GCMUhPvpu+PuoAhls1SCwK3mrzPU
loreQU0HRtPxz+65VqV21JxGCopci0wkqRLirddLgJcWmWxAHxOBATk6bIXk2gyHvFJtnTKLaVyx
UoNouh7kYU9MkqE2xSi06U8tpgcQ1T2BCElCAk0iGoZ+VECTlrwDxzM/J+5oGO9VvvHfYfqW1pRS
RtDv6tqpHbnVfFlXicBvtiahHQg0B0r/lA7BUzid8XiIfaa7+AQhGJnyTlVO9KD9nNsSMVmy2iK7
zF3XRXcVhWhef4EFPL00zhvdsen/1w8fKBR/ouBLIrxGwMkvTziWfS+NSmKUZ/I+1jemiCXP9U0V
DJrgROlrMSBo6hQFqzw4xItoVza8gqVIeVO45/HbRxqSWhLdbv/CAJDpMM+UwlLJF41VwShdQ8Xm
IS5pAmnMiJYBBeuaabPkh2aY4NJaee4zc2icfHLpuhAhf07jKQ4epJMuTCKSZv24EfMLw3ym3gDz
3s4ycfGOGynQRRM64/8ucnJKxG/zbGe0tqQgfFPqFi8gYcoApR/a3bH0iXa6EEEErOCHTNyIssd9
ZiGlW0p92dGx69InfL1Q+i6mvPpsdIQYeRp7JsKZ72m+ufDO2fZVbRkos1EorTAXbszQwKP0B6oT
sonojB60bVup80XpbwgnYvrDZP+c4SFe73vEkpfodZfRaHOzJY7IdxpLsFfI8oUXIcnD9JZbyJwg
A+81zcIhQbYw0tlE48EeUuUGP/GZAMuwH43DQIar77APQfFJDqLk5SKw+fd6wYEAV60t67ctRn7E
J5/cfHTN16IEro67Pzwg8IO9NF74o70coNENlKwHO0Ru2M+u416zeVOh7shCn5pifNxSYJtyGTUN
6sQ56y0LOf8a9v1JdyZZMMDo+SSFIEejzegwg5eHpjBJyljUh6DsM0n28sYBYFsyaKWyYGgLtb4Q
dXn4sh63ZEBIA4JV0VVqNolw+O/aZxrQ9HnqZ1BJcM3waoaLIBWgyCHKcGngxQvxm1IN32ui4o7d
fy3lr6A4i0TRSEiekKWmzcPmvtOZg1PEF9cBWNI0G888oq9OpV5NEWFThfGaXmOlN35fMT90i+uj
bazFJrMTJvfE+w3wG8oY1OhKfSq1RzuTPcUJJ3fWYDzf3HCUlCeGWt94qh4ygAZqpbRXau6xp1iE
M8K/iMgbeDnF1vJStUjO8hlFcWeOZtBMQ2Aa3iC1NbqBjofLVWVjKWdgHJuK+0umXRWD5FYhgJdD
pcaJJtulxCDGAlBWgLkjzE5vU96lCM/wtule4x7eR3WfsD8Ido/9cR5gs7JVMo+MIZaU0WxSwgfR
snVBEh6wbjhVtSwSdBrt6hJbKSLV6W40iuD9OY7HzcRrKAs/hfPhDYtMgRurACi6mz0uxzS8dtMn
N8sVf9IiOCbwlaaOb7xlZvkAmoMXolWPqwglp0aLveFJpPzPOfOobFaECqMbt1eAyVVuL0Hr8+IK
viklNWNs4XrDDJXaAhyB2qvYt71eL/b/3nnnjusFOb6fob51CSzmnJzBS1z2fWIX2Is8O7cwRRbt
xjeg4vUBf6scgSEq6kmxvIuBq8LmmVRYop+4fDW7H9RzRDm0I5ZL5OBPp6xoVhbCq8pJy83a9wvS
VzWxL+dwB/yYRamzzsNKaYNqL+2uxgPhwNaQBvbUEaDvAVyb5fZv6wFcMVypzA7jity8e+8tHa2i
yhBf315ADpLXSFQXssRGnkwJGdujd3WObpg3d3ywQh//Cu9I7I2SYqpnY+QRmHKXtYI4gOuE54yl
DDEQWHI55CMZ9iCaa6IS7NcSnOJOhPrdZjlABf99Zg/hzufD7bs7qakUVSS6yxxqwRa0dKn+SQ5R
FQQSv0XLiBWdq65hLYOEE+epDv4F0zMiWjX0xK/YCOUH35D5aG/TGDQiHu30p106+kfT3xDCUNgO
SGAKLTYObI+GcviUT7tRK+Csmr7fhtYaz4ddwZfer66lkcQjf9Jx1LnsbkIyUq0jFdI7KN/h5h6H
L8/wQ0pmOVBICp9ph2fVjI7+POfqwWPcvG11V7E4Qs+kq6vpQHp/CMtW0+4yf3l7e+pKyg6aOcUc
SgyoxhacfKcMDiihn3QTuZytogdKIHDoYKrpetRkLpoAwU7WgnjNZ1kme6tLnplVsegDZsdSrisE
UagmptMKcMeDWQRPkyB1Ef+HP6Blu/78Avg4KfYfvryQk7WcnjzrWYDoSMZ0GM44divTf1RZ+3S1
DHJT/ZeRQt+LLkiYwpdr9tQwXcjZAz4cPbPOR4zdbWbQ9YoeTrQCsj877e98/Vdg/6PWLjI85P87
vyO+e5nOgkj3U6ccqP0ECjKauY2UIVrFDb8fFW5E8vRzpoCJCfqYxBo4XuLmz2Yz+UVhlAHUZUU7
8IY0dPv+fLeYkES0/MDESjuMx/DJS/2hleH31uuG0edUXYbtHAM6c25lBPqMRMGvc9IH+LaNuzRz
cKTT+5iq1aYy9ymaj/dqV2jeXNY5uS6sgQfGTsZDjj7hFGzRFPhvaDUlDdbYmRAun1b5/BdUfhQI
oB6fndqp7TjKi8sqga0JYtkQNTgbcZsIUEGMGq5Zg1NV+weU5dDYXKUVoi++owdcPogqgadwQnsQ
ILpKvfhaqgi9HpZEt8HgDkOfYuPQt7ssA2vVEagCUXWyHwrJaB52ehlG772vGaKwY8/ifj80JndG
U8+NJzHOphBpgY6JOE0qFuRuGvr0/Q+5bSU9yxv69WTYELFQ3dYHRYhhrgpo3G+k0KBpVw+A4esU
9W094Mb4Ukznsa1SRoTeT/ckaOx47XLqGk9aqJ2OeZa4/aMcSdlS4I/7N6y6P4IaljnJ0pft0YCo
0s4P43oF2LuYf1P1n0b2uGhcTOpS+W9jF46g5D3VPkFcSyJ1UzM3B95BhH5rhBAtPPSFnlAaVyUO
u0aCm0fCFoGdGrLrkHmDlqNNRDoBj0QZVG3aPCrru3zSvij4g04glMWGaj4l7Hv1LmBqQJcPcSgG
XcPq5Juo76256Rg8fk+RveKrFMB1hTNJS3VcimzNBtWL6+ZE+eBklaJXc9n4VKE3ROFLCchRgWvn
thiyoaQynnlIuWrsxzBW9yUWX0B34tGeKygvN1q5FDZMBfUbCZfdBWQ5KuEbzacjCI9flRv3ji68
H08HnNQ5DxLwStgkg84J/komA4V/p8hudj/TVgZa8MoalhQKTyunfoSMGMZcAtm8Jo67LrjX5RWd
YIadzQY6xWAIPk8KYsxVk6gwgHLT+U4TaeVfM13qkufjwLQ+qdV3wkSBPAanuzu2WOqifdfPZKYW
xIpPYlTQZR0GcW7+yMbyuwKNUEujaZ7hgPvso6Xghbe7NydklUv8xHILLHM1qu7amGPQ3Wz2rrx7
Q1JTFPrJf/LP4N+JaYaaS8MQa60aeRYFEnT+vsS0kjma9X+WklHJsWOkkmvIAzeH5HDaVd/V9yk6
CUeqleM9+Wxq66vmjZfrIgxYNJzkUrRyBISi6A0kZa7l7gjXMnKaaOklHy+srU3H/3SRHY9Icd/6
h8LvLgUu3rvZvEfS1Ww6aaSHbp7Y57C1qmCfDU4UUDZ5P0VPnWG9mDpzKdQoBoeaCl+OkVczfLIw
mJaH7GoSUfooGIp36cMDCfRuIbVPlWxbupo4b2wy4kMaTBMjxPVMt/Ffspr9/8FJWyB2Lqm5S74b
tU2R4yifzkgAZDOap96LGYsVgBf65y8tUxz3UK3o1z4SrCyqa8XpuMvWBgYc8HSjikUcQYFQJ8nC
EEDMOe3jgTwOQiJytKYvTO25XXDoGM4dO3fJ5SIeqdj9jtQNgQZluT+AVbDfBbDMDzmzM4I8qyBK
JZCgxdzf1XcNUUQJjVG9vB5IStLbFHToppGnzYI/ofgpHWCGzl94T11W8h3TIe4cjTjMfuzGg0ak
AIyzn2WtIg2qPP9sx9mZeHRaql162zxfLqqo5mNbgpAXo6NVSS8nzviZhq4Kt4EYxax8NaThVwLB
PyFXsIQUqq4MmELNG/QPElZyV3bxoH/AIgo9Jvv8fE08bLdcSdgA2Ko1UNPR5og0ZmI2nJYUBxu9
aPZ1iOYxpNcepMaeLmjxg4Rog8h1L0/OaTuJSZo42DQaQ2PSTL172f9u8bTcQztZprZz3hmbFTgY
OZgPbrlgjslwMc3M1nQjlxybjhanh5B2avjOXPO3Y1dqFMgP9bDI2DWUjThobFHQjrcSlUoNJfIa
02goD5IDKl43XEsZOzaR80UKpMCFkE6gLPlE/90CFY0Q0KpqOXBn0Cfwykjrgkh6pScU9nEDMe6V
GNjH6tQVU+7MUEUd3gumkEx5HgE8nNh5lzbBk8dmUEwC+0aaXzzDTrgR2HROyn0Q4Io8IWWEkzIK
LAWaHJkT8jy6xnlKEHzvTanmdiZPqeDZR8iq4t5dkhu/SMMB8lemfZNzKxiHdSrOVfyznfL7G6t+
B3xkZTwp8jd2KC1OUY1GIWFYvsYuaWG46fP8Xjb1PxFLx9MR74u4TKFUcGI5sDi1irtgR4xhaKNr
HNwO5znbewBtFgzGw6800LPyInlQFKAqOHcOZ3OHqV4UMIfMXgU2zXGQFvSIZx4HTcnlTgNOTsQi
kB+4oGZzoJN5NhT/jdvHfppPzjoHVqPeVJ3yIHN2XBdclRLuIJfhreJBv7s6h8rE9tB5WYz+5XVe
PIS7Ti5CTMmnCZZDbfM+VHdpuKEWhut/MJMe2cumJ3gSrUEvzp/4nTZ5vrUz7Hyf5YcJKGeCWN1Z
SHOsqnT+ihHQP/DXzEpEEGbb2OESMKI5X/9JtJktbzCGWKcRErudAj7ddohbfMmhsvfyshDZq2mC
qDBj/lNgAe2qhU38nzygCGJqAAcQWeFckxLyU1NrNpVCPFVtX2n1Ru9jlDxZiHqwmAgTcQgZpzVn
zj9ZLQprQhEsaIsktdSk5Uhmjo06lsm5kSfWWudPp3TeZoj2vJw+TCdXqlWktEH3eBub/zBe1C27
jJoMzlUtlhmHS+WMo8cwjWUPKxBK1e0WL+Vu2dMmCrkG+n6at7A2kBxudPcPHsFNtq3FdIcH5QvR
z1x//YYL+ZWhyE6dBRFP36z6zXKyQcJMCfV6cM0ekryj8MIgU7nZxjH/mQizRwBTbCHeFVwShAqU
f3EUMVoEGhcjmt/mAPWzCf4jmxYc7WoxNjf0uxJ4drU7JpOKzddqWuM1OjkojNu6LGaliJeQxmRi
H37VSbRSCHtXeGmFimB8OBtMwmmbE1RCSn+3FC6FjNozQMEdRyy8uq76TyJId6LQghzMXprsBm2O
JB4YV2HW8HRgU2MjMnUtLs9Vq1izvW9IEMo5ytWQCr4Uei/3FcpMlnZFV34oQNDczPJAwxG4gtBG
Kd60dSC0/ghmivz+XRzdNqNtnsiMR8gLaf8CI124LJaG5XYKTgSCdQeRmqhnvE/1RGz8a146WodG
hnZSdU9gRI8dyni736vj6lXk92IZcAIXionkhQ2YYX92qJBf2PHTvBeF9puuELo7HYSRBASxgclu
czaoa/z+xVOKz85LI5yOd4xAn3Rzx3+0oF//KaE17onR7GucMSxm8UmW79hLj0fp56NRBfTRXNp8
GwHr+rr5Tjbt+roRY0w/d0SmAMPXFZa6DiKmUwBZcWqc/2GWziKtdkkzmRXdGCdDqsZtommJS1o6
InmOKADiuWvwoEO/UZKhyUaB42ywwJml2w+3knw2No36AtdrElc/S7IOplqKNtYuiOxyFamOoC8v
g/L3oaxSSGjJAFW6KebsNiSQZfoSDhxDMYRk3XRIfzJcyI3anZJZFVzPQ6uXX2OeWmG6IlAMV0Tc
EOvnrOlmHpCA/6jJRamKEPHCo8mP+LyM93B5n1DwolD32xfuH0wGwH/Tx1H9A/YdRdFFDn2MVbNg
EBJxI8UiBEa9bSIxHlhxmge4MY7Og315MbaaJyrHebPD6QJnqn8n2ttCE3uACcxiSoTR09JtyjKo
ijqDErZ5gtVcR1TacODSSMVVw1yNEGuVu/TRNg8Ekv6lm+gxOi+SjCoUJxfDmk7AuQOxGvnS7iFb
Ue6fRZ2Yk/zQm4rOylzHMMZ5U/bPDmy0JhGDG+UtbNX49saU3K/ig9wL6VfdDLEf/eDoibwtqGJ2
2NOB0YCeAxZgkDCMVLkEzAivBdZUxd9e736A0PbNsLnVlpyewPjTjGPyTeqv0+ZXqVrrsL/CGRU2
1ymROq3R98cFRPTI1BsjTsbLtPJ7zHO50urNyVSXV0GYU5ddmtUVtbQCHaBaj7Q/drlSCKVteO0p
DeC/hm65xYIJ0AXC0a33LyEYaGn1h/LixH60cU09W+3bfYq3N70jyFg3QmlpqMjLMvCMOVXuSNFr
+PCx3SpZP876WDjP2nfT0aow8ym/mrgdmFVnU0HmDZfFvBnzebyE6JlHkXKmf112+OKD02gJWcaY
HwUOlU3oe/pSHJO79zefHSpCbi4geY8xLbvAkrP5KIMntK4+o4Ia2DT0eEaUHcUmVcYNIMI+jAXO
+Q8Z9e1RxzIo4EhXvzsbAc+cWMf0+4vRq484b6Sdd743Ze+aQicWeLYvT2YLX9ISTKBrJiHCpJGi
4ZnqXDnkQTPKuArC9I5gy0gWwyIvBTHVvClgvxD/41lyJ1T/mQlVUdQstQM4z7EaPjrvxAumeSFu
64nTkn0wT+CzTjmihYMhJGfOa/Uh4ILnEFJ8BGPBjsKwty0+Qo35fbBuLywP/PycJ5xYGn8iraol
yfZ1DJ99/Wyt39/fKrvsY9bRR3Ui+yBvbYgfA9vSX2KBcUA4KO2hKezbuREqz7ldsSWhFQkp5F9y
cq0rLJNuYb6yb8oTQn/R2khL3R/6N32LyBuSR3iuX19AVzPzhfvO5b+XHk2SSIeXi132+RMGpZXh
6mF5rlQM4kfy/VCpUR63Cy8ECg89nAKtW+goYBvsek6WPni4U358NXDS3+UMENbc7GnI6wT3Uh5C
WzkdXJEbElUrDiYFRrP9tQk9FnKHmDpO/P83/dkOhFxfQfxP8xTTa9eIZICj4MUAI3fariYHEDTY
9X1Cv6ht1hOEUMVxgahAeBOKc0/FTtAmPUTRWvNhtRxMbxFd1MllPGVItcrfQVEUDyzFECH0MCvv
0emK9BY6LgZhYDwYqhdyJs751Y7tuKVMI5CtTRkSdEn/gYxTUvwdJoDRyttBXtIgGXOylF3HaRSJ
djurcOLFnwCqNXVmDogcHAqT7YN/nFb1Poqy+XBY39ZHAPUSuN7YvZzcm9MaEgh7L2kOweLUjCmD
g3eR8v41uSeqFkUeHHy0CTjmrZYd5sWmSnWVN57pXdmiJ1YGdfCKTyM4IqFIyaoIAF0w7sP0Hs3y
ShN0McvlQq4Ucpo4AA+3lb+Ca+KNR5wDk3ZyWYdMyca0VdMn5XCmnhyXqeTp1xy1k+cyjBhNunjI
0psyYXyTSnsQ59nJXOwMjqrou6Tm9KR8bC0dSBzMv4sNYDMoB48uQNFvcQaUreUOOaim7QidR0Eg
K8jCvsoP61frD20TFxWGHI92U7Zth5EqxbfcLMjfMDucSC0ChROi0+CqfeTgVl/7lTg9oP+PTvaS
4xJJia8gO2Y8ZEFyOXaL603c3y685LZusaHPX1T2ZdlDjhVvNmF4yJ36lWCCqQw6blboe/wsIS4w
xbAFXQPhKD2pfKySFoojj4qcYqWuB9mwNQEsGGJpmyqcrnyKmw9+M91v/ESjqQpPLanoeCH1VeWI
652JTlvftlrOAGTUitngRMwgqiRDkbbDdOcA1eaG3VeihSk0GVokjFNXIJD8iJMMYHPuGAhyNFRm
dDZwkVCOTh0qBBaUonFI8d51olCa1XeeOb1kam1R81kE2RNZemsr2IfikgmVba4K1iT3cyK7vUaq
uUrsT7w+2VsMJe7XFecTTLXs2yx1PIn7THBeRHEPdV/44ZnnIUnOaGh5RpEXJswDnlyyDDUjVboh
/Gm3sy9ojDPFQOTrpe4YMb6XXEZLr+XFvd4+2pYXlrfrYdv/umcA7XG/FGHWj32/9F/LpUPpLWE2
n1ehmBMyWrdBLBpCU2srBf7iYCkW2/3107GM3ms4SJ+X/0A21yQyslKCvfmx2q2sIaFpPXB56DlF
zPZkkj00deFaM+RY4RXG3lfnaFyA95qmOrcvdX301xt5Gy5IJuQ+OKHNcZ5tSJQpKXRxd8GxVZli
Lqxw1z3i+liNH9NZ/yluIxvYj7/ejnHyblic9WrGRp3wuUPxIV8vK3Nl3m3TsGcPO1joFOhbgM9D
cVUAdYqXBKzqnz1i4toluRvOyy1c7inhBf17cKaL0xTBjqBj3b6k13uw3l2PQTsf/KjZ1Js86V//
W+tzg8Fh/emwbJezk5OstltBlw+EFzLudehVhh+/xe110DH6HifcywUY1Pn3IEEQJBSbDIrKmyl1
Mm7SYl2hMSCJx3RZ5KRsD/VeabcOZmIpnIylTZUhEpI4iOM7dxn3gQ7rwpsvNgvoVHyLbHXokmzj
odo3Gnp9Z8EQvPln71Tz+HvY8lFKVITK1Uv5fm9TZkIgg+fX+n/qSdgZwxoKgOKOK/uUmbY8FG3M
ecBaMutNfaZuCAwm7FNw7qbSPaxMi85EOcALREFff9CdTap3hD0tqnZpv9HfxSkmuPh8/8GBiUdw
DusCEvF2fWU18MA35BuNITk4b/eLxJoX5tViNRjGmilgyRTHrGeUSzAQlUuWBc15e2h6TG4yvU86
xWnzwk6b+LmfSthpEB5YlG46VwmYDdkCxI5CL+oHY1em1DKHvTX53MESE+R5cuUjwSKM6tjrTAe1
bii2b3pscVJt43Es7PX7fdezT6ESo//PYwGdpiWEm9dc3RdqhPEfyEwKzBx7huKGEC65Bdk6EdCt
D90VkA60JkYs3a5WIguci6+uoexpZ4uz3rTAFR6As58guwAgUOEZA2RHiud5itFp2Dd3RGTbFqy9
MDdKTFKAU6awdxe+wCcrny5lRDAuaQDGiNt8RxsA3rGlITZUgI9Lhba8Yp1uuhz+YTQ2IGnwpWhs
nDX8ezALArQwOHbwnhMCcqUQKI/ideTmYx6gXzHgf5wwqmqxMBvOHTzjtY+KBFSLTJpD+4w8AxTA
PNhIld413sWMuMjKFieXhBnDY5gbK8T32j759tlLN51VxSA9yxsjaYcGO+p/QxykTIsffvYCyA4U
yY0duqtqrtGhM7JUA2EiFGk2KRVAyeTgiIimJlMNo3dC146yOpiZOiq99+0VWPsD5BqvmFN2olEv
+jn1zIcinWBzRvHvF9NLbD6NmM0VvwtKZ9StF5cBEgPumys2uYVirYPSE9z0eHbmOgT/2hcGg8eL
O2Y8iaKEV8Jw6DVSxqFDmQvo2KL+m08sDKyCtoAolATrdiO7A1jctWv/Lf2Ik0QXr6+5Y8ecN+4V
bPQdvoIDI6uQLm4rPFZliKc7HHkXgA+VlvXpk6XcsDmn+4sG51VkUHVrIsx3bDS+pnoO77gPNosv
4rqSeQj51GmNafYMM98oiCDR+2qhrAMGEAhllu904ZVKDNXKbO7LYLEU5mUqQbjwF3A4tkeXsdje
HvYkidFazFE+2d8veaKtIMjw1hDLB65bD4U2Jm26lUGj7jmq3vvYK6QCy2401UDw3nosSYnGm9uk
0ANtLzq7lHqX+mxWVtSr53XywDZxP9Rzi88QrfSbDbO4jvYRRrfhlkpcLqwydPe0a8/1burgqCxT
E+aI2JpbT/YZjvdhboVOzE4QNTHuKa8IfVjV2iH+ZigR69qQp3gPCJ/ElVP5k4VmG/16n8tx7oDy
QoGo89QyeXk8ertXFO+rEaAVDGuQALRYIdtsR0a6gSZQKivGGCY16raQpC4ttb1+wOqpYX8L5+Vt
tStCuE/hjdPJddzoMJqam8bC72/yZKm1IwCysGRBxhM8hbykwZMhhNO47JvYeB4J/XN/BYD9LeO1
K2RY9HsPFtMLHADxvAazUWINeXHURGUwaz/O4na43XnYCELZVO7v4kwo05HVs3OHygexnuWgrelI
23tSyJmFG5Md3/m7SUjXGeS/LrmefxG6mCjTAm1YRUXPhzMWw6MhZZTIW69lGglPhj2H9/FV1Ejv
ko/5Ny+KOlQq54hPYke8xRyPzDRj2EejbEvJfjfdWMOWNssK/NwTnaLfCTeWnfRhYNQ1ZGuKS8oO
rxlSMyc6BCD/tp7xh0ysFpuF7ude8UnhZNuPKzy7i/KHrR8KB+JItoGwxo80D+2ooX+2O1o4ptb+
hPMU40Kf4GypbkfyN3gucEGbI2RNsjAL28qHbSa+C3czpST4+CmjSBvSdU+dMwRnmsZOaSko7OBq
ht/iWws6FudE/geX0360c9dI1ZT5+U02yIJ2AB8AARQtlhabHAdvWKjHG+AXbm83+VfLcnrr7Ofh
r9KzR4wS5N+h5MxQOnrv11cBH1dkAN7nVnAK+uY2mIHISEQ1DuR0SW3oKSlW6JIic0XVNTKgzBjR
4tr1bjxPOY018IViFt4/3d/TwR+OsgzrFLKMgHeMh1nyxWlGEnIGWcxSqb+YRQOhmNxR11+48H7E
b9eB3uU6Bm8M2MSGgNFsGBdZDjM1/K/906/bFaC7T68yKKtm53IGeC6IhW2dRojG0FdvW+TXeWK3
0jw2G3Ypy/v/iBLYInOH3qQusqbgd0I2oM73RS1LO8btlbGHQFLmF9HyX6OWB57WaUnZn2cukVmB
75DkRdzWHi9gmC9e3td22hEf8InhxHucTUL/di79IaOlKBlvDN6NjWfh6089H5+t3gLZYSlFaQPG
qvDz7Tynqkq+pLvi9V3appnm4LBTFO4o2qNPAxM8zss/QlJTDfF71u1q1Z1ooNGAom32Zbm9RfET
3UOWhp+kVMl21QuWiHZcpWgU3tdXhgvABIhf2krJk75oHWENys8Ck9wiWAJsOFwPTBBPc7bE+bpE
A5SPFGCiUpdxgIRDN0w0DSxsQlzaoE2eSyjlFoBVJ2dDQcgngaLjBRYfCFFVpSnIbFNVpYpXP7u/
K+0+wzh5/Vrq9Uf5RI9vJ1Hlh497gNa2FtILYnVOA181U6tZz7USxFbTHfr+29JgW5cetI5bwVog
kcnafV9HSXn/dV+RAOCz5Cjm6nycoHenyN/m/ZJV6XlyI/qE3+coywwoPXeRTZVzUaOh/JjCXeot
3NTd5VtVOz1yePlnKWz8/QN3hAHrcFmeBS6uc/Sy0WsR7cJh6axyalMSj5sYHo12pOHy+ADt0BCt
hXPR2LBs68mAv0cBaXydRoi5s8jGydOQBAc17j0JDem5xsSZ5T8OXYJFjE24wrRMpTd4Nb9G1JQp
g2o3n8i+oXlJ0WI1pHypCgLyUHa0EzlfWbTNDsJS/jpA8ZPONOurIZ9gMmTEGDgGKAu8pvH7APvr
NLProzkai+PS7QyiF9LQN/OKcH2DIEYsw3t9tZz7ZWCKdg6XJlfTf9c6KweKSGM/ZWIcRxzH4wF4
lA8ghd52iWoGBOQpTHEAuo19xvaUUiLD4LBfQW8iOd7YTTMyiimThObbXjePEhQirvu5gFu3+Wps
nWxCPndqIoSnbLPlnz3iT8F4qL+2QO7ncWE1bOtIIJjSI14S+Im45ScMkEEfSo6ypWjFl3Y4JWvb
DMmq5YXQZXS714QBGVqg+FFe8iEcQs0ZptSTgNI0nLNAcrT/k6+VKv939qvEIakFNfgj+aP3NtMI
VtvbyLyc9t3UiIzz2ghgF60AT2wWcMR8GcCBnJSjIXWxZS5xwf1AjUsErd91Zfk5a6jXTQUReIwa
7dYVvj3P6VoJFQiKxDrkdDol90h6sPJNxxF/8tPpey3Nh6CFcHDZspX70J48WZQA2anzVEKEpxqv
yLsnBtiP+hviZwkTUnJ8Lt9FkoCffnthR0v1EH5cpOBldO6zcozrU2toK24XgITpWHvHNHdAPDQM
imzT2+kDIXAHFxADQqmPMHsbrpsXCD2K5TBzzE2bR16eRUbiQacfBVEG8aZLGEtqZr7iP9joT0e9
wSKNqu/eg1xlBNvONWwGBCvwrzicpVTx/IIBypHfFQZmgAEnvwZMNwizd8wb6RUfOLgZ/xalDzC4
puG/aToX9VUd2XBg9PauJ1h0C5hGA6Evp0+Lr/uGtOKMKAGY1duIbxgoBwZk+ufcetxQAEhZi/vX
vSxeP3P9H8Pcj0gL79YatUH8NmaVRuJ0sxUktovEBadUhIdVyWcNGvPJPdoCWLIofcOuaOclZOco
hVrC02Gpi/kwffV3txvmt9ILZFQpqoiDtFQLZV1WXm53tl4YQl3SkMmJSOsdTpBvalpVv6y9AjOF
xoL8M7y2HMa93zFVbzVkaBg0ZlSB5ALl++gXaT+gqv0gbA3r1iN3Cr2oxo9cU+Gv44ezG3jY1hyp
JqbajJ0kw7uI1ykp/P0ZSW20Ht0HlmJi2aE5n8PoHFyllZ1bKiclcbnO0PLhCFyotZIIN+mZWX+q
w4W7ALoEJUYkv2lYWCwjKpYyGZRly2MntEifzf1TzxqfIaI339pamjikLsMjdPw+MPtAMwziEB1F
vJE2LbXWe2n3ujQrEN5K/cDzcRhz+/aEPz/XjmhrbpzUGvp5P52IZnkRXH7yy3NE9POkQ8veThMD
FOMd3Lqss3g7dgFOh9J2E3oB7NYBa56Nj9C9R79RLit98gN5WiVKTuvVzUsM4q6JrrtvM6a2n0/6
2VxJpTOt0dHxUn13G8G7YPjE8KKyWoT/sXJvQ1I7awf6GUJPHyvyqcYpa/NBqzK51Yi45omo7Z5T
vwiBHcwj2ufHUJGUfEfDrOWa28mpJ+nxZAwoxLZebBKuhgn8rBo88h7WGoLMib7J3XR0aif1GICB
6+BFXxwPKt0Sx//kI12gx38ME3imtwTbpj7CJkO+zL6ebN3Oat1AIXzKJszTn/juwZJE5mAoRRsg
gDLfPtPm65Aa6Rvn6GAjCCjpUGbQWrtyXExm+pg/2MBWqceZNwm7DgVm5DCoLpHa3YEBBqrjZHD+
wPgloiyWjSAX5J7FM+ovV2wZ7YW49ypvSHqxpCjQ14dprU2JWlz+3TW5yY3yqW0KPpBywHbFudKI
VqwhIkLScciEDOn8yIQ0H9TmK8RrXCd46GkWtFDtvs2kRE+nKiwna6sOcF/x3eyuWhKCt0628pcU
CdK7wCFZZ+ZkLiJxZvqa16CWLu8HVRUxzm3pZ6m/8UNhBKUBMKKp6HBhR5/U+KKCoqWhXl7bz4q7
3QLaqEvHGSN1EsjJh8rr9MWqS8z90PUvD2rP/KahIwVHTHfjFVjwOZzKP7eexxfCxS81mHowJVK6
FEwtqDi4g9l219GqPBe7L+YxYT2hniRqVos7BHuJmXhabAhu7V5fOGbm5mp2PEQxe+KOWMQvPOlp
8jiJPBMMhOxdL/dvrAzPHC9JXIeCll6RgSxIjQ35KkvYM+XEmh7k+/AjpvIncmTh6J5jLc0tm/fW
7jPJ9bj655cuOzRd5dz+KmtWTVCqdm3ft0AX+qOe5UJ4fIYTT237ju5PEVw1tpnIwprMd4YgRWaK
pJ8/wbbkxzekkJIYPhJUhRUfMDBmfOk21Drcy4bRXI3drAlP5kaMac3Dkio5KReXxao5BzZI9eMd
dFx08TXb+Ml6dDaMnsp2v/wPD9f8FDIUqzR2u/uqPzU21zWWlsgYVUPumTFMb3DMXIfz3UpdEmk1
3CEGhsJAN9j9LIJWcMghVUexvnsla94HWDUCO3RqFn5R85+b8iwsc5lZNR/C7M9et+3SYStIqMDa
f0yzQr4JyI0/Jwxu/K9Qd6HlOhSj153K4LV5iNWcratUDdQ2xozI0yY3AgsxLXFbhq7IQPJd0AjX
rQvrw8+SwlCl/bMhFMWPfZqtjwUCXwr+yAgW16mQEFaQerWf57YhU/gcwPiBdWiKEpS/Jv2GP/oA
BYghKt7JIbNweS9+5BNZ5XG3s5CBsuIGWob2cEXtlVeVpjd7XDa/WRR05IOWJeLQWkAjqqBahQgt
2QeUjnI2H7AdQdqxJbZutT6B6qy0Z1IaIcZQks6Y5dAugRvhIPpEqQPB0jn63qAxZTQYn77DPCWV
03GoqHf18goVIUpL1zMfolliOZ0l2L+CoBuh7ScYIEiXD8hGAtN5Rrm35CqXvITpqLFSYsaNYwhu
ygq5GNcHoJ7z4tI5sh3NAfA2rvpBIdJqmauIrwcLFImGkahwaAy8E093UahcYDgLVoSaCH97+bPl
LFDPzFr4gmSWbvZtl2htYod3oysitwyFFmlZpFqH8ZTHVMwaUCPdQliEIkam3EsSgcma2pKHh310
d+JP1FvnMuXqA64LjE7YADA32l1Tw1f0uDvP6XYjYWbmSJrIppJmV0eRxVKXlA95mgBA4Mq+o9Qx
wjSiobZXas3k+u1FfA1KVkQhu5kRT/honQ3uWoNBFzjYNG/Li9xd7MqVf+qbL+z1tgXXKdacZ0K3
E68YBxV08waStSQFTeHx7A6mLMyt46l87m8PIzfxwgkVAau2vfvZtfr5J48rsgROnMxfMvfgEmoo
zcUXcwjcIzIA+xjyqGzjPbZNCxslE8KIfiDC6kyRHOifpoBZSx+Ar7oQvCjZpqVfqn7mYk/Q7R7j
Tzhdj2KQylikJM5mfWEcwgQ6IZpwedYsEV263wXD0CZXGoyMuI3dLvkqKi+qZoOhPJtRNyk2LMgw
mtWCQ1Q0NA3wEaNaotPOAqTZpH6lMKWEZbPTUpoR+MkV6RFiCGr+wgPbW5JvRaroYP3D28wnMGan
0TboncOpcPC5/onS+xlw8FULCBppQOV283dUE00WGzbpM7BJWNc5SdDv4sGRo3hE3bChHQmV6O+k
h18HbxJjrk9z6jeWDx1yoEAOtZQrvXuXRfzsIjHCf4KGtXHEXPKL1vJjXI9ZvEsZsJe7DWR09g0r
1q042mRoDXqTTY8fqL0YZsjDWEwh+CS7ar9kzwrYBRfMqnSyhVGkBJ0jctGgg9XoJgQ9xwQXeHpT
liihwBNjYExVY1HxSWOpk5RYT2vh+riMlcgGx2Se5ic814pwE4dLP1GIZLBM1WPKIEiXu2BAQcm7
LCC9rtKds3Q9GZ7Kdvc61SR/86hjjGiTuw0lvHOYWCUocgjmGeGnsincdlzlDFFBYJlcIR6Erb64
IWBKq20NNYyKpBFAQkjITOQwGOWsZB8YKDCI/f7mhmQg/w1o1ivUL6wIY2F7uYkxQP/9Qm+8u+mY
Y+dwoxdmMeZRJBz/Gy62bpQBKAvx6T9bWMr4n+6it7TpYX12aTjNfv6+CQljvYRvDVubvk68PWHK
U8pBUJrxIF5SlrfGnsY20NBQEomVopkDVTptWnSgxF+OFJ2EePitjb1Njp88mv7vNowiIXaIkl9I
uhf7hot43fGpYn8N9RBsXZ2wIaHm2xIwfzeStgbn5wlDx+6WMU6eabUvbul8kGNyaC+r3zMiFW1D
AafNLOGKn2309WcUFcDVgkKGOp+4446vn7qDKGKSVhNrLh1NZHQ3+m5GG03tQE0GLerjAT0bRUc+
wgGoyd/jdxBXmgXcg++/vE+Tmejn9umD1KdcDJAkfNVoVQot5aQrK0HAKR0W6fI0ksyKTR3O/GUR
8qIC61a9tA1LZjR3gSDs/ULS/Y5V4wQphnC+hnT8XLR4NlfLUoNZbj9n1I5tafmeMyIKiaoE13NM
+B5/6NLmDrNs6jEi+D+7ocnjTVFsB3gUfwxUHmdV9BxT9DFV2j3XoqfWenllJK+WAS7Hdq6ig3iv
Vx0lV4p1hxhEbm5u5klIfk5EfPedpZnj0BMCtpBryaN0m6OlkWw5XJHtXKDyRN5GTQPaG6/+R67D
52FLVqpNlYLhAiR0EWw7EeyseLqCLMX6L3bGT3OvE1i7y17lsedV6hkTYoG775YlVxJ2LRR5gRie
3rzLgCEvalD+QsCUL5cRGl0QxTtFAYxMnESA4pksAPs3pLCVbrlgHb8Th7nRrXIHBCV1xHriKkRj
Mx+RAigl7bHAyptkcWXAYiD9WUjHv14gwSgOKWzZkyfKWF1ygR4sqKCWp/0EM45vFlYcYexEgvpe
lxaPs+TjjXQAI2bjrQ9tm7QUGt81esuOPdXnQgY4b4pmdwRVc8lCktl4ESOiilwsUy2EEF0+o+lb
Viwuu4egdf3TXiOc46FViQyuduQQxnv4hb73/PuzdpuzLrE9VIngyhC+JFJYU1Bjg/wXobEorGhh
bQzjZVaHn/6sp26YRdZx1r72/UlcXSrPHM05Xs9RDgkzy8qfjlC3DCupmIysQ80MnIRCsjzUXHnE
7L/ausUMwBULAUN5SdYKYXKOcQhmcYmoXEqC85CNdaXQ3fcDl5Yy4Jh8ZGGwrZUWY/K2FoZnlH+d
fyoy2uJ0wzXJZi9WVogRVxsn+SraFoxCLtYr29w+vu2CdhA2088P6S9wgrms6lMLQ8J8GZ6qycfu
0OnV59QeyhggUidYL95eAJ5Efmjlu0EabYetWFtBLlVP4H8TQ5r6nT1YklMNYrf1T/Dx1BIzHpA2
uH0CxULKbUlEsFKc2PB7HhCIXrYOQHw+TKRn+Sqw0ZcuC+dVdHNH/HpB6uENZXsNIPPKp+a1vR4j
DdRtR84cjY6ynLURkYpPKqYKGITikBvRIFd32ZXjsQ7yht3OS25Jx9YUkydV8G9aeTaBGPe3M4Jo
lp7ZL6TGbxWD3lMYGZJy4fqgR54I4CYJi5tKPNaza1AYhogTwgGQLiez1GJuhq9l4utl4/30vGuY
bh7dLlgOjDJctyDudXfVfptqaDZCLi1D89mBqdCAd72InFaWSSF0WjBJQQQHdG2QzVwZovVXjw80
ui8J4ElG0/RPUmGK2Xbq+iWiMFXhAujDs8uRKfJzp72D2jE7EhXN2tbLmW2mmf29n73A/aQ63q6g
IjYccqXg6rhjwHvmoRs8VkKIcffIftNRbJUWo7Pvq8VB7TMfgi7vaa0X84QDXffBjupQ9ZUFGDhZ
MvOf8AJCQkRkvTP1xUuoeEB4li2tz3ro6sYnu+r16MY0+aOh/aajtXyAGL6VqtQKamoTsB/3cftb
5ws1Ig6pv/AgAekDf45JbuGDrK5vmEQM+yBTAiD8hnxckjQzVuNrenBiR4sw0VGw+Nk36C2TDNet
cLeZcAsPrj8p4xtj+7pTQIG/O2tpAEn8pCnHpEpWChZp4LibeCAmZm2JZPKeann+3nKRHj3KnTaU
rIrRNIlNOq4gxWg2vGLiRo8n2SjmsvbqANbrfjYGkfl0WRECs7ORhodDUsyJ2XmSYh49r7hvfnIn
FZeLX/qmaI+UHUkN68AZd0xENF7fQsyeqen9U7af8hUOqB3ZcjDsDJMQwTnC3nexEaDYu4Uh04Ru
pcQmfgwCmzyie2c9snZmMWHcQfYC8FnuUsN8fThGlBTr/X41x+aNEqpYJpmy3HjT6xfoRqPjxwlb
nJFAKkFhFO5F+lVc6kj8d2TLfG0Qtk+CdTSv9K7WwGyk8F/eFPbQBKeIEv7yVzb4qe222/2X78cc
HxUb8Aquz41DViQqMX7AZJHurG7WnZRUBJDS+PfRzsgbesMnm9OKnZilkWq5dMzRzdmpIv4vgcM+
NYPeMUbNx1d26WWRXBVdTvjv8ZhM6S/QmvhZ7ygiGKBe6k8fTNwGR1qwf6232Llo+0incYzAKNsE
9F+zMXvkIq+xS93BxbqEXIVsJcn0N//GmFGs/OxXvQ7h9CFeyCWIkB0eS7mk3+k6Ibkd8UaLHA+6
CmaBTnulyywWROkn2z0w0+Sh6oOgXIEQOYKfTrsX9UYLyDJnPuXBydWcWV/6ES0+0TiMawYjqZ44
5W0yau4weTGick1OYiwuzD+qQrFefHNVLLX9LV3ql2bw++bQgfgvU+BaxbbK8xK8DRcuoT3sg+Im
G2GRT/wPhQvzlf7g0vUSZKs00uUH6v3ojxXVPSt5zcR1XRwzGFs1NFoZBfdFs5neXEEXGMrqCc2n
54mpp8wpYLAM9IKtCNTRULmZjezuN7pIxhSAufXMawR0yxb2iskSxN5kf4YwDKrkLZSZEH0NaU53
7bvxFtTJoCufFljEjBRspRECSqOPzhM2nx/Rtry8pTJluj9SNXFZXtyLZVvIkIkcHom/QbcHFUbY
61vgmzVNQbU/1/S/6s0f0/afDFAIzYGg4YU2L4VGK05Y8T+I4yiOqZiT/XbY0F22usOCG+FzvZny
5oQ1ue4sGi9h8vF8pcif+GiAivmOGm278lIMk/QPtawuu0z/jIelkRWomcuzgz+/wN9H3r1K0krI
AEzawyXHrVSyE7GxS9S7BqigzUltAdK+1kr7sduXaEoCN+eigO44WdFloJbp9hRxkeT4tVR8vbEm
lnBR3gY5tKY67p6xBEgR7wcBq6xnONykydIaDWVU61iBXyn4oJS5F21LclpzOGmlqQoZ7o/j0XVj
vW5gp3m27NqUWa7xOrWKjAty1/EdQEc2ubeW9zgbUVYaXpWala9oikLKtu1Xf5UtR9l7XU6zO3k5
s5R5Xin92a0QzmjblzSDecD5HKhnyHUWZuwIkeZc1GLUOi6MpTKFELDsMFx9NaYGhd08wzNE7ciO
mG7E1kGYkAPxQbRIqBqDuLxoldn8n9H+HinYLGGktucU6bkmlOCzKgGXkV6KYtic11q+eCk2QDTD
dK1Jn3JD4PqfS0GLMQI7VWc2uqYO7y2WUUBu5mka8yW6RFJx2Tt9sx5D61bPbkrmsqq5fnZx8Lte
oA3/5JnCAzdtOPZyC0kjGSYzTl8QZpInWfnWPoS/groRzz651TSoOHe+uYuPJuYsPsSSbPYge5sT
yssZ+SXuWt6RBvz7JPXUjqVusZJgs7DJ2othJucCNkfE58oSm7sn+eXfcjzdAECqaZpl6gnrDZ0v
LNAtLd1XdEEuJU+MqG+u5hFMiSaZkiluXtAfUxY09BPiknrCysoE2hMDMD8rI85SS+jznjl2sZWS
aqikRMuouTa3GDiqrCfYCdg8xU8MgrG+4Xk2u1aJ78lG/Sjce8c992yfBdvWEZ2yhtr7m5q8akjh
FEfiqxX2Jjf/6z/rY6E6G5Qa7pspj6HP/7HbpoN89234rPh+ZCnw0a+H8Kcm2Xb3tnce/WljqymY
5j0aeKptPj06GpC42+41SntIVwggu2CdIyQmhXVU5FZSc6ygAkQgFEqOmwlXyyJiutZQkS4GmUuS
d92HFz/4h15WgskXFf+qdDqe834hWTKdusaj9TRjg4J8SV00xcEKRoNk1OdQiyXcBTQdMwnKac9k
yqz3aDu5+EMBCAOFhpaCeL90dAWvSkzPVINo+4X/JCWBhrWJYGBUIbS/444WlaUUMZI7wLXiWROR
OQaFNsNxxpN+G9hHU8fmUqTbR2HUmkJ3KMeNEn1hwAsgpZX49ZKr4VEXSLIskYBmWs0iiFYaHgBo
69XT2+156yxJSnPapgssoH8JiYve6B0lvLzC+VqRmzihQIRCD/XqPdAFu7F7Y5HffvKvfjZafpB3
pEmdGEHL+SvdPINLyeEIyhud+p40AZxWYuG7ORO7S1Kp3rPr6tx9g04bxtwT3qSoTk1W/xRrg6TK
84nkWnodZl8hM2DPgavePmeG5ysnrQ5fw8V9H0YXAr/Hkuoxhue739iXfS05+Ct76WEI0PWQ2kR+
nUqRi6u5i/43w7tKlP4pOIvzqWah29wGkGfYc3r90Ds3rYEcOYX/1tqIxIwbsoi3ge3wIVJ0cjML
a97Jgn6711VWN/g26iu2wCRde1QIURMCB+/CbIsNW0su9t/XMYEWvxo85gvd75YmcUthZ62MvJbm
3h7P8s3eAFKN1RQTYcjgyaefzom9bipRDOk5l4LaxjnK0ZtSEJgznR95gSICesn0HTMv5ls30PCV
P4MEYmx+HY2tqbYA3j6tlB8hjkAF/PBub8dIyUkxQgTk/0TJ3mxfPhDF58MiWc0Ot0YjcHZP6ZzW
4txjJY3Ws2aDbMAvbSW1YzI1vbMMjMJ+Bs6uuOHEgcMy85dffkpfHotaDT56s6CQHE2z7xwyGdlT
51Al+iru+gHkZDGwQ6pJTyd+N5WkvFK/kcHiiltMgswX6pnXpaGq6b87XzsLHxGHUOjMW9OaAim1
RrQfuZ6wWbqC+sjDa4CTekev5+8/T793ddPBUoogj0KXZxWx7hPcHI/M/PhQOzBFUho8KGCpn8t/
RV5+qxJFr6w93jHNV4M6sYICmL2bzwC16CTqVRjVm86JRoDWngTE5QMIlzYhzOEb+q1Dy/zKzfGk
IMwGtj/erN90ORTliVlWaQiajQWiFd4R8NgBkAHB9s+JWJ5N4tFogEu5ZrBmpYFTeL2omGkHap8U
j9nSqjyYxaBOQr1WLAuR5f4dUr2HwcTy64a9X1rpAwZMzewiz0hlpEKs3pspcbN/UsIR89k4R6if
Ae5GWGLulHpyKGZNn85ADvA6cBwjz4GOTHPMdi1TMlF/wVtdOdCu0pBffTATNQmj8HKpZXMaIFhi
8T3EJu42Z9ClYWIAcR58p2gpgbCMPOgdZnvVVXEmubag1r7eatvUQnvMKEhZ7n9r0empM4ivF7gW
SwUkAggil85Y493FWqIIKVJrohsvv/udHB5/6AY6H39sxDe5tbWur8XhzF83Vkl7FYYJGCKI1Lhs
LyAG7koOuHGKxDK5I9+wTVL5R3TeHdr7QgfAw7Gvvs9afu0h+a8rbNT23Yqty7Y1rwzgOw2y9y5H
hDbaJSFWRHn4KGDj66r7OEeDXp4jtBjIUKme7QbuM2YryLHZHCd7QRKPpQLf2EmKkczlw/NEfHez
yqGTO+XyU6sNP3Xqhq99SNdPooxiUZXbg9on3EWYqslAO6Yl2xu60PvhDqrkaGkMoTu5y28Dkfpk
adgPNBwrFD4n/4K1CyVIimGPhJEbV83+nJGrDi6Exnn+/i5qe+QZK86WSVSMdepcsbHA1BC3Jp1j
c+LOHMFvY7KfHLI5ukpexMgTc9156Kj4AmZ/kvd+9hmQa5p1pVbkbG3lKRrb6BPK2F7t85sa8Xcq
ZD9Ek9cg1sYMWKue991Uyun5w6CGA8vrYZS6rC/hikPT5d+0D00xfd3RjF2zkAvhDOwYYHHzdZV9
eULMJvgEj72N/HQ6zQ8c8L5l9DpDAC9h5sH2+pusIoE+8afd2S+pproC5L2BbW7W6h91TMD4Lvsy
r8GFJg/I3YMrNazUX4hrfoC357muAKj6ju/lHTybsSUvuinvh5qjPSsPHm4CWg/Tx84d2d6+MS+A
U66KPOt9jQU0YwST1/DzUMVIoBokiAWGZs+Gkm0nrW8oPlucFhuU2Vkf2tjACWiQ35AflyzA4buA
aYjnxmpJchxshiqrPjj0Y6P2tulVvtq06I1Cd00GP5E086qydUKnD9DZ6hhKpmi5ANST6GcxTNO0
yUVAbrXLALobq1YBZEf/bQbKmH7dzwE7smmMoIqbEn1NeWc+QjFyf2EfLbXeHdkRACFYeReZw/IB
Yc/dqIKshMj+uXp+onW3qjzLgJ7kM8h10GlY+x/d3J8bA6+mZiDg0rGzSR43Vhcc5CjjuLQspx1c
7XaCxyvLQPgzEsO4jYz3f1398xZkpqX6zM/W8QZ8WEfpXPF6YW76f2IIOJaRyX5BcCgyjFxlXhri
FUY29DWAn6TieNjSv/kfAQSm4ccv54evIe7uFVuXEWkTinw3P1pgUs1goGlYneLu1LxK7ISdrx9i
cWZ9yK1lCW5R6LBoMssiac0itF6hgGu0TlowUMVXmAAAbsr3lUbdrBT1X9MNZozvq09t5DR0mDIa
bXBPjmBcEPY75xbvS7WBF9ox3x9rj76ved9iJq8vAGq8gZR+DsqteO6NDiQarecP64Jy0YP8uqdC
6faMr4Zs91NjUP/ze5CC7ZfZ5WC0v83Z6RTCnT5CyUOXm+1dZSVYAyjOkHgb4qpNA8mCkAYKU6a4
OKFpZ/uJdhOLkm1lLe3nu2nZdW/9UkLDU7T4FqRRrTxADtIIkd4puOBAlN7p947nQWVjtjMi++P7
3LkByGnLnF5fqjJhe3TqT/rn8e4q2uuyURRVLsrUjP+oHStd5XNUmg2zYZFWUFMTh2tzGM4WJ8pU
tl+vG30bnhGUmZ5Dcoddp80t5WqgodKBILmDCALHWSKk/EtaKrI5b42FxwZ2epTy67d5I4zdlxVu
M8vDw1T5nupZ+KGACx9yqzhdjZcb6ln90uV/C82Nw9dvJHRfRhUBKpeaJSIVE7U/cuuKtK1Qqx3K
toXci6tkEEM0+W0yVaf/dXScSuw0ABIPfU7zrrjxWZosJqQXAiZ2BswztjGtxRwmg3wZeF027jes
+yccZGy5jCxq4Bv6rAxyJ0fXv47a4P+DByQAf1vzmX1sxSqSCoZbVGtWhNUTo0lRaeBE17iyrEbf
FwX1R3adSQmnSrsIodTujZurJOLKtzMVnDHuy25rcAeAJZgNspi2DVkjFA15ksKd1xux2WG6m+0y
rxtev1GWSKDDaoqDouHMqDULX5oCo2JPG9eW0HrLNh6V+zYgss+TM0TiKq/me1fAXrL56yKG4MqE
QuF4ib2a2llgysE8vu7a0e4eY9OmWFqg3jYgBOWwCZYgiYanSiqHN9os0YQj5g/FD60N6Vokz6y9
5ljKfjb0ACMWcCkwKmGkH4NS1D4o0OPKpsK+p0InRahTNfYMy0YczEv6VwKXyxdL9gQ0FOchXxPe
4GYhI1ndD+QoWinCzH8/DmZOIsbvIe6lO7KIArKwT1nSKa02KYIPMj5dw73NlBT5EZBe4zY1dkBk
17eOAriBy+6hQ+JRjmnRizP5H3Nrg6G3H6p0jkEGJBdqe+7kOshjy00yrgEXb/2KKeAp+a7MkXv8
svXIk4DsJxir0SShb2kTWhWJ76VKYmOmXtTJa/2UIjwER6lqfCmVFPXgNdHe1fJS9EpNSiPYHr82
ubsVdKFuTnJGsuc0LP0CG3dKrGfd0Azqjrnq91/EZFE1yq2riaeiIAqWlo4reNC+VpRyH12qmLdu
j4mmvEat9LibVXPTgjx/yOy9oat8v5zv2TXiVjNSlNfTTyA174MxEzj9SOljighavciVOTj/PFU6
uuZBOCLyGk7c+bFVbqwdjQ0mklObwkO1TrU9HdRhLr72mWJbXpt1H+QV5K8V0OqSSsmIWlkv/acx
gu2bCaarDsBmkn1RtGsqdqzZSfMKq1DjHj8MlS3LAIiVZcH2cUipQ96vzp1/302Sct+SjXtBWYfU
zKF/15QMXPBMpEz5jVcbjSX99+9whIjJ2o36q8VDhp4g7oe4LqhYoCpaiYy4TPgJmdOr2fzKOUbd
BQyzXJOPID3UNPURNz3E4GV7s9+nopZ1bUZLNb6rSfhkNekUEXG7VRDiLIasOlSUMjNChCgKffuj
bR+QH8NszSfeWIN+sL2MTPbH23e6ULeX+CokCIz01nPacWk4SqaDiybJi/e9zJVQdQ6iNfRlXrCk
DotusDc/CM3GrSaud+uMIsFSycTlzWOI9fETTfvCT8e6TaL8Tw9EllQYoMT+vQYXMYsDvjxqvXLv
9jvRur2bADCC1HeP6wtYDX9jby+ADQ/g/qFOfFXL0BAo/dhnI8NNI5TP3g9XDgJADipAUst3hxUu
6jP3nT//3qKGJEI8IlWdjLWJV1KCNHfYFYJwJeEtTwusRHoeucxmjaTcqnUwEchnRtW3Y3tLHNV4
gRX7AasegY7aWkCcY27ptCXmrnAZ+5mgquVUwPLvKD0YED+L0qlYqnS4wT/2j4XY2b5VXBb/0V6M
UB/Q8BHYgqwcB0gLs2EHhNQwhdmKcLbNRZuCPSzQ82OUAi1y3un8Rtrojq/QYGChN4YPqZsCkOB4
58ooCEaRqGMAszdB0jR3ZloZck1id1qtkZ0+XGK5gt6klf/kG+GaeYggzlqEsUpR3CEOWLLS6lyB
uRlJVYLX4uzle5Ja+qWy4+CoYROiLWirDeiQAbYQuI4+NQg/7xSl5aYnmanUXwUCZNIw/gejRCZb
ytwsRpHtbmrq0zNgs3zZxPzeacKL4rS7FL9gx3PWK1Xdgmt1U9KkmxsbfFIHXUAJpNd4vM408zv+
BcqJ29Sc/7qxizAi6DT9nKEz/4+p9XY+iX8wapB50tberpmqEG+3vZ9XBAguvgO+UJ061y7q+RRV
vpIK8RuFU4j7cc7XTn/MrV6f9AekAVkd9MU9LZDFwRL7m0tdpdB2faT/5/ntX6bj2b5ezE4FIiUM
iPSH/Ya5B3/Ff6CzM4VFyiG5JgLN+0Js3JK9/rin2IQ82s8qC3aGtPEgp641jWILrsP2T5SkE5FB
SZI04SkekXG1pi93mx5r+x7P3/4yrTsCrpFhj22upyFE7gC3Hmz+vFVUdIdKAHn9qWAm6HhTsXiK
74fM3C7IRgBQeihYE4a90PvGYtcEhLWhNpAvDaEY4DCWoHiorCFAp7DIikP64ASKL9FY4C+KAuUk
Sa3uMQMa20F98StgmQgoCqcXA1b5WmMbzxGThuxW8BobsvxN2IL9rzVGutGu/zgDyuR0cEsfqOb8
xsDqPap7jdslRBSShqIYUMcpjH8VkdvTEoDQW7NRb+ZLLxDMwmG+sgmqPfTs/nABtgaI1fIoSs6W
nS6esixwqdOCfjLJ+ox6rW9S5lCiGD5hb8TvzY1D4fJAY4D+eTWew8IQhina2nREUpKZw9zPElH4
i1BmOgP69rFQDgy05yOo6sQlGoGAhNddU0K48qXPQrgGOJUZmoRt160EerFo8opeWsiqRte9xu+z
mEWhXC7pQGbZ/8QW7ahDvhFXAqpB50a51FvBjfPRlNtv6C+H0Coc3o50rAvV26d62YsfrNYdBqRq
2nTlSjle+PM9PQSOGdTkquRS7vMhX3IqjTGQPYACxiksXnFw9xT2Xw18cj+oBvdvxWueiSJbK3xS
BWmLdoaISKueXjq7QY/H7m7gaccKJUhQZ519eA1WRvVjbwp9WiXYm0Mlb0jHGYeS7yCNIieK3m7J
IIs4dnm4w7v48tSd+08+NQ4GFDaJ2xXw+ktq/A9jVAgS6gCiIy1F+634pRkxW6Nu8XBAjIrZPvls
GFh1fQ2mRCeUHuZyKCUIoX02g9C5W+qIDr4afWtONeNnAPbMtpc+YhzV0yUfqLP/L3VgU8VXdN14
D5NWMhff+gtmRf19gtMQjDYaGyHNMropdE7YTehWZH7O3hzilOXpEowx82dADb1CWHlBGNbpArWZ
tn+yLymOhP73bOp27c6rVi6uGx1voGdHA+N1+BhpkPSvA30qf/WGFhX53cQThlJNlbzLBL8Gscej
+TCE/OZzmylL4CBnUT1YDSw4G0lF1XyZ6xFY8PmdEGWEGlk5LTi5sv15OiYkJwZP12iJUev+TR9x
KyocXZu9TEFr47NUI0dc7YmdZc7MlOI8XuIYi4cgefbc3XJis9cUJoCJQOT8By72BUH5U+weaZCN
vqrAJaw8vmB8yfR8S3pogDxsYSKzGGxUza7+IhI0PgnN3jzk2+Y1CUp26Rm8hBfSabJJRbe2Ovmu
YKfYPk86W7piaVAa7W0MvJVW/MLAjs8/X6jU6n8ilsAUlx6LGJNHmMPwyvG7e2dNZ6hB5dv1LJmz
Mi8uo/jxVE3ybo+B4QwCaFJHo8BFJPQVbRcegHlXLrFbPEFf02oCAeN/WiSzSSuIJN1EkPdqXzKE
AwtAJyh/w/FpZc4S5FnL2rJv3bGfVjEhXd5f7fHjOrZ2O7VcBaMgtZGdN4wqXbPcEIkwqq1zMGHF
kZAuYpDW2IkRKIl3UIwDCuy9GIA6nvUtse/ZkeWwG4ofWLiZVlYVj/Xj/ekx4azqFz/YR6kQ5hyr
83ios01/jCkzkjNMZEuSnHjXhCRRxVBuFNVFw3xWwZTfA6/hntR3JNYDyv/WwaCJathd0mA60t1G
z4IROmDvXRLmagJSiK6w2tynRaHfmrl0KQGSLoh9zAC01++1Itlut9L68AyxXUb2ENOMAh8I9r0D
Izexxn1A+SM2UEP3Yeq0rQ2F7zJnQyp7oaGsT/LowxDiCejgvDkc2cK+sKG9CN9IEkdrZ5h6ABBa
Ftq4TiB5a0Tvctvv8UsW8+b23cBC9Pcp7uys82ef6ngvz1UDVMsshYGg2Ro+kisKHFqkTklAk7VE
CrrEN9rw2ib6jLI5fiRxFOqRrFlhNtpjipqGgyi0ocwBsV5zjtt9S0sHAQ0mSlBrRg0GoGjnCut+
Fy8eYtbmdSj5aXtfP4RtGHxmp8Kf6iIHkfd4JQ3dAoL2Xsd8bR0DINDez5AbhP0f9/M/kKW9NZf0
cpUvMFoO5lH2pwf4o4IuG1cZNL+IbTeEw6r37L4sQii29L0/nUIlZUJkVgz+Z9ZbedMF+pMKSHR2
wysGpyF7dbactsUgPhIQp5mPNxBDFWBxyQrTJII9QIQDDU4F37AbHw4KQPvy2pUtaC7PmnFOza/e
a4t0uH1aFelazHg84tPiGpNfIOgNpa0kDPXdo8MTRnWdQeRm/d9GrD+pCZn0e4795+sBPX/J7pOn
3ySW++LC5ZqZg4c+efYyB1TUPkJD4L7Y6TDWPIUenz+Q1ZV0qsv3u28v/BOXk5dmYHcggvZHD5x9
T2L1LDdHXdLbj4LI/cBl+fAQupqBVGEWSRif2hqDzsHEvQLgu91mfHdDPy1jV2YJEIRhEN5XqYtL
fRdw0KyWxJnFwO4e+HIJQezufhA4t4xZLtzIJfeXQCEyuA1D4Nezju39rOGrwJ0pVrO2CEcQaUc8
ZqtknPNMqxx8FbteO8QQGsCVSsNHBXebg3IxeJyB+THbWBXELvqVRuJf1QO9VQ80DCV3wY7oERZS
T17sr39yQoUmx3WPHq3Nxoackyk7pZ70mQsHMCDIB0w9vWYdmn4CwMky2Yp8G6Rc7Mi2crzzRrai
ZqJZDUPSGGkIY2M17TNFnCrXttYKsN/grFqYHXFqI6xlPROmcxUNP8f/8JipCH58Dhubtl/RSpMd
V+YUlQVn/a8ZCfrqiP4WmLxtjbq9MW2S4YnJh0z7lCdL4c7EKKMS6W7TIbCQF7RhMj8nxY2y9NPC
LMeSZ88FhO1nk27DH24SBzPVlsQr+JlqeAOH1XTgxxMQSNTUhNPBDFMRz7hZxIVvXWwmgyzY9dzs
OdZYvI/BUWhqIaVw0bTODzM+BybkMu8YpgjgsR8EgmzW/933o3Kc0tVTNbix3a80Oi3n3TghVe9Q
+qki81qW/+Ibi0s/+m4oRclcVSo0jfFGk6KN8T/m2W5iVIuj71kO6A1rmsJXoGwGPYU4+eoHkEdz
okKNhZtbEEi+9s7AdMTCHoI2HpkKiqoc190ArK2uo7ACgLWKbuapDVPDbwJSDBknNxRMxYsBlIAD
Zdc1BRNYzoXEctgKiogisBbmT831B3g4bt+jhjFw8a0tlRstwa+WLkCGq7FouVT75tQShDmD1anG
20MSiPx1K7U7kMpRYzcVR0WGAi44hMJUJQwjbnNU7V1rU876RLhqL6ZVDcndF6WHs0H447C/WQnN
VnZpehTGmUp72MmrlP26F/Ku4+M4HlQOtB32b4+sAO3hrpsrG8QHyzXpLqlN60snmJui4qu3p0uX
ab4qx9Dri19OKV20QMhmQ+O8/U6Odtse8J2WmhET1X8iAbhPPjVWOnNz797MrkqqzO24LlLSl3v4
DZi789jlcohAcwlWQkdNJNCIGXZUr7xxnabESHfT2HZDs9siSBfl0D9Fv5dDtH8yg0TuCKcnOisU
h28VHRg+9K8gXn1nitmaYI2rM5DSvqy+miqhrOV0DfWUtpNxfrkjTw/QYjJ1lLJ/9sm/BUWkyidO
Wtx9dj2rYQYr6qrTQISqXpPtxMgoX+9Yk5zTsB0uWnz5oN45TSlhjLkTjKj3mzb70cRyZrIsco+o
OY4oj8pnT1rxD9lZkhpa+btEi/6s3CEAEu8TQ+GRafDwj039E/rAk0qCKXeNGEYgZYfcBczf9jJ5
PQo1O3bxfedplNMvmdY2Sdj5IYMG81CLA8LEyzgpbrRlq0bWzyLVAIBtbAIUdjawURbu46LjbT4Y
n53Hv5RdFXIjz2GfeH7Gig7s3tOFt+0IAzv4Jdjp2ANzqRmoKLcJzGYHcPXX6v6xbRXSFx4w71Qg
+ZPp3p7/LDEOnvAAjuJQWE9olpW5+2eRjuRFMW/vWKMjpPhdqDiww/p0fofKnZ4kNZk6SBrVz1DP
wiukz7XEtC4op8Z/gaQRYPG0DjoTehoLUAkSu0kv8NVXXi1MkDwMhfJshWeeJoDYYlB/xk5zP4Nk
KXr4lN3s3nVLI4fy8iO2qfK1htrW1i68NRkNUPRmTWu9+Ptkdm7X3eyw75WQ3RImXYIAporz4nwt
y4ILeWalZuk+vHwRnAP36VNhh6/aIfWEl82H1LXZ0IWmg2S89MI9lCu5PdV5vjXITcMhlm/ODR8R
MlU8uhjl4QKIeQkhs3tkuiOn1SXdk3XQaCucB1vUMFCKv6USssG2PPxSb0sInWzS/nCvnBweZ3o6
s7qys/JSg770coxGFw3qxXXRX7njrQqOVMGIzqN/ERhAQXGh0yTlCm/lpnDP0ydtV+Oen/Rce0Kp
lwGc7cyPVnPpY0000xAd2xFkmnafdok85Rc3/pZGMdqgvRqxUhzGIvuLtmQk1bS++HY7nJcVwwoq
tKIfQLdkJRNVMTf7vF0ROQKkAhfXqeecmxLzCnyhtMxKwA4Gnt/yWoNSjTNxIWKPQJR5GLzpXAjF
AGrOpLM/Ni+FVcy/djlDKHnitOwKkFuYWRR5GXEjAI7BQ1OfN+xjvgQSF3DatSrqIQE0UoVXnHgU
trJr9exjDqot6KCjRXBnT0KEQXI0n82cOgck7375GCvT2GozQyQqFzkhfzO6yGFg/MDC+iaaZwce
3unjiESY+jMzRSIbkWGfZI/8To+hVj4ShOuMAPyJ/rGX66ZSU2L0sKjhFMK1Z9WQ2aN7XMatR0mk
h9pPbSrvHtJPn32O/Ni4jHg9gcogxW5ksKMFhm+yX6zopHrMx5fAMBjHJRUulP4uyJlj7cHT4z0R
o8eYJyKNY1xHAPhXfGGgjByRKEuAjkNCDaVRxUESv2kcblmput5MdyKuyctc2vi7g934gsWUz0Av
ImRsP/tVzfvVIoKH0s/WHfuYX8xFpcnvqrBd+m/Vb52kxvsIANvvkXddq8eDUShT3WNpaIm1vwVj
wTwxWtDR9POhtyIHy6Z3Wnbmg1ByiRW4N00QWZ1/qxS0g6hnIQZVH6OpLXf/YgEnSI6y4Z/xMcUo
i/9uKCxC+wE7WsHuHjPBMVd38orudN9vxfRhN8By564cLTBeXfUm2G15BrgKyz2AkKeyeMkP7VJl
uyJkf6fGgAN8K6jZVzWMjqDw5WJqFff8Mt2ipqsApRbESdftYN8hClBgMpX5MyQIi8dGsKpyq3UU
IUXKrkirmIXImcSrbdBOQinbx/g+JACf+8XBncwaHeCe6JO8w8dNOWPciowzLET63SekWky/1SMg
dSe+O46hKRI+tvI18mgUUuNVi6wRBFz+hnS1SYycVI0KT3v+xqDaO6JoAQrSoiRI6j+GzzslHnk2
B3pnfJ8hUQx+fTK14VEBEuj3zXf+oTJ4LWFzCqem1MoFJ8qQG5m7JXdCAdwOFQPghglXGBQchFaJ
vE667dvth5Pe+ntfPYGzGF70baiVcLByskKTHaGFuuVbo3ER9X107jBUykXZoSJ6ZqRwUWxOfKIj
yQ5fHRzk48KIAypZyYlxnXRhH7+BZwEsjbNWl48/zvmXWsvwXdbQiZL+K21HAumYxqqwL3mJFvcS
FxvxR4ejoXN+3Wno1zohoK5ACr7ee8qafyoQYjLMZF1nK1JGpVZwi7R0wDuswum/OqjBuohvB5W+
72pdT3CJbbxVf9vZyMA9GmHoktGDlOIiDf7K7HklKelUnQDJEMrSixRnbQL4eCUoGwwmtKYJ5Wwb
rrWamyPwAQ9mbgejyopJARFvwMX13Wv9Y7izzPrFO9gOp5CLZUISAK2ZX9C73qird7ZipVFzcyqs
rlEnJoYsrrnyvqqsApkG4nyG4VrEtFk2vMZJblmJKOjsYlvfehbJXUGAM6SlBSRXrnTfpJXEE4sk
OFH9bNlHz0Pw/Q8BhPC8PuqIU/8dyVlEnszGFWotPxztSSlkLjYaF+JGxVKXp/sy5NG1XyGWdyWg
Hj6aSYZZpXcaMdDYipsSqy4SiiRuhDG0r94wfJz8mNis56GVE6rMMH6zvCF37eo6Jr1TQ9X9eS3f
74U0W+M1tvnwDgdTklb4IwmdD4n8kLcKt+dEfeREBjlXVegRPuUyaf6+4UxyOKGagYRdLzLMHQ+y
pYJrW54QbIjU2iQLeNFzwErb/nfg3Oiau6P5LEgYavOA1jof5xVRHr0n4AimEFEcmb+/RKfoieWJ
/okKKyQKmgShCT1wnUOa0byimHB9PbeMfybWvskmHyqy8owYGnoWjm7jCmTCxbjY+EducitFZ4gz
Iq+EkkzK3YgLNBFZO3VVZ5L4a/Oh1N0UPOL14IxjR4xcNRVwgHpYylp8TFScH80wiyjxJTFV2Kd7
aE8u9xjDWbbuOGsrftqgMX8v12Cw1vbPpbFLtX4cIJLSxSCPpkBArNzbd+IiVsFjFxEAP5Y7WV3y
nlHCPJDygdGZ+SscYiD1TCeisHjDvHlBWQ+fp88saJuazC+FiA8ogiqFl54S+cIIalAu46J1EoHs
6iHPxp8v2Q83IhzwBM0JpZ0p/EYfwpaZKCqtUNXCLzaq8cMsT+PlowJ6Achj765N/W3Kae5M/Usw
kJ3w5ckDfaDPgiEdvmwQSeoudTLudbborshwvQY39pUsXJxXNznsH22Wrau3pciPN3JukAIlHdXg
ulQzFVflYQHmXdfTa2DR2hnIUEOOwKPPQYRn6jCxIN91GG5cPWD5SSBfCVBSLbz9JeUsvwL+e2En
jdJaSJd7g4rXlLTTQlEIbf7VIRJrPU+m9N5fxx08lI4dN8qZYEXeJsIy/S2DHgzkg/WPJ5U1A5UH
VQICCnbPrBlYgocmb2Fz+nvS9REs0dS02Vew4BU80tJNuEAEKQ73ZpW2I3VGF/xU70BOytN15dgQ
M3bZG+Op+UXW2cTFl4dRcf0DaZhNwTZYv36STyggfVQ8wouM4NHE6RrSrhnFvjHJ3zflFeyHQqZu
RLgJ9rK9VC8HHbxfRO7bMgW/mZYFuVYhPzCNC1ELjqtmZVPaoxrR/lqpE9jbgi7uUyzZPcOudUbt
VH1UvqpUzpzfpp3pDGJjQ+XjuzKOTjAxq4Nsitqc7FM1yZyLbsCS1ZtlvDMLQfaXtUqX8sZyPNlH
pnkB746WDkQ1CvO0xuY2DgV5G69cg1Y9SJ5lBo9ncbS3viHMoCIePyrkBmxDYuyBb5kwo7ERqWpW
iiLBdcfrrZkqtG6t0gMtBQskmS0or1ONr4h7rHquP1ORegX29frqowC5O3KqiIk4U6cLcmzaJnUs
+ycw0POFUN14lO29LWY0TV8VCDWpgrSaNciBcXkkuznII6XKs+s7rVTwkOESj9rUMcZ35qT5ENHJ
5XNayxfuNGOxdDrJ3GAWxbgbc4BCYqmuQHCpmR8eLwOUgmh1ccqsGbk44uZ32zZalheQm9zviGIZ
VsGuJ5p8UO3ivukFp2ZaTDg+e8+EceCq1QqCj+q6epD+zZaBA1Dw3SScPeqsHEczNOYRgPcrxqtm
xsxWCSzNcEGW268zlp833U7nSmmPhRUoEEjKEvQ265CnnqXhMQ+KFwnDqHpRvw8kMcslBvJO8geL
NHgrfz9dzC+vDioIoe/2q0mRNvylibABeIKjRLHQeHKF7AheG0cGPfKrkYIs14I9Xs63ACclLLxL
CKmMNVBoAvLp7T9V5HjWbJKgO6nA2H3WaYi+9X386Ll3dsSHXf7iDFKc5NI9go7Lr70dprDUyN+E
PGdp/6H/+I6no1h+KLwqT0hVOcDidtPruYWU5hbnozSRTm0cN/ydVx9ulQdWEbg0MhNFklBu8uUn
rYMMYShoFOI2/efwG0LPSvb5qbTQeFX8r8K+lNJYspvyzgrjWxLQuV6OAsaVJdu8TmsIxoBCaBcV
T+iDf9M95DpVJcQMhFIFObekfe49/O2wZ1QY/E6CtxAMS1EZtXti3F0Mq9nw+3AEGrUsiVXRfaMl
3H61vtwdSiIAQrbGKLWPuyoRy/DjfNDshRab7S4GpAnEEcDrCDu+XJcV9mLZxiP0yAcTI+s0xvwC
IOSRQFb0ig/3icYS82GbNCFe+gAPdf2OBwx75dTTZQ8/yfZhfoKhVKWgn+34tJMsPhlOPh/cIDy2
//wqLlOrKubSdBND5i3twxeOS9OYCXMC6VbehYMvwrUxF/JGTG/9VTGGHXVtyW6P0BeiWW7BWghw
4cfJU7P1/1EoOqRjUXYKtEmi7921KFbzaiqG/T8c+ICyFbJwGASypbQZYIHdM+qXICfmjuW7TQPa
DoPlMTZD0N+JMcdTiGm/Nud2GxukYa4JTBRktrAKMlfzDmxTNiu9YqyETedVnvo9yHkXM86nZcvX
KrOTutLJnW2h3pMQW97xjsNC9+s1AR+wZpf8Uiq1lrqooqczPIzpCahaTpn4R+lWgwH8Te83cRF3
/Nz8OZi10wb4xY3gBJmjXF3v775Bf1avuxaSYAfd/nvk2QNvUnkfvH5oSXN3zbrSogAZoyTCmGv6
pwRwcl48B4VwXHZCYnowk334KAEyt/TEsuvSXfhZdQpOraGL6yXNvGRsT6Obk+p4GdkEjsOdB0Nm
EfwnJirLqWRDFfbcJVLIvCflKCpMmRZ5D+7Nlqmvu14Jiyw1OvfaibLRQl7InOMYnJZ2hNAx6vju
NLLhceIdDpRlSg4jF5w6fU4e4TGLOlepLIwBGViNMLy3JCmgINf+Vn1pz0srgIohamUEYbVcEs80
zrhC73AqsZFNDFXRa3Fmwl5L+BEjULMwKd19VPd1PMN4utDSxFEkA02dEBwPqdRzDSc9+DpoeXy/
AmTVt52MAkyk9TsBE4gEkrmCm1E12CyFURMWcwJKSk5HaIIwOIkLmKfmYmcRj/yOKeoPutEah5L+
9g+UZpCHLJLW7t5nO+eTEivK65a40FOZXbqjw2rWF5ZttfOAgvFloRKqOKuvERJFtuSuJNxZFXK5
rswADzvx5riA5QVBNtruBbibQJV+E9iHDh3Ht/vbSk0iZUm/vfqpsNRcovyo/eJJqpuZ+hZQHwLN
HtvhYGLWbA+2NCM2tpw1Go6lyM4+AkrBfRBdXpcZSzDXbXyiMPWj8DKxwd//gqeLuX0MAseH1afH
WoerBlLj9IvOHBR3nrut7xlHdl3RXCyeR38o2okDWUilJEQZPxd+A4dZzwshiVBqe1trACduKHnA
PtZZ3K60TWX/OHWLtb1TWrtXT83g8pozm50zn/7fk8BXbTxtdwx0UIk3zanfa18pmbizbfihrT6T
13iuXfs6OHLXpZJ70wW9Jw3h5ExNxyRYA1QkNqTy1ITu3Uj0HJdlWghu4GpaXdj/o0L7JQ4kQq5K
+6JZimRksrVvHZAQkhVKu6so+LqEqgaj7uQKKNIVkZvwUJd/edoni1RCbY+kJyRGiCMHHLDbU0P8
M1Zo2+FUDC/K/buWrn4eAvZLbIsXllSCjpnfoGJVCwg3mfHD9BWZh8163VRun3HSpW3C0AVZV2vY
P3FN9vqJaUntptIJGabEzSygvf/+X3F0YPgAYL0M7qN8htSVzK2/ku9j4TTqeShdR9OQdIh7J2n9
elSBeTfv+UIw3gQzXRZTpqyuY3vy5+IdxQJcUYcp9Gfnv37a7SQKz71extGRdRlY65/kaIYWbPVg
HRhsibM6b9KhLwFUOlKBWJBofKtyxePooXcSysYqyChqdP0AGqCKVO7bbRHwmdlm8K7QbSljP1Mb
gmetb5ynlv0wW4DkBCAG0we4nJV77yTcUcdBxcn2yZkm1vv7qAF27p2Iy7RPFlhgJW1hy6QqxnNP
aS17v4qkyvsjChCTxbzDGmL+ZS++0MdsGBiN1ge1HuO1ouJ7nwjec3bd7ajLu3jWT8Wvsp0xqL65
iMopLM67yYzJ3e0qyr+05w886mUI26oeHBEJ9YngtlWQtuUcTVkS2QTrLdaQB3kW3byLB7QmzfuL
Uq1BD3PMqHl38YosNR8ee0tdca5dcjwh2x218OnqVDR0T7Qq/wcuZoRUp4fwOv0Akl6mhja/RCl/
AUcc2ENLKhG9TSqIgChNqw6emu5BeJglRT3ibYsHfP6te/UBhZrtWwMzdtwDEol435XvmsOPIWIk
GVfBGhpqyCKgro6YXDPjpWHVVS8JJjOM/WzKklyFiGRN7VsGTePoPUX0ec6ibk3rkG2kjL94uyT2
XL3wTDO5mALr/Xn2yjOYWLW5SvSCPyx426xRJUDhAiUXZv9AA9oVhljqwuFnxdCp1dmmnCXdJKra
gqQVsGpKSj393GdOzZTaHetTIIOMBr1ua5Zpgwp8GMMG6XalC5E1O5FjlNMEGlhbpWsArbG18T/e
GdzqBbOlyvH+gkp6Px7tF8Sg78RWhlMWeg2MS20SLBDaaZ/nt9yOEGDdc9/p12eRJNya2MFqBs6V
CDFggcCc9DXeFITiJd15fYged/olmdRcmE1UeU6phnJCWBcmilDuVEKfWUEjMFd2blrz7YVRMZO0
u32M+smcJmaCv0jOegaALKSgCD3aOOJgg+6Ks5Pvlt5r95/XkLQz57J5AcM+x7fuVpT7+O709hzE
aSjadZfUNhdUn8koLdJSW3/XYmRNsR5TH7ADMXw/SYjTDWlKU6EEIcuq1MlV2yUGA3YgG18aDZIQ
R01rla16yShgQ3Rn9OMDhTe+6RnrqQ2DsJzKpNSjsmxBuh++48kTscHj/H60vCkVfe26cbMGsSPi
Q2Fhwsoh4TL98Iu1GOGfnGLCeLzVQO5YctZbjUT5M07DVui3Q3ut5frR61cvXkPOY4uM6ydQOkxL
CMI+ql7Gzqze3FDJg+C+dhTPPNb/KyMSOGoJ5FepMc1MReCSPku9XCr/PaGeqAQYW0vGK8G1syjd
gSwNkYHzzEDw42EAdVP/aremmlxyUobiKx0ZR/U00lwFNWDMNK+zpf3MJtA8GoqualmHMk7+tY2n
v6eShpdnJadBhacOsvS09n7kS4hu6Di8RVlYsHFJtM3pMZcZLNW1ADRQmyWkxdErQyqx2NF/WMXH
wDhuYMF1FUoKkb7GHjh9mTn5yT20thHLCRestDbg4JJSFr8JWKzeMankBvJhKgb1WP8ZW5sAgG5U
QKEMzAX2oY9/UmLv1QEVmCHirHBNZYFAU5vqlYIohK7oPus097xEE5HRRBh0aVYLEqqFfylZAuem
wQj7Usnu/DPeL//KSAVQyKNufJTk2gzQeGPwsVNZumRkp55VfoeMp2q8gV4h1Tk7ND6ugPLp6PF4
TXqhiCrg39hLuos8tziVAhyuExyM1Zam5hlV/lTocurEeccBO6usi3uwjnUVZpfYIZpXT3RsMEM7
aDcnev2krXJ0vr/0hjsLR+UKKmg6mdxuFwx6B4tfNxlsrKW7sx2cxT6k8n+c5HzsR883mW52un7c
kGsivTQ5awY2Q5NDtIsa0QJtXfffbgIXrA6oDsqRreujweMUp8cv9DV0Z/EiqUaxdlJqrKQUF42p
BJG4XcKCxfzYvYU3ppsc1FPTyRGAeEayFVsHfttjwBTPZ3j5oKU3rnPhgm0Cuht+XeUJX79m7EQo
hE5ioUmtwuJIon1L5AvG9cBweThYhAJrOBwlaidYZ8DuMTu66cxtqMlkWY0EAQOAwCBTzssUc+qJ
c2c9c81XJvYSU1iQ3QW8+3g77C9evyXB04EbmFfYl6m5/0jFxcfWHToHWc0VQQUnYn3XLZxDQYZj
SGr4BFiPqKOr95hLTx8tZQVJ3OASgqwfxDvL7Ff+buLkvJVZnXZvBiMKI35ewSEInBatZNYwph1V
ZidwLsAJgVTlKKFUEAbizXHmh7/utfx01jm59aAwUzIrTVwLhJe6uSkf3S8k36sYCr5gC2ZjV9BJ
Ak8HXlRT4/uC7PT6WVIpTYpoAoMrkfgpCxqcA97m63OTkFERZ6t+Ya+UfYD9BeQgqGF9fPaLCEqW
oOzVcFWYJQq3QPqqarwyu+ECDaias6a6Z0PGSbLTq1UDKmvIVXutvt+HRvsCYwIE98Stux49cz+B
XvlHk72bzoLRQO8WuRG3vuLgJPfjD/O0mbhEuFDOvvcN2Sn7Bjr5Z6EwBswTjn9Y5dLg7IyRrQiR
nXNo6GXzHfxJw3PwBXF5ItZOrdOpYwJcONYz34+JAZI8LSdRqJ/gCanGA2zTReytoZfYjKVq19ZT
D3acET4O3h2H3+4HQcyx6ROuoQo5JF1HKCNzRuQ+0MzKTRPJ8+KOH36qK0Ti5d6vzEdmav0XEKBd
TA58Vk+7DfgiRQRjbrCoR6Rt1LWQLMp1w8Bik8vwzZ71oRjZOtsShWzHI+NRA4iwLLrJCj2j7cT2
4iyuxQt5f68cGOTlrSL+sOJ15yPaaWDnFfG2dYeHr4CVnQHNKj5xl71mrhoqDkEohViQiIy9t3uD
TsDmlv7+HC1g4SHfzEWp538pEbGpuVzKl4XT/SycFx96UO4TRlFcoiUkhaoMsL3aJrJIzpQVVRui
HQQoX7X+iPsNOEMXOdw8DNalYyQVtZ4sQ2JMHpemWjEuXVMNEc2NqckvlvoD/NaLewsLuMP96FIm
gCQTmOO3zublBRq98hDAaMpgq0fW3kB0SR4MrEJEfpHs79WikIQvFIuvqzeFcEy/FYbDnHIGfquL
evDHF9kERzTR6vsycZ/2DxXNrWQf6Mj9jddxHDVvZG7873cCHkAywtsXr5uMtDiaAh2fQqUQpmeM
WQXSS31T8niJODY9l3IVvkyhWdMiJVPB7a33RUZUdN0/DnlE41RXHabTWB7fMF/J01WTFIe2y29o
NiMAxKNua6LGB1IYa53dxWMEEi8f4J8RtTimaKYbFpyR5e9iZky2fhoEKphDh/PgE9I/WE+we30I
fA6KLojAGm+BMWsC6B7zmiabzHgNB11mcnhFVeuA48azxfYdGGUj2TWSP/HUsemHGpPUDssPR0gh
pH/utTQLO9eT2uSNeQ5+UK0X+gm1NKobVdau0q8jN6pp4YGCreULO3FUb2nOTYcj4rK7csHy7jDJ
/+huF4aBKny5n6dL83xWCys4QB7eQqN9HTwqZYvgpLTe+wTLsW2wYQcXXG312n3g8VHDSn/dSzXO
2VW4oBYxPF2CvbzrZLR/aWxD5jZxSJIGh9+4AfGPRUDmV6PlnD1x/rPiBXRQ/pW7AaA8t868cftf
yjHWuQSbWHcWFbtXjxKgtB7adyzOdZgMcF2GWKPboBpY9G4nNtEyXcFhvh2MdzMnL4Gr8no0OX5V
B9af8iOeBv0Q2D18rxQqTbRW4Ko5z1F65GeRO8jPGzvw93YShaPD9j/uic/n5PVTKdM4ZV9fNBZC
2aZrbSKe/wKnWOo+sn4hybWiWSKbFfSPHuULVDJHe72PZgoNkbFkcOg+5A9Ss/nvbsxPZ2zYYTSo
qYFVpOP3dZYMSAIVCJkLAwZqIBDMzEV36kw4K78JGOio4N3DFsJuIQrAZb6scDETvDbEuyMIsENQ
aFZpftprJkL0rt//VoXcrAbvmCVwbHjAZMH6DYFmzKJSwvyY2BpbSXqSCtt6De2nox+R9iMk0fAH
BVWj+/BZjJLkL84OT+WEWHnk9I8JuJkAWnpZ6oq132vB53dbUapCTf7KWD/nvJ31uFxQTy5gKbcD
Z4i3pGiKiAbnFyI99x43eYl3J/fATJTsXkEDqS5d80/LH25avQUN/n9ktjTcktCiK+64VKdUjQ7O
GkaaPVIfWMJbFNIjb7nUHu04yIupwVKoUmRHF371zqlw53gVepmPg1G0IZuWdpLAEyM9MJnXYqVm
3O4VxIapxx1+GkaZ3QfVzu3wxQb5tnpIxIXe/chEapwufPV0RF7HxVM60k9JRFHVrG+aRn6H8+B1
0fACPR43dK0yiPh+HWZO1zUvWrIGRbAMtVWPo7ehcAatn1s3bM5zgTlcgXLU4hLgYzm7HnuHnguO
Oik9XPf2WpGB6xhQwCj7pTC89pkciGaUPAm+2zTBsAoojsud0TMW2AiBLAj+/ZihiANXPz/ooV4J
5lDLxw8ok6YBl9U3BlF1FbonAAO0oXkr3MWljUzF4IfVY2XsEL97Gou6cnhvvVKQkSUbg51ihZp9
sXQfHrFG7CCcePME7IbwKGIxd9gFcfczsAkEWmfJjfnMetbJHAgWV38gNkJX42znlw1Hu3r3LRlD
i+Nt+B7L3J3PCFDjsMIwMimgme5sKvRm09n1UkRaV43XqSvuUflNgLnCqOJU6oN8iJQTLsoDJmUW
pZfqdSj8whXyll/p545ABVqn+ZqjqkpWTM7veVqQy8a1N8RnRGsbD6mVuBjP6lEDAX6QQ6+dEEpQ
DDb2uOSH14aopo+UeGOLcBRK2OMQVmKjOowmMIqM/kBXClmSLPNHpgAVk7AnwXblfgIT+c2CeKvj
P6JOQFSOzYxvvD//3/c8mbXBMTByrJj9sUWuSTzSnI7802eewBrvmYcz1AE5F/56TZrGYh0bWshl
P7NdJ4MMU2nSZ+/Yn1VkzUNVSO+P0xRAEomVCBY8GDXNmsYpTLDHT2q9nJ0SmQDW7WIFZHLAqww0
Vlfqh6YBM2MpsDx2PzWo8YvA3suhT1orwOd7iLceem7+L1p0hlZEBJO2As2adEyXo4RBi5eWoauL
Uo8sUbgmpkg2d7aF2FhdMP9vsYKo/Ff+A9ZxMB6giFifOzBBTB5bdnrbkfjb3xy5LWIkbrs4htgh
0Asdj9Ixk2ChZlA9d+Dn8k6WhXYAh8moat5zOo9vEu8N55jHlwQNPDJnUtV4l3H2lY6WKwihYUBr
ELqm9RDm9alROEjobcmv/Cn4J+6NEIiFsUkvUDQUlvIKfX4k7TALThiuMGycQLN7rVLVSW0SUI++
EkfSTgrOhv0CAMhbc9ZjAEhZNb0FOAFNcVXilElE0xjk0qhlQnocnh2axegBX/qzE5RqcqRKg4+v
EHkkeDEXQLd8avTMhfpb9mkvpBJVoncjio1u6i+DQeeJ7Hzw09H7tKkV47lCNjBJCR0k4hVInJ4H
q+6otc7w9r0htbzHVHJ6Idlr9Vl5NP7sPNURu7g+qSADLxZClkLv+cBsJRz1qHxKgSGU58EslrVq
SBE1GbNu6Eo2D/IPlotgkDu1TB7kXZ6XfTnszGjl4horBGnq+EogYOsANWfTKwMwA8J3hcecCRd9
D1+kmjCPtdca6Z6rQ/GSTp3EPfWoBXcTUc++aAE5mMwC/YtLp+So2RDVQCK3Fb9tmGChb9y+UqTz
PzWFRkPgk4tRnBJIPy+T2t6D0lQmTs5NvkILUJBHlUMZBpLeb1zUx4jqz4W3sdFbR/y1u8e69gVg
ErsTpnaOjjEqwdAqFgGN3PChEu+D0LoQ7sapt1uB6ov62DqqzCGUWx+xF2X8/jCOXbjMLGaKaZ2F
hTPzo2ug/NJkTjRKJDz9pZovcRT34OcF1GZKBAtxBgdg97KdJ4TAH27PZWQqcvjFvVNGB6/VrqVV
aFymar9Fk5+WZkwQqslkx4qlAb3UkAPevBiMQLA05zRC9963lvhQqZs7If7+c57yvsDC0YpJd8OG
NxuscDPoQb9LHUeF64gtNCOS3kTArqOUSLyUxFGKEDH1nndO/Oay1juRYu/ZZzH7qki4agbdt+MD
CRizLXtdYo5+Jb2s9SsCLCo0nj0hpZwW/t+1RP6bzshU2FLQBr+JTfQqY0LAf1z6JEbeEhJDPqwT
y9hH4Txd3GdnEbocjkoG9wwEkfNe7XOhmS7qBi2OhrqIbwvK/eB9VnNqqVGIJp9aDPcwznhrrL+G
z3rg+8z5sgU3bZGuw1FL1O1kAM3ETJuCr6q45AfFyvCmydXk0gG39Lj3Zs83q8lnSA+Wg0DLde4B
zxpuBYkHBPNhqrgKq5+Z2Il6J6fiC4Di36uGqJ+SVTwREpWY6vBnvnE2RdsIbxHmDZLDxF0O+FpP
CESE4UudeW0x5KerJIzDbtKeavon5XMgXndCIBqqN3YPnb5PEJNPO5fYDdUoOO5oPqeopby2OYIW
84gedtnhcKvvZjTFkBK8GQ0xXhh5xzLY6CZSFftr41G3Mp+41kf3Z1yVDVVWU/cdlVtQ7rv10wIP
7BtSXIi+CPlQnGAT03//NwDuHqhtjcyHXphKQfFmcJ0zxPGeVD0DM353Tw0qo5XQXdhvwzwdtTFp
pi1igRW9yXfQGOb3YKtiuI6mjl6IekqtieInucylTYfQVY3QtvJQ6R6z1nwDX6ZZ9ZY9zPLsLJHm
z0SMFrxlhGMTdbKm42VJ1FpDzMQN/DXxiY62NtWUSNRTDoRLa1NtREAQEmBy7PAdyloFm3y+iLou
UltdaAKocSzfPakC8Kq4OSidakrtMCFXJAGIsZ/W54NWCeS63mHuX8qUsG0C8ii8h1kJBiTTE4zB
hm6yr5iJHU5hGNU94YOqTxSHH076eE56FG+U4KGhv4BsxPjCin2rQxPO3ueEjTA6JqPfTeE0X5ZX
rKaZ99FwayxayILPr0/7AzdkJnYg8o/6t9gcE5lgVjljmIiVAnDTfjAI8Uo/nWDDoqoqda5j0KqO
lCFWCxRcIZIHmIpvJt0eTJXDjwJRQEeuOvi6U0DsAcbDdKLwDtN3J7UsHuSlkrdLCva61pSbSNXe
SQ4/olZc5f+6dGIRTsFJgNEZAONFEnDv8L8IMrBr9dAW/pWDgpSXdR/CujEliDUzcFXqFqH+Ky1R
CU7TH2eT5o1DJwClWGeLDA2ALnzH+sUUfeYp73AaPTP/GOkwokLZHqHqnUudx+wNLEaqmN7ZadXn
JOqwJ+4Z/EzKxtnMdfu+iynT3NDp6zmDaNvOO59RErDKWX6D0hZHO5GP61YgM2eWEhH/rLHsMnTu
Td3+Cck+jtHDzNGe49/o102BQPOui/Q8p1Cs+29a7WZXp7023O3BF0nXWV4USuMZszkJ6UcvZqGL
XfSiK67g4tAhGCLbqaqQLZogPnS8+c/hwzu5NF90HXZ1WHOIyBdim/Wtw4LxnOLasWJnquzJchmd
dn2OxsDNlBIojevftBaWIMzxYMGcloaJjDqSv9nsQeE9O+Ln+pFS3KRBDa+DOr3Li7nY1+Bd7x0p
HtPuilj3wB4jl6ra29ceJRXdEezxUMu66wEBqlDlZndSbJc1eZ4u64YCwD9T2rQ2kGINpnu+F5U1
3UQIy+pVvfFYTBWL0G4DKoF9GAvpAokxDinmG5UtldrEXEQuufq2JMUmyd0pWOZjrlemc2d7ypvT
OFA9hH/KI0bVdqoRe7JBl0Oqt3+BZKuGggPZKSnJiurGIT0NDJC/47zGTFAHd/HO1hK62Djsr3cT
b045x0SvcBloMGjHe2+tZpmX5PKQl0lA1zl9veGlIhuhfTWGvCbQAfiqcw1HiCTcJ7rO3BkNtI/E
v9A3Bk9P+YixrCXQ4kXeyDRZD1/fPwlERpt24L0F1Hcj8Qo9MS7HG+Uh8jCq7gPF+F6cg7ddEgdG
qbxVcA+wI0bga8e/zwjHXzaktDSEwf1VQj6tA00QZ3JBRX2rd43EDn5yINNE9GPcDICBSM3a1T6Q
8o79lbuy4TBbniZ7QuSscXYjhZlJQe5NZptrIyAueLORcmhpETJ/YQ9Fr7vlpAuqvtMnWMSv2tf3
fglSGK4ko+5IHFhGhtSGmDTphtx0KxlrPw7rqI9gBn/ksXwa4npNilv0ZQl9VCaCD9O1LL0Yt/mJ
uK92EqRmWPc4j9vHlgo+gnCTT4LxYL1PfVtJoGIelAVJfnVa9dPQcAhdJcFhx6397mszZIWYsyC1
EAgSF1KWadlsOAm0bGBx+YqpRNaXm8nYrYycpZsq9w7C9bSja6g/jpYCB2Yy/1c9Y2xzJU8bFX64
b0+TmjJA9sXaosshak5UAP7YHnalm2gT1QyRJocnBA9NLUfKD9Nr1dz36e4QQzHuhiw2gD+uGK4P
l+lzQDSWGilOGmOH+24dHQZjZaflVYjFJeVHrH61ca+lP9p12BABQL4ooPeW/NY0BeaWq7Io8TJr
RUvWgG0Vm8gxfPkzbo8NV8Hhk10XsNUOH5QQqgSo1wTjUzxA9wRStBzzb0JsBnQsdfW7oTWHpMe6
2Smaxe23HW6ryIXa/hEQpOG9E7UL5tIv51Wuj/bpJq5Azvs/SQsfmyCfkI3d27RHOZrwPvSURRsJ
/5o41lxXb8UJsO5TKw3y0awy1LYOq/lLDQWPu/yMeJIhbX7W0+/LlZAyT1xIGcT5quL+5IQ9mwvz
tR4anljhlvxzxewCX5Um+OmcjaReOEgmdjs2/n71IMCVQagj/U8C+pL0f84UpnTprS9nVo+bYrkX
XOIRkom7iYigoNUd+stUt/8jIxYPStZFyEnmAKZvcq2lA+sN8lL0QMoRjb6ZGXVsEKb7UcVA8Sha
v73K6oORbKwNZZ2pv5xduy9VE4zIm+kdbLK/EDjZRdzvvSdoVbzokqgbo+4XTiM0tGy9MSpFNBfY
zsjgBh1glfTx5cwrMWeQYZnfjJ3hSvTHWe0Y0sZfh2sCxmYpj8cwPaFlvhjbMziEaj8RoOf4gNbx
W6Xi2HzoRGkU0972sblVoEd5JM7qKFHL2JeIFGpxjcpUXHl7jXvozqyAQSDVUnRAEa1k1K2dqMYN
zzmM61w7+h5+uEB8khqWHYLTYF4IPTXFPvN0VJGC9bz4I5XaOlUZM0CsDiaK7fjjg+drJirxRLEL
cI0MTn3+44xX/6e7JmpfKyamVWOhTj1m6TUg5JDJd3jDGQLApQKGvnbHP+oFIvhmgB9EyVBYTVx3
EFXUp17auZEBHSYUc+i8WZI+H789ux3GgexcZaWRtgU+TmaVRG5HAGwcBVinmalMrzMCXIiq/7PI
NwP3q6FH1AKnk3Gik/h2KsrXSXTeE4f9JzPT8noJBPr3Gx/e0lQOZD7MS+BCTy5SjrXzcrIG30Qi
lv+iWE1foiU8vaGyI5XEBll+Y7+sQqk7/XOJgUhio17m3046axD9vEdbI+HhjxDmnwxqSJBSUG0W
pyHuf9iSllcFihbOUAnHd0apNy+Y7TiLGbZS6ctZfcKaItWNSgtKiZZixkubF6brJjAmAeWyoiwN
7ksj+FzPUNRjIBTJoeJBo4OeKTayKacNO96BUJ6G55Q2E9C7WDQIF8EoiIUSeO/yZznmC36YRaTb
b9jSyy4xLsjvYH8VkSNoFkKdXdUlOi+TfuNcBzSkvcMo8sTjeoJHW1Tf8lftpPmGf1YSg2wlAy6r
NMOR4KrZI4hFNsKG4MEC2DceslwghSBxhPMe0sDHLbkeb1J+12Yq+dizprqtb56n9tYEXl+D3zF7
aA9DTzOu5NvB8aCn8O6yQuMrzhcKv0819FnUZObyMlejYU7xEyLTUi5aytrd70hjWUmxbeY9uwNl
kbR1X/opa7yOZccphWbAQgVx9XwcezHngerXGqAr4kIVaWxAaKLqnqWfR5luhzii/kLjos+A0/Vk
kPh4E/8YxsGDYxWCZztqxuYJAIx0LcO4QbkVupZfKk0xyF31wlip1UCtGMfI47I+5yEIYO/h+WQV
Xbh9m4s70Jt1H8dea52RA4bTiQb9bJo/pVS5HC/dz3HvML8rkjpy5Li/zoBDYOoiZ86mKHmAKXbV
MXZqbPnq5tSwjz4zCzoqnl4Q5g2mpWpwm2Rr3GyEwxkKyGlh/6kfK7Hj16oFYPpKohqZTDIo07p0
OBxBuObECvoeG492wL0Ex028Um63ajxU5lqaLsMpPbKt4A17Xj5VOPAWqbhiXjzOyRDtAEYE1qwB
vhH2reKuXinufJqGjvD5Fm9tARhUrRtUNSSLRwklzF3DCNsMdBW/+2Q8wDfEBmQXtP8gnEX9iqP5
n4UzSOVRM+QzVbuGTDysaT24IvwLFrNv51Wu0ZHMfICKe9N+WL/B8sJD2bp4e0sdYir1mNs7Fjcj
OCPnpT8DNCMvcXCTeSK1Vho5YWAWW6MaFjZmF5CLmyLzKlPrXaw46uNPL2ebWq0cFDQ0QWcqvv97
oaWQvM0/sN2xtPWhkP5VSplcfBRrfxbGVLU8kpgougirYxa/ExmnLTR+nbCmnuTuPdg08LWEmj0J
iAp42g6iqa7AlQXZdMd21Bd97UtQrIh/wJftGrBbzGKWIillK/2vETuQ4QYuSf9LD+aepxa6IA0u
m1NpHrZpirijkvT5Lgshi0MSLa2anpx5T2BUrT4VakOLYdY9QfTQjLjuaqcuEZF2fM4pcFnkGA2M
+b/PnfAECtaj8tZ0Spqx0WyBhNArWOMZE7IdGN08N1pGXjl+f028xt/O2mDieyxoqsHPYeLYqFtu
EXp+vODtEHPQC+voEClVkApXytbULTL+BUE8RvvsbUpcTrEjAqKmXWWESMVbEe+OPIvqjg1J8V4e
g4OSf9I1WH4HtvfxtGoKbo86grkyfPQHs4NKaEQTs6HII0qbdzjST6VHBUdg+0p6g3RSmbf0NI7E
99B+bLSGnC464V64hx/z4Z4Xtd765Ry5YoeS8Nag8EF3fP5YDJf44NispP+Img81zKNENipwebV2
UsTJiPfFHQ0QTFzTyZGTlmlrK4oGNy1wxXTv+DP2j/RjZxnIAMW1QAz1oRj0fRPg2CbfYVmfrxwa
IOXVoOvIoa+208JjaeDLoctp2nhfHdMNqEV+r2xelBaeBNLDo8Un5VytAGSKnACWao7KWGWwWYBt
a0EP3tQ8XgZQbd8bLHMyRYQpkxTEx96nkuvgdxbCHFsuR4Z9I7HBPLQ89WcREQaVPPNBTQzhgQ93
7bYmeYb7M3rtyR4wLVgw2OWZJuvEzSTzw3p3W8PKaSSWU++X9hXC+LJIC6aDo02E0M1ufKGG0Vq3
RnKgpJJEfnDjWQiKtVjqQK2eBv2r0t3YreWkZur3AgFHdB0lY+DqVtYR81mUnId06J5ap4bneOMV
4+qbDE6RibmvzmDm3utxz9zSyZa+vZfLLs1eyYnLhgqMYW2KHh3RIVKhYWrA6g9LJVl/61XBxorC
i3TJ/k1PsZm48F50zgs8fWp+rBSGZZJkrVBfaCz0Jq4u+0ZpD1G38Tqiu6Bjh0RuKcickgC4UEuI
iajosGjADlvyUvg/6DM2zkwOm52IqMCPWtVl5mtOYsm2GfHeTuGy+Zw6+4AWj0pyfieSj8u4oQHP
TYissUUjZ2bzD0uqzZMNL1ZCSCN2T2t/nZju4yG7zc1WpiOshI0Ai83GuAV8Lmipi9qG64bdv+T+
CYOcKlgsbfeREB6ixAF+NirDjeKtZ401LOwHxvsG5tUYWxKQqPERh5vY7VdyX/V18rf8ZWzcoU1J
CMxuEl9ALAcM+p/mzrvWqQSMbDvxdG0Kg4b4rygIc+9R7J6eZGSfeRKMm76dmU1GPOpO4KdApG5d
52uHjKqua6m7wDWvfnq8uQxjG3YzcBzzpqn+jmcKuclZGE3sFadCUNwaaC+YRoQx+/TB2Dl656Vi
uNSdBxNNupvtFIYh1txsrNjriq5fGodpe2hSi7X+EvYX7F0e6Jny4f4H1/zYD1EXz28TtbBRUoXP
4/L5N1Ir/+fJIitqYJDRc2rPCLNJid0MV3Tzl2UMW19CX1dtg0Q7DsuApasei/CxV95bLFxE2j0n
lK4Uf3Ts5dltmED6BRN2nCzAGEgGu2Fn8WLL3TcrwXNXPwinZmnzuImmt6SRaMe1zUa9LsIQSaM7
iUvZkIuvxmjjSBIz8MWrdmVhm/mr1XB5oSNeNGDxdFZ/TTb3xobzeho55GrGsDF8P/Jh5wc/KblW
cjKbKFaKwQRzzzmmVJAO1Q9X7lDlEBhjTrzkSocQi2S4KfuCraToIDUoZYH66Tpto1FSAepOKunO
qPxleq2APRQLZg1/tpro9mA21qzZu8SS++U6y3fzIB5IevA055Dr1YZS5u9dS3ivRupmqXqeqh1O
8Vok5mrTy1+NG8Pc0hSNhOzXQKmcTNyfPO5udYMfy72VFdzVMuQZOIsGMVGsMqj+HQWZmtNCtk1Y
/w3JxNytnwygbL8WURLo31+sF3SCwsKLS5Z0p8zX5jKsQ8qEvicaMFPOPTGYTIDBzB76n51U/TGL
lg6o6fFALKrj/cZPbcr4vBsbXbZ+GPhIT8hb0lNtF/bd84iikl/XFenk0rhL4BOFS/9PHu0+b8hH
BPVWyDzcR89lEqv3hGytXQCj+1fmBJd8ejygMxk1ieWV9830MSdBqv2NOX2cSrNA4DNlXcNEuHv+
6YZTKt3ZwPBjK4btoMspKJ2kJxk7/EIJrBmbGdMhEo32Ot2NzncsAMjLPnpEPjksuAZBY2davq5j
lUUzlsM+L+XeolkbZwoEZoMrdjpj19giRq+3mt7DdU0pzttJMY4hzAyxFisLNLUnyFmbWtDHY8OB
bxlmrYNHc1jsXPx/SK0ApsN6Y7iOUWOVwY/yXe09aTlG1/8s5qyEeKmkJu4AksHjL7Ep+5zFNN/o
Azu10kwqGgLkulwmkeDnAqT1AT5E5UZrw686clhKgEaOb3CdBLWlmgJwirWdxditj8GIIIY1St1z
SMbcuNJHnN0VQLYVLEo7K7BCV11/8TYrJpStSzRu9egFjPX72jEBACW5015ZTpRcUGy1fsmBpfIY
Ni1GZSqAC1hg7plP9PKHtqXohgca3qB9bA3RF50tCln/EcgIxxoGMnQctnnyGKApM9bc2foRc/z5
Kz2DIDxWLUgg28Zct68ND1oLlAQH531FZjB5XU8geeJJXjNiLcxEDlLblQ+KbKbijBbarYzY4Ey3
5LIfVlaUKqQzJi8kDLyLB9VgmAQNXuoNMv4gILugEd9aMxjCgTg9Q+UFAJcB21+J6ulaVO5CiwLs
G/Qa+92E37Saxz/fkg8+jhpYDEgGZCgEY3CgjnuqISVZqp73qQMHI+iGA/hj4BDhsQpqiUce/qd8
WeHrffadImEkcRDHP13pnd//781065deKuCdaqjBZdAlnBah3/8MofAFqagbQNrU+24aTG+Yt+nK
UbJ3trx0vGuHQ2oCbN8+7VWb6uM0MkJYhGxVYxd9vmGg+60cW6ZGAaUZun1gHpv4yFJjPaEYiu9B
LDZWDPFiAw+rEYZmmtucHyMDeGt9B4xueBoP0x00fTnaUbo/uREk55pL5zYO0sY0euwxaCL+Qhr7
TqnmVkp/aIQ08Yyz99Zoz4xuXFQz33bHnQ6Z9UHm8+eo8fCkhN7oAvkequIAN1YBfFo7VVWB6CUb
adz1ETiKoSsgNje+0bv3TjEzmuEN2v9LhR0l6dEMo6xf7rO97NL41TiOsQPn8y+qF94UA11tfrpG
egFW0MAmxvBUlcR+MUTTZzqeeIEsNlE5i3DbmuZGNmOPhqWlJmZRoo7dISicAsGPqOVx8JZJxmuu
sr1r9cXG1tBmlDYBFb0rvtd+/I/S7QFTew2V2+s+3P/hpCN9MVuKFuLihvCiFUSAwusSEJN6gfZH
4Rj/ij/9I6TyQeUpADJESI2u2VJ1CSXlc+2H3mVtQCYrTDAFqSxFv6G+iDmDZHdfBNSsNJnDImqO
Cgr7iiBOEn9SH+Wy/SDM34uHrk3ySICY5wcmurkuVvd81XKjlxHCgwvWfZI4CRnTLVyQWXD9gbbK
hQYkiziTEqsF77Z6DTCbQ06Gp7kcJ6/kBH7ZtjNAyJr5B30Y/Px2zTcT4wkp4z8XVZt6n0X8hv7w
kncgaOrR8hd91D9a0jFPV5KZdTpLPMYYdI5fmHmDSylovYvCMjV+ixKLICv1LDOM8TxzradxKmo7
Q71ev7cj317v3+WtiHAQ+NY5fvdufkHREWVvyEulg85GJ8hXPcEzUJO0kgBCDtxJ24bJd9UJLR1n
LvFIUl8H9acALeIIE10e2jU7iGouE8JT3gidLzWb39ZBhh4HmFBUbNYggdIWCZo9OjBmJ1k0jtPX
hQkPMLchzEdpAghxWgipw5LoF8yUoWWs5jPRNkH1w8XiCSMXyIdr+R7Ks/0h31/5eegGiYEorzgO
4jJrhxT1/YtYO7EAXfdwJsaF56BdiZXJbxJzrFy4TGbdx0FdUqd0xicYkOWPgaGIxNJBs3mtma5Q
SJqdfXIQd8UD2xjHUmue5bR5tpUpn7yw6lTHRVSk2Yt/fTrDCAxFHYKXN89HjvX/m+TgrVgB8EB6
T+vwt0VmJj5k7lQWyP+uL05FEzEJlCdVNDldjOgmFJy1diDaE3di2iyQZ8QrhOXfAxAZFvcdwQz3
cjUPMZiGnEuXpN+ZwuDtOnS6mo54aJYlPftlge0IX0uUEcoA6rQvzRchvsyB3iisIckfmBDKfmqi
jkWx5pLCHkhlWUZ9HU1Gel0NtliN67w3ru6a75kat3T/DnHJss7NxYyA7sriPoRJHCn7t2wa8Ede
WaIfbI6nVYDTcs1nnYBo2xmyIzeYgJRQUQKslAbvdZ0mdnA52aRWWnTQ6kgm5mathNWnFEoAvKtb
H1yzGfnrFxE3eq3yJS1t+hEu4OlJMLHaM6Fj0O12bSIg2j9ZfHljALsxIlUwCl7KeTqwo7AuKeXM
DVz5zJLuXPGbQN81UbbiCa1wLgXFIh+IJzC9pVumXNyWYk0QPs91+oNypYDOWZSK46dRB41Acw5w
ixSMV757SxdtPRYJ0sdJpYS/zqVeqCwgrVM23CeYKEo6P0Reabv1/tkqABPC4ntCxS9XzBPw6M3n
wTBJT2YLabuemOPJ8MOj3Fij7/MU29XKhO+nKEqL5jRwUlS4Vv18YZb6kq+RU3MzMon5UhIdzGuZ
O7Q6z5eNtFjh+LfNqVwLCCYj4ZEoW+1ef+hSrf7vGg8BK36vY8l5yWICG2Jf+agKZKvC1+9iM1hy
5KF7bmvTmrhMNMOwrNv0Bqe3OW2+Bfdh50nv3q61qvFGJsS3T1SaDnaMD97EXIdKz57K1Z6t1REu
1AbR5mlMBMWkk/6QjaXstpV43npbW7oiAt4Ccs9Ul2zM7UXx0vC/cGgzgpOOw9qArKiaphjVqmZ3
bGIHPY8VUaIRDd6wsNsWumY/PXzTX38MIXyEzZByBSV0tUrIBl3l1bWvHUhTEMd6SMeD4w/gq/mh
U885JIJpZCdYZlFImmp2MJppJKO4CrtGxZ+n0IVbekaVd8vkmT1ZOQTgbD8dzJJVAw0oDWhefctL
m2D824yVCC/nLSQosUdn6qky52hT6/XqVgui3YC5osM1mYrttv9bX7vB6lUveOcjjlFjrwPSB3dM
X15KKH6iPGnA0/2t6db3JqVjJovrqHZisoqGU6mLDkCr1ancAwa5o5zGspKkBqOIvn5fQ2LVLUT/
SYFJb5+7TqibwoxRpuF69IPX5gesrMjZluGv6tKf71r9YzGuyBTbmL5Nq+qTZRWH/pn6Uim8KCS1
ZeiAG5LsG8PytWz8NounsUiONbiWdxIon9lCicZ3ZYZOPh+kH3oy37V7/OlAqMxuDvzZFiIFDNpj
/5mICUBNrtEmpsKdJCbOzopsRbaXzsAL9u/5EMC4GHvyLYmfYbcYw+bDrJrlwUTCjbWHS+AX7P4z
J8ylCwsHbWbJPFIZDDwwfx1+XwW4vN7RjF4hQkq3LYkMm9AUsrp683fAkRm0o790rjgcUTEkpec1
ttvEPj/mNQ18AC+RnnpPcVI3dZ6QgCozA+6IMHEiUWNrpo7/m39i6KIAj9vNcJ2TsiccTT60FqO7
v6kxjXvVk/uHDLOsJKz6I7fnF9YcbKLgrSzDzK7yFanNIVN810CrV+b3+07Tfg01D5DYIkXmb+zg
eLUFrEwsiuGvEoX01dzSb8DEU0sbMCZLjYpfc53hXI46TIuAzOGZYGFFMcWH7V2FdjWkyu7VGjbE
juF+3c62hvByuPD7Y+9HPRqkcPqoWuSIkHi2jQ4qa9b8g/ZwGovAZAtRUECjkVCOIqrDVcGj+n7q
+g3F4dnOWa4QzKlrXTomtkCEk5cz94Br16aG3xECkVrx5wW4yGjtmo/qkqeSfcsXgHZ4z7DJQD7D
h6e1rD0JkMLYvTeLYHlAVEdN2aqetiifEH89UJ2L1Y9YRmPXwvQgrCtGwIaPIAXybgg7SHaearMY
jDRfNwZ+83cdp5wQocL0R78GBNCQ4krCqQW7m5bkMD3rLGdB4sh/s3FSoP72o3rVADtz1bqQflyI
/wi/lC2un1XUfT0dU6Rp7AB3nj723UXmrZawGIPJaNkpdW2/q2zYnAcD7tvwUfAKyLlkxFro5VXJ
8VDlfz/3GfSROvSsfxV2XZCG0thJoRRZks2k4Y51M0+WbKoujZFfNeC9YE22n3YcdwKrQsffZCtx
svHKj/s+p9DpHB934wjbu1GAOssZg94rHlL6DXRZu6pE2MbHK2o47tJ6Bo9qRRs3fBtiYTjhcuJB
auRFXF7KPX1J5EQi7NbcpLVEAW+587fBtyY7YqBMNj8l9+sP2KzRJeGtzHvd/ERPhMWhJHSlhoxD
IuoeVCAKcbb3Lo+pVCAKFLAEolOMDLuH7rCTS8VVhybXQJjTsZ3d/7vrBgWsPvvb13L/C5CEINRp
9j0UTzwEauFhrNeMCWWVbaXeoJR5ky5YsgC1U820dOBxEre5XffgWDA92MfbGKpMs9OSu0tiqdj4
+AAQXX6ujIsw0tP+/LCS6F2PQXm4p/AxoGMPY45fj95IMPKUW6fbwAHM7ipZdyTXFC1QFz6IjHTK
IH7yX9yJdH2h3xohUeN7cKbs60dHCVqznRRyvk65soWGP97C8Spix4BIferrx+hmDvikNk8QypPS
mUamAO6XaYRQSivdysMV9I86XtK3H2bTzijuPfJfkQ7H5Ci4r+xm6tuyW4ivDPi9mebaljYO/OkW
kdAnATsVk0PMaukQnOExtk4DgSAAhJ1fuYgCB4iVhaFXtHHHudGKcF39Qyhmr8Q8FsuguJjplofX
+C0vY65AUdQaUVoAMZkegXsvtOM/LHDpgIUq6GusEF5OafSjGGotZ1iAacQHpIKgYVwR3KCnWYyL
nDo50k/QE+gabzfuUmaBzTQrawf/hnHsmpLaeTOtmIx3AgJC4sn5wS8gWUdecDrZIFk5kZluoibi
dUrxBlpKejFR+W7Sw7puoqhFGVNOADhXPs7k0UUHYTtV02NDEHzJe+APwcIkarrLoiokAXHJ6lns
l7Y6Wtq3A8/uaIZ8YXSxYpm8IWT8sMKSHz5iVHrAu/Wck8eiadsND8zBcen4fFnYPorGtLfNh1dm
CM/TcFr7pKn2ydFfYoh9xinUt5E8qqDsP6RIY63TbXQ681tVZoaJzFk8d1dsAV+sJfxR6rUeTuol
a9VfM+tID/CuiyaFCjBPhIrudQ4Y09PLweDvwFOQK7IcavxAG6Ym5SOUK8iO4Ic4gi7dZocRJ3gq
qyoGlryLelkgs2xw3PVwM0U2vzKCuqgfH+RIseRjP4Vtsyq83NOFqfP7HOkAI2KdlpG7tGoPKN3E
s0VvHJB1I1RqoXWBW0flGJpG5oUWsmZMiGWFBh+ZsgZSCr5+necKFYqD/6f8RIbJB7gn/Y7Yvelc
cAGm+WBGUtMolxQ+5a/cfqNPgPLgbm+jTLtXhCqlwsqELgCxcxsOx7yZ4f+7KuZ6sF92S6eNWI89
+DfyGi7nfhCAYwkdbArWB1ofkHQr1vsGIhbntpgFbpFQE4fv+phP/io252PlRsmTw/5RGS8UeStz
y8h0BJsH6rtqg332ouM8IrM6ihRZSeUvszNtFommlqIMURdOQW8n/6Fhy/VQSgnsvPC5tC8Z/lXJ
BLqbYw18rj+m+/dMq1vD0JpTl6IitSWwZ1opcp4LpVXm9GCWhIPPs3gCY/d2a/TsgpQ6u6I1rHac
v+GYk2CFKOgu0Fn5SxTVYfM6IpOSu3NDitvYJW24QPabms3D0yaM55/lnP+xSr4to4nwSG7K55l6
k8m9uCiHe2xFuPufPcw69d/jhpEcx4WS9B877xjCUJMndyKuYWVymtNYmktYq/iOFlLDY/+94Gxu
nZauhU2X+zyzn2O2z9nfJzp0EhtfjiTGdv5yQlmXikLL84roSOSqd0XuoBQB3w2khRZeezLVPW/i
JEhc/vs300mWuMvR/wEIG9o/4tlqge+iODuMMPcbYLnTbYKIh5uVyA4U62VubjbRAlmgX3TrtD2g
iTpozAOH5IP75GCV6wUfCpAyVkB+I4lnjkGiTOJN6NM1lrrLNqko4lvbpS7dCrRIfEngtefmPm8I
+0NKR7qeUV4AKRRLN0oTAQuTPweHKOgpfGNkw5teQhknyK7FftY0nLkDkC/N6N85zi0Qllph9wkt
NDf6jAIo6QQupR5HVaWBoShqrryKS9fJVI6nBBhB45uFBRMS07l7JiCjeLUJc7ooAV6EEx0arpM+
KToU3ZJczt9UqD6DP6nABdbf49Dq7i5lzxKcTLIbQyhHSFs4XDrSlelYdZExQgQQ33vwgheyytA9
fmWrL4Myvpm3AoB28iRkQ5siYNxh3ZJa+COnS252yoXoCS+t7YzT1Z7bWKUxSw8ZNPuFd3H2FyTW
+ks8GKhicrXIhdGFuyofSQmeMTKfrHDbQJ61VOkpTd1kD6MGlStxMBqbAyfc2qDbJOyDadl7CkBM
oc/KQ84AO3revo+rtHBLCvGFatOTq6gzu2vhXpKPMEIp0ZRjhgwlZzR/sMaZZnpdrI0UHa9l6CJI
xXmuYflzH6q3JQNV5qCOgMpoNIpErsclykEZrG2t/3sopZpPn7Fis//HyKrUnHcVddXZHKl7EZh5
g2g+qyihQBeiIIKO9msGyopOSDkzVDAmrEvNfIMzrWOTaLftezlMmGaoEZQP4tG2P1B9r7K5/YfQ
NlEUvJ9cs7CnIK2TyVUFD27Gp3zOUol8JLb5TVP1eQvbdqwEU7VEX95rIJ9smYf0hrDVDjFVVoVa
TXB7F83gDZoDilp8ySbMCLIryYe44l65pqn23XNBn/RR7Hx+waf1BB+Az05MhNwV5jjXk0w3KAUk
YlOuYmZWv32GteR8tXoJ4NTu8LweH7NMsJxO9cqYRq2sRJoeZrTBdzhan2fSnE8Wj5odwdZOekRS
7cC7tU/cgaUXSB6rPesP1r5BFijKdAB0/j1bZCa0Wt/bRr4wLp5t1+hVf1Ja4aCEClyWZVrYV8gx
VOPiIjSnkywJirqVP5vcsLDBbnTG7t9ADd1gl+3u9Sz2BqWM2TlhHcrEUP4U5/qC+ZAi9CS3RuTj
tyFtnnZYl/sc+ryxkxRMkkdsdt2XYS3MpKKx2uWwefeIk2WDOrUFTLQ3Zjpyc4+S04qIg9ly38eL
47E/WUXDdlxzOmvrT6AmnYt14OMcrH1+7GOfJjG8qicPGZBM5TbAxuELkmqrStmhQdEbhchhcbFB
XFaiZlThh+n14P579A4457HvdA6n5moJ1eZdszct/kCnbQDonqD5czR5ekq0Xqej/ZWcYpA8dx3z
jHjx7RL3YocxbJDhniyWGvYGoAfWLpASXPxgG3BhCBkt1B7NmCxGlYm5VkUYIvM4ue4T0rde56A8
wbS2WrxMQaYiQdwIB1Z31IWz0izG+7WvRlHtSx1QMu7wces4JPsVv/mElS61MRsniqFyVrYZ9zS0
p6FyQqtkbpPAe7q3P6Y86KTO58BhyEWENBsh1c1E6tP4Lxx7h5tYzLkhCq0uR5ArS6gjovkwD4o2
IVPq38aCoM2jY2SETRybKNkv6iPqDaljO1UFNLzeZ7Y6hc8APHOZrwYN1Iokh6pcDgf2lH8rSBUU
An8Lu0QU+83z6p8xHZvV3z6BbbG51ELJCVqMkIakh5uahm+fP6IFxprLQjZ/E0XXMmmF52RQo2XW
/mSETJPFBfWV7r5kGuFefVz3s1/ch0ARs9EJBVViQD3spEr7fU6YmnsEYU69YsIWMqVvtRBJKNzq
tm/Nwjguyv3t6zZwC2Kgu++IJIvo982Q4PvcFcZWFLnVPdQFuzMMZhhE3LUX6BntVqpCErEM1bXZ
Pu1XVULONeyoldLOpM8tuUIxmTWI8IF08oOQ1ZrFiZ908lhYF8e65qmAcMRc3BkR/oWgv4e52jE+
Zpfb59X7u+OGhG9OA3SQN2X70PFTiq1XTi4UJj5gaQUgxLENsZM88j7c6Mjkmgv1ubnLu7X0dUQM
bwbT/gPFWXMlIK3vOAqwAO/QK7NFaJ8rrQe7uimXaf1vT3zHXSrJSv0OJDltkYlvO2FHT/c5+Uu7
E94iR8VNnabCW2fd29vgaNIBilDi6NwtVVgWRVrNPoqSe1IxZyr2JcgIn+/zrwQ93Zak8nQxGncP
ldvc48o4LE5qs8o5Z28T5OfRC5r3dyVIJnEmRi955ZjJq+NBwJFcYsGO6Dc+PYBEoU6HauZwvnwP
6dBFSIwp4knADHFMMwRKag11CFjE4d+QHKywqeb8EVyQxi5a5Yxbgheg8zB+FRqJCLog5IdTX4WF
u1hZMIS5WodIHhP1D8CXLrfj4y/kI7Tyza96wEn0UKAMMPXeR8V66auhhPFuc1ALhex1XNph9AKH
H/+vsk5nGrlXdnpv/BEjWF8n1fCFMKm5O0erHYuFRYTJyRFor0kjzApxjpWISNH3eyUS9LCLmea4
nZyfks6HtdCc2FDmYUkWmSQ1yITZeM+tKpvoz8OP+maAM8k0wekK70Fnqf50Prbq6+7dQomI3tPI
xdniYfbiURRSGughDBm/fsffcN5HRfB34LRe/d+gc2BWt6FNLZ8PFzSXLxs/X2Ym5Sdg3k5wkGxZ
QJdfrbkxYbL29L+BeZfz8HX27mJyMKLcComI7tyytxVOSVwcM+zX5cXCEp2YKgFKiFHNW0qDwBDr
EVg3j7GYYl7ZvzQFdBIIYuuc1XURRXqNZ7cVSDg920b2I3x3JaH0CZhxEoSjUCBZTxeOEtUmXf93
+qRmzltw7ymTNcRaU0Z3KjMW6JcqwbzN/aklUnzmW6xWZzRxbGA4NF+/HXiteGawvelmqCvNIOFv
JDPJGFoQHOmfbAywcSExJXAlfP4HAMpXCgXmB9GQFUOUx2QMEUALJBoy2IPJVeSPEN36xQrmnKOa
H2ENMuy740btmjEJ1RhYIivlffXr1VSToNXCkj93paGwz7DEoxYfCm5nWk8eObSqUOlgWT/vWTw8
aNPlxjG7GMl/1pW6IBHF9GM2ldMH/0EXkMmzTBrxiTogGEOoK++d2PYMXSlQAwTTNUj9XEp+Xuzv
E+ToS3uuan2YUJfCwzvrKBPJGou7MOK+J6ii+6FwTB60LlQYpmH6W1hqVseU6NRd+N43Xn3kt1r5
muAwXpw3IDdYSYWsthZIhfb0BfWW+iw/leK9Mox9bu/oB7ntRRvO8ki/VvKzTjGk9DNrudb+ApxV
c6FplxKotZS6kf8sMstxm9UXHVVxeSZhD+bHwEs478tbrbc2o8GtbtF6hQ+StB85zOCip/oYUw6t
y9dvchuoa9VkLA2W79hLi2+Z4spZPeY0dhhlxtkbNH4rgdWCSm6Hh5xfiYHyjsOQJcLNYwgJDwxu
5I7ihH43dPNMoT5pl3P71ZN6ULBM8ht67xTOOi84SZ2BkYFtgCVbaiFraxtj2ItB6IwOmYMG35Fl
V1DgnxBhXQYOmXvJTeGEkZFrPenBxFb9ObcbZxyuq/LCgfeLe8nhv/veQA/in7EfWPb9M/xuzvl0
8YIpL9F9uvRSn2/psIwPu85kP0e9PHruC7rOX4DuK83Z5KmECmcvhlQMThnfAdXsOvyiDc7MNoyC
BovZhIKPOjYfIs2YM/4h5cKS1pZgTOtvBCfNtEDqTG0a72icKnfRhCFahwsnpQEe5E5Ob9qfWaiT
9F8G21dNa1cKhFct0PasljlQmXWgA1jrZxWGCCcVkY+uMRW4VpIk2b9b2KO0UrJIb73BTSLVywDd
WUrO5h8bs7NiCfMes9X5AGFrYYrorKXHrou/4vwYWe3lwlgcd7de4ysy9mP1GteOzqfheiwrfu3D
ns9iASfNIsVjeidw9yMvck1S1c0Y6bod9kDCVO0t4fBYBIhDtmZebzBU31YpbMc4DHQzGvJhg1R1
yBXOjaBv5L6Jw6e/MYthWdy/0oAM3hlk/86qiROceTV7qZnxZeCi3lhm39JqxXKBoy0cjJ1ofdEw
xMPD4yiv+QGpQaCoU6iXEkVw+KhEE8Vuuo27tmQRHr5jA4fzcTfl0k1v1zZrAltrWrCfLG/6tk1D
JVmkP40Ia6eB0dNRG/bjtcD02PUoIjMaBiV1yDwnfn5jTIQPT+8RDFd1V6V67HcbjL5ykCCAIe7U
pdXcjZVzxru+WzI/KwDuOxAFNOEvdJfocFgmxoM8CynMH5lQR/EYHC2x9mjmicb+7/aU/+dOuTi3
spribGzyKRuAQ6rL/HF25AurFHAMZhGezk01/wLd7Ph3Am0nKjg03LQ750J1FXZKyhFQfI8uc7eA
JTVw0GuGvRf7M7mwM2lBhtLkWCdtUunl6H1omFln/N8V2/fyaUzY9E3oR1Jqe+DG01Qoxb9U4bEB
mQfUH0fe/aq3TKjl2FDFKXeGXIrCSYMduTJz18QkpWu5TdIobCnj4YvGPuf1Q7afspa92U1jVd94
DmX8ROYKwR+eoI6w4mkcHAhPgminUkVcdudg+XpYBe5Nak4ptd6VrPxR/psxg/IS+kb4c9r6NJld
tVWwequGPJ0Xx8aT4G8XCBmzSug8WjU9DD2TReQtL7M+gDSHWna9fVLRO+xfdvTjhn/qqWhFiOWM
5dM+JEfj2aIvp8eAuLQ6F4o160lC+Mb7oCxwa2Un961NpcmrRILH4iiMoKDiKQR+LUV2MoIPgA+4
oauoN6hKopJ++zyqstWqhGT1f7WLd6a9z+NdLAzMEpfDl6JgQIZOxvp6BYI8EsI84RiVwhZ8mjEP
LFLasOEIMSF7lDHMpni+V+gwdNK8wlp+bQ7i1ylfUCc9wEvoWYV80F0woImEZTUJ1wRfNung5dT+
+7Bbp0qxd+DnjS7WkrO4cBtzfBMm3bGmJBAt1AteqClomghQeS+AEuRUWno7sicYtTDEjxZDd6gf
1cn6LLOsJAA1wH/zidEu2kXYO7wEBIYwB7X9sMvWWRx6WmLKOYqUxYspog5t30WQjfyTxSXkXBZ3
WqnlJIXvMkYCg6QNOJVzvjH8elHQCxn1S5LmLupRQQPyDt9ofgygIW3lbWT5/X7LFdmDvtzZGYgs
SPrIHC/5xJC4S2jmtcMXQTp7gek8iTyisNlP+m6yHzOzBmiEi6QBV9KPgJtTYR8qhxX1K8adV49b
QA+9ngvkgWaC6Mcyq69tVeLN715bBWROOUScjB7RekIL0yUVPyY/E8ejHXDGoY8SPeS2smsKDk1x
1ZEwhStAihP6hrBw18aTjWihb0RJ7dipLspgMvLVvLDFtaCxUUwT/4oYEP1ctnxWOFsP82UEDiUk
4/vcI+6MiF3LlxSvCxckakY3mlz/VE4Xtt/76fJUyh2A0aFJieOViVM4pwYZeFCRVY9EUCCSs+Vh
VSKmfTMe0sNd53Bst3rAZeH1e7I7h5+i/8aivTyS/UayphzBephOyigv7iZQzRLRvtYBWpwvqwvn
XCe91GGn49GEpDrTPBbjtlWg92lZwFGIHaA5EZXAEGcZgWlNtzkh+UFaxLQfvLkTQM8FuLSo+Zm7
1xtT6PG8tQi9a2jauxe7cIdwfUTiJgmgZFnScrObYG0/yGXMi4KdsjtT1c0Aha36rB5fBtk1MmPI
NqXV/IaJ++b84wwaBpwIBxts/iFmpEBEU7Kw+RhcBAKVQ/rN0kPAAJsAMz5JOenmUH1vAiozYPae
GmPF6sKqhJNwPQ1W1rsbguxQIQdR8GNH/TwPPApJXNkADNAR5vZfKUOKiS9Vy+HwcmhDw0/Shv3S
2M3WufeFjOjoHeR/TIbuJOlJfVxoqxJfTLTGEnrSFADaAPjhIDWE2ToAi2sZx2urTag5akwMWozd
nQw52QUiswP0bvaVAfm+O4zl4DB45y/ltioITP9BzRJY0OkZzAGFNiUzjeG3NY+Au7ogm4tF8weZ
VnWsx+dqmPyzAmDhqUZC6CQioivZVbI8q1C/R9KC8JwiHXwrPECVDVaw/cPgBnOsXZ4yOkRWEdo4
YiG3TJ0KWtKLhT1uWNa6iwyPGqYKHKhi8arxc0m3dLPyEcLd2gFG3iVEt6TLzly+QttX4ndQ5faq
07GJX9FmkgWfw5qkLXkaRx8TnzV6niBCQhMHHNWEDwBkWrnDsGY4tgvyir4VTIo0hQpfGBHTcXD3
ZbFtjOaEzRNP4mYKan5MUT1rEodbqCJ+KCk8pyP2qLv6nqubU47UHOFKfmvvWV717bCDbgoeRvQS
3SwGC6Ndce1eCX7YmhXGvJbfIJmx97rn2DLJhbed34inQssEKI8jBlLuVsv/HDTEhjQVZ+J/BygX
ZjXi9otlroehomDWrzaepO0sBnNqpnjX7rJSWxbM8I6EKjyATTom0L1j44/TfL6liFZWr30axEYm
uIlLNfPlzaH5AvYtXKLuOKBgdpjmuYQtpg5xSaAeX/hq+1PHFEmROkCtbJ23lImhgPPjUOKFxfe1
982UV8oOpCp1mZBtE9yzxlXr2ouB7FXpnPzVXR49s7IkP9Akyhn+VlYglXbQZofm/rGWRtaAudfb
Mqhr2gyAv9XrKhlmmDRxUvyFJt0YT2C0esCzyUZ6OLp4u/8H1hNxzVKCogR27GdHQcjCHWcsCMFd
5ZReoX9pgfgLoenrSJ3wWTU0zb7heWoJGJvH/QCWui05htB5NbwT5MFMj/RPy9vMyqEN/WLABllD
VzNQEeZVCgkia+fj0BeV171iPB2cBwan7/6JbmTQv87Vg4gPNAd0NUYy9ILsel50/pvHW3f0PGcT
VeuSC5pYX5c4WRtcqrr9GYttioZTvrygcq5mVFfyY4qftfBqcvP+lrPwuA8CAA4iTpOLdOithc/9
cYZYyvApC8kLt81Oz+OPJBYvO6ZDshTZF1JzIdHOkWvhKc88EZN7CABnSL7jwb4SBFP0QQKhnGWc
L2GwE9x7n7EA0toLUtmz3RJcbVVgUK2b+pIfLfiogtfVXpvaSM+x8aASe5QJZ9AOIL/BoXU9Du52
k0poqecsSGwSrLrMXCNmqS0TBevNLFz9oQGlAviteFIYP5+xcd2rgtUdEe0wvoDwM/eFWWo3Q5P7
dnaWv0WBfyFj2e/9INaBU5pa3xO/bbceC9SIgPr7UQ3sSUdLBog8b/Aoq/nnTZJQjjYqw6tjY6qR
g5pQYeRm8LyWh5qAwsS3nBCjaeyRjsSyXo2oJ9h9VCbetxWdfDygE0du4+I9y2pjR2RDZbMQ1t/Y
zOaT4BY9FoUeQaLq8VakLMzZNPRBCypNDh9kCeEKE57gBXiK0JPcNRTxB1cYZN2A6zKCW+SIUg1y
Dv8Sn2f08w+jsB8WWfH3wPOnIDgNwkk0yKxdgMyL/Uova2xjZypxRCdemprFuVNYUh6t9oSs0jEh
99gfMEffmztoAaNiLV4gH0x1/hbMq7su79MMSRkna03a2EcVqe1EyjvGn3hGhAjBJcTlO/IaQOQb
KyszjrD5Uz5yXqtBrhOMo9EPdTOn6reodzK5tEkCPGshme6J5iSBgmXM/Tu1KhZyeFOiHxx+B9A7
6VwgKz6/SfaIBXl0Qlz0k9nStXEgwf4wXa9LfSaCfBNDNCiBl/JuW2xjlwZtGmryOIVJGh2qW4Jo
c4cxX6J6dTeF20A6uKXnRFRRouAMgtlu6kiMuk6WrjPUJV6ZntWn1W8qhZwBoqpUQahrabywn68z
4/VmTTBrxfkGyJ1Bv1pf95zy8QMeEwSaOluxUEVmOK8xxhkTP4hVoFRUVHavoHC4slvCjqykzXk+
oc/IxqnVDBa8kL/M3krNuqXgEyZBbUxW09NsbPHPQGkY9Ic7gq4vRNnd6ZLeKjPBIVKTc2NGIeJw
tmOOPCMBgMv0ianQrIcxBw2z3xpjZPCjkzmSJHQp3U+H64yfRIu8+tHQhdLxzZZvUGug3rvpEkAr
H/u+/LEnsWYEtiHh8wpL61xWtqCZpKaExbmEO+IRzfr2RSPkTHvJaIia9Gavx0x+5OKF4JV1DwtP
NWsz+HqAHuRQDLfASXhJ7pDWaSEnVSB9qfwC7mPmVHy5QvjZLTdE94YT5pQejPnsWxWRUJLdb2uY
wzkpt0GGE2v1t8g8c+PfkyQ9NTnx7eu6LYmQ0SijlBg8Dzq7RLcJ6apFFkSwSJA0uu5mdj6im2AU
wOMxtMuoNW5ekzS3QXa7fhacx8q32DU8nipbSxxLlsDQsCz3AWOOcdL3r5OCTViJCEk4yaBWGgqA
nlY+3r3S6CFkPhixmHRZb+zLJeD3hSJBo/WrRpr+6fphC433UTy3MGQ+XGtUduYKCirtn6K1dS4l
ubdN/nEwJOfE5jZbE4MHrQPwnjNuiDO3DFELHuimsGpOMJrNYETzR4PAa78lTvYiwgUssCMGmKQ+
nEZy/uyvL30ABGF8dErG6JAs8FhtC5GFFqLPw2I2smVKHfmTORGMquiUuZtXsZRwtFQIqpnrjl8p
Lw1WvdXa7iQ9uzp3aOI21izlzAa1QIokF84MmKP0VcAPfuKfj8Uyqoedy0I8Ct0ZnDFSmudNdkvr
7sFT0XxTdtHjLK5PpXS4WuRjKkmynyCdx1X96U4/Fb9Ql0AqSy/NcASUjz5ubnsMFTQddttbXHub
VMpzCdUA9Jg5d7hUU+WjczdXkD7Af04NuS2jrfkEzlvD61yhPk+793TE6m9/8t3h3CihmBp3r3od
4UIPUUunfZssBRMwCcm4OUYrbN/Vwtsu/KwGO+XUWpnfDCfShh5O1Sg1T4Zq3ZE4UPV/Ccz9SBFv
SvPaEjpgN0NutN6CRJSMxmH0J5WWKnPinIddA0vhVW+l4uIbpn66mMIR8O7Y6iqNpD5dp7HzBSiC
crCRNtkh5wPw/1aS71DyJz6zQ8akjHZdyYzXNmsmINdS0g3b90a4R7NqIzr4G6Polyci1Phc1Ex7
GWjwCJc6bccUTHXnrLykdMLMdUw4nGR/ci6x/Gp9uWx9tBQW1rWoJdGZbk5uiLntW01H9LwL63XS
ba7uMyeM7A/5h9UIX7oWBTgZHviHsISSiu08KAEeSUN+BE15fHe6OraMi34J0OPmPStXs9azd0aV
JkT0ovhm5dQSDbacpJTPbtxqiBIl1+sA0fexiGNBHYU4WL9WZpqznH9+n381BKYJC0S+y1vtwpTN
NbjXYj7797kMaCrKJlmnUenDXqKb8nTqcCw6AoK9p3huTxISVkyj/QHZBQ7Qr8yk7ByXV9nKZNTC
oPLQcN7suwBFAFQBxYoifgTzk/VH0s+wixoSX18TUnLnWdbaLcoD3lCG7cZ7fLIb7F+bSvESdwMu
fQ0/We/yCV/D1VrpbwSzKOvQQyO0ypzpv5Vmm5aYX4xl1jSqDavQJY+OuI6HywS2E0I4YaMVM+KG
M6sUsZ1/UYwvyQk5zvw5UNC3z/1MUoefbeO8iMEqPnBYwhZ4/p+u0XB5vC/mZjoO/a8xi57q+Ven
4mJofscdsEQU0zrgtR13ke3lYUmDR/GflrpAf48IuYUIV/CMlMG+qGlCG8f9dFjPeC+6MLk1PlTf
dBJQrBwkhPxFyVLNGvKF3Dza+PmpPJMNN6DQ1ivhE8/OuspeFg0oX8qlYDslzhbvEqKu7Bw1xEji
c2b9WaeTYZmygoSPRboZ4327x60GoHi7P+LK1e/ztH2lAO90k/qWRV7wLOnT7SppdjfSWf4JJ/Qi
SVRSVlcH6h1AUdiW24mS/zVu03E+YJTQAazQ98st5DUboAJbf63j/7pTpRYaITbIMszFCpObvVH+
9yxpUmsWFx1lBq1t4cxtUsbRRCppzNN8oxzJXT2W2+ION/ap1kuaeD1MTD1mrvfAT7rB8jZ/wiJq
VqqJHin+6VhyJzwLn+RC4da5UQwTcKwUoB0boWF2+QsStaSBigKBxynLkztJMcTLZeQOn2U0iNYx
HkQIfNZkuMJUXVFmSG44orrTv6M3xoI3Iat/pZP7EKmOL27pRWfBjZEaOLduwydGuSbYROWguDPJ
ep6+AvYZQHF/GgsfTnJKKu79iZPpIXPmFnSbO1kHm2cSKapm5mkVu7KUq5M8r7eRJXI+ypt6hBj8
97KzD9hrbe2kVY2vEistMYzNJ4w+uhPSCi+sRxcvw7Ll9k8XV30TxwnH0kOnMnBFpDrKzuJ1hk2/
g63vgKvCVupTcea/T2eRyYTPqgtHz7k9m2ER9StQeWkJAf33aOa/97oGuoEzSM85L/t4xVMCeL8s
M01yEX9CvWQ3Hgf/Wwe/RnPyGb56GCW+/b5Qg0NvneEA3ugGLnJsK4RneK8EWozydV18gjTgql9H
CI6Xb5r0ESMzzNBjZr4h5pgBx4Z5T4WkrbjBiM2m6juWqjvlV27y+tGDt/bkx+8a94Bh86Box4F6
PZIqVRBD6GSfJ3Dn34o8JkmHJM4OxS8iWjPcM3QBMvocteQ3pdmGBzOlf893ZvPlptxaBb4FXZJL
nfWmKeWOeu2YK2rcXDMrdlprrUTIyKI/M8iIY4wqeNpcrxTpxgst5IFSs4CmIvxv2mJN+jXyV02R
2PkViP3GAi0/TWQOs7nUwwIBST8fNjXTDmCvH/eESndNP1RiypdSkUGMal3U61bnYwuZZ5DUl/IJ
AjeqNJoxgz/WwuwbZFUAQbSmk8nqdJZoTxheNpxPBBbP+fdwb/r56+vNFEAFcNSNA+wOKmMzyRCk
THQRMICT7f1Sn5a48N96R/T0dgoNAxbgUkj+A1LFIq/bgk8jIgXayAsV3a9xjrLJOmO+0U+tNKoK
zdvvSKtFU/dKUK2vgCc8ke8gDUBX5O7DxaXL8kFvTtfE18y7PRGLSeA47+IZ4OBx0FGLk7o2hUh0
nE0KWol8Jm6qySYC8IBUVU5B+FLnjoo0nn792fCgY6exSypzsvevycT1lEtudFOfzHS+Ct2/fIkC
aJFS7/0QJCxTCFKZMBnd8DgpbXIkDYAZXl6gYrEptS1hM1PEz75ezlT5YAIrcwwyytLIeV1vq8sZ
vr8gBFJ2vww0zMFjqU4CI2zdHdG5px9SWC1qtiTU4q73KSV4JI4Uheh6/h1/XidIz6dduZXjy3K6
wIdO6a+7UYQzKEeRXvQyUevYrIsBOmK4o7H8t4WSEdJunBg/Mu6oYfyj4PtGwcB9Dos8KAlHRPt0
ILR6Cm3+YixHVEWR9FaOi1QrfA7dD7URrTtGNnXhAZvUCyZw7U8T811gp0+4FzezUDzUqp8Jyfoe
XzCm7hgHLc68ERNyBUPUWNj9DSCk9K2SCRIhSbu7ASAcfQObRfNwvxFSzIVEZ74cvoDnnQK20WGS
vzFnq62cW/LUzygPHDyhZ9qGP36hwSAIxaofnBF3pib+b4zv3MuN/uPPayAMgAnWYotgKk8zNJ84
lPWo80OJqNVTCfcZCrDvV616fxDcl/2Ob7xvgasvNj5AzFNK9YwMt5p1EjPZ9ag8BBGlCk4ouxo1
FDp+8ZUrkKqDkhylcv7RRixtdR5HRHqKLZjv43UDpIjNSkoDTc1lStM0ESHNb1XCvQJSHHDIYY1g
MK3pbeCYO3SVUSmZPj6CcHBLjvVkbtORlj5uEmWdiA3G8LoCVrsWZ5nYDGv9r6nD5lGOoup/yRQi
6VRyNyJ9053mXGnHA6XbPZ8xbM14Rq5IX0F2pbuE/zLKZRZKiPiN/zG/hJZoPgCG+i8gGazYNmsF
mG7IeKE8n6WfBCz+KXIvv6SG30/39aictphxZEZxTNfg5rPJ64T5w/pSyGqx2Ko8xgtXJWOl3Ppn
KPyQHCZpw7sOsp8y9e9sVn2mE4hC9Yne7rCwAT42iW8ZA6wwwqnfoV8J7GDgKcBQbbGM8laIUp/r
Vwx3UiCHOd2EnJDwMtvJfNGC2+1b5P40kySVbkQe50Z9trHMOcXiQca0xsDx+CfhoRbipUxJBtA9
Apw8Ol/Uv/rXjHGWGOTzpsmbDgS90gNg15yZu64Bpzr0+HeNz4MXCUOginRgbpZZfyOuFWyfpX5N
5UM/WTUIHZwURiPsRTPc9aPXczaWV76X7QT1WBktNOnWn3+Gzdl+ox+zjpCG4dnk/aMf4qC20KJ2
a4p39Huo73ulCI8QfmBlR6wTx7K76ZlSXG3osmDI2rISjSdk+tCVVdPJAt7jWu0XWEj7WgVlBscO
6iMYSuhPkTuuJLRHLdzoi8oZAWihuM1AKw7TVB2QM4qDBLHpHDrttQIRCUuYwjSP3QPZFoiCYmZx
LO6aDkwKedfqT91SIuiapFkjyeNMdrotGJujdaYx1ZeIMjb4fEHlGCH/wZ6eTbhByQiNTKoJNMfP
zZhBA2rUVh45QsJSRcGi6W6jSypauXNFGIMNiPAOsIBWmriQj1TCStLONYFHP+VSawRSJ47MY1Mm
qFgEg/9kd5+xK/fqA3y+xYXYkroogKd1qulNOofYdaWpGEB4bPKL1Ak2GiVllX1C7mE03RHtUpJZ
gEQNJsOhRM6jXbl8icht6kuOVKYdzUbc8U8O1Bx1sUapXX2Q86f5TksUQLV/lbDcq7+39UqTThAn
fwqNrDMYb4xEZJBBEUCGHF0KeOLlMrQiduQsXA1t7u4vkYnxptDllybadEeM+HmtyH8YyfnvpL63
ECezqOVWs3eKiQz+RrsUV0sk/It3bsnS2gGeE6lOJ331lbHIpeb00ICAOozF/3FJGe1AkDKK6dRn
3tNmBFpMWXPuspn+bwl1CANg+qpMAZoH5hl94e1rJanONVw5gvmMGPD9BZcdimc3mWJyZhspejRk
ubt/oAzKHmW4mAeGBydNd+T+KzzWuNOkO/EB24O90orG65Zy8pq1fsPj6sPdmwFa0bU+ATcE0eed
QmNE+uw/jNBXH8dnnOyP61KEoNRqD89hwbO2FKROh0gyKXclA6AHEgACFf8ttw3hhbZZtGp1juCh
SDDU/CkSGTOpOJWk71esc/7T8qROmyLmRdn6vD2805vZCQmvSVQFuQW3zETHZRNAJd2gnjVOuQyO
Ulm5hL2qBTe80efN/vnE3BRHTDyVRigZIvylHWZaRvZSzVaA6QZFxqxeFNW31kD1e6LLF8toCFkF
3AVFaoeY9dcg6Tmc43P6T95U8dLwP6uLfCX5JJkfZQr34XaLPBEypIONbteAkQtnp+0W9U/IfQ7R
w4DpppUY2aSgRWa1NF94lsyfBP+UOHr73DEtxiBxlxkbYwm5fiOLDJ4mQ432gn+paKYd5pHE+LJA
sYGMXM93wTxOoc2LZMI1z6Ralpuo2bSjg4+F2Qh/PE+o7mrlizDWhIecmkqLpa3boBjOGitrfT3+
K+PyrAuiK9yXdDmVXqgD3k6XY+yATvge9m+zYE+oQ4gCnc/RLvJ9/qEjfSW+DEikMcfasvuhY+1a
WcDwre9SHsm2qI9b/k8TIwjL2V/g0YDygNggoONUq5/9EEFFgfjdrHw1LwQIJQ99tLv+Z2MTBDyG
lT+KmWrngocwtI7YHZtR+2ygnUcpR8b5krT/YhwIdiwhHKzxwguwcQHq37Py3gYFom/qIgIrV8VC
QDRPF9j2TabPU1yF5JfyH4Qtd2Yfx7XRpaLVPBsDYzM1mgW0hJVJOu/5iWxdzvXPLIA65XfTEQwc
ArvklU4pcGpf3zZMmR66ZZlnvQRelqpGYmpZuvWL7GmSS7u71BGwpXoOOzTeoZc+ylGHT6+/DFlo
hyPOb9Fh98kbjl4ugloY6HTLN6F0QbYaCzBri7LWA3Ta94Ea/EcKlYKC3wPLUoDlCAj2IUySEOfM
X/EIDweHC6o2eS2k6EpVKs6fEbPvDDPBeb0RejC4AFmtpqEKaG1V+RdyHyhioeC/CjJnWGaQhKGJ
1yUC5J+IiKtFGG1GfuXmozqnhc+Fh41n3nDZSlNYC28/AtxX5FYAMAbJqfmL4SikUT4cfntEgI7T
Y0OiJetIm+UdCrONOavPS9ZZOZQgSw6q6SzPcnL8LODO6wgYiuMw9ukX4L+yqQNws376VF2TdwgT
1LzY77fwFw5FdSgBX8m/r0e1hL8IQmj95YTiaojwOFKVt+LJKkBTlJKMqSEjJZaU1eDkRQSs/YAo
C8m0gdS5VyYzSDm80DOY1ey5pE9hZsOe6dlqlhgqifk0Yfv6YUaSPe92w9XoVQlORXkQSDLY+TCO
iqB5nr01SJJboXKpHvIjM3nXj2lU/SnnNP4eWNpcmJL1bRbFC6N1Lk+yfdePyWUZ7vH0H5e0qCX9
+3h8/H+c2hGAS18DCdLGJLcnr3xvws+BUkmHnWQmHFhxETTQnGdV60IyJjuUtWE22JUs0qFoGqUa
z+oEGI7P5yKKtY8V6uHGeVOkkzcwji+4bE3oaJDCHpEilDR9eTctz02t/IXy6h7KEcyklE0vbif7
htZAO6M6OLGAEAMb4Qq11B3/AN8gbqDOmgOg0wjm/gjgMb7vzj7ikiL0y8mNZmvmAoLDS84f4uCM
i5U97W37HlC1GkOObpT0GR5pm0vxyoiYx8BGVD0vfWUxbja9mi1Ji2rwsJy0H6QCX9eEPtntyjOm
FCdS5wSd9wHdwl8IR1RQYVNKmd5CGItWAnOnhA5Y14atlaQkyzc9a8FX7xk/EBylORGovgEehwuP
2xZp7XNR1ISn/e1SpwlSi0ru1c/lXNxqiWRkhFIB3haqn35ZAqzKAqd8D6/B0ZCLQF6Kl0MZlGgN
fWFstdect3++2oosZ6AHEoQrb4NEEwEzj06SDQ2DMgDFt9NJb1RRqq5qS5hswOljN6L7NZlRf+/k
uAhQgI3cZ4A93cNp/hebuoYAvRaOBK5v1id79Mm1yDjj0sdBCxOYNYziQnWUc0cwDz1iCvmRL97M
m963adtOQCOwV5vbpvEhG2PThbn5Vr5wNnMnEdl5MZ9o2b+loqVve4saM9OFJLGMQMvA/6RoFqGI
B5BDvrKhjxO+7b0Tg9h9tokXTL0UKpLeg3sGG6rd0tBtJWtv0cqZ+30QAVmvlAkC+RVInYRThVSZ
M7l/oWwoEE6N4izFasKkO73+ZvMWNh073XTK1AkTrfen3N4ZbAJOwrKBWpBcveAg6LLDlr8qvgfY
pH+MuUamYt9egfveu4IF66TOalnW9rScF3rsZr6Vf0HEA2tHIp2UFD9JF+6YguSeEEir3XzEqTyN
k0VEpd+Jctew3S+NF3mkAMdqZAFzjXlXXeRDyqfbCoJJY3F51ZNy3XpFXx5yyDmBiq2ALXX7uKDD
u8RyEQsBgsEE5nJKXKy2yV8jnoQBOoojtmOGSau73Ux0XWenvPOOzz9aehXGj0tjElt70+UcbvPG
uZW3vAFcSLzZEyu70pBKqTGzpCxwHVfgWH1GIbF7JGN+ka/F9yuL7PicZotoVfe5f6YPt2PaD/AR
7p6ddgbOf0TzMBa3hDkrw1vB0gmNyQci6s9E9LbSlmMLvAzmAHB9yp37/AUNmudoEblKNJ8cGsDX
MVztnwb9iOfku0f53+MXO0NV6ipA9YYJLgaitzhum8WdkeZVTOY+jFENCnNIqLMH7brEF2b3e5/P
GiR7cac0lH5lg+pavwHT2+YcNdMGMYTIglAVwcllysK8X1KELBcasPR7qwQClzLzJaUQMcLpBbLt
VUGn/UF6t1NQGsX9n6SP3StFZNODxRE0jGie2hrQm/UEn66LKxEdvBe5/AsEGLXbAw29pUfqJ5M/
PHNXGt6ajkikxy2WCdws30ZVl3GQBcgUGO8rvBYaeXxVRCpWu6XyJxAhYLhsiCfWjd4HyFledzIP
8laCedenVxilnWFJ3Y5iAc9SjDlWScOdeA4JxvQes9ISKnN09CEE/tMj4WzpzAnu2pdGpFHSyA1/
YRDkchjpBeFFwDo9AuZbUFnUInN5mFBWQ/regBEZP6YUFc7+Yb4b++CQwjPJJzKQ4JHtiyEyqNuy
7pC4abFU9VHXUE2Y+Y8ELrZe5XaLnNfN0efPBliKoQqgeuMdgr8GLJSeAMEzB4ZX2BmfgFcDKz3J
jnmlCrzP7WhiCzasgr7dCmgMQiGp+mogikq6ZQe7adi3ciR4G06D8FEtjxLIcMk6+/DVpidcxxVJ
2InxabcPVGGkY5n8vBFpxcHkcUco+CysWQYR6C7oDYZEG+eKbfyGdYZvMQVaaQBtFiIFUEyKDF2c
6nQs/hEecnaY4TcybnuFrZFHw/nRVC8VRbFR23sWlffqRJOhi4JLNpvgEj+oDvGZ+GnL3iIraFHG
OeseWXIQiAyDtAlXSOmzIJ/0M2nLjchfceVIZOBTUxYVFbTDtUUDO6u3K13PjR93q1Pl+AqN3n/6
52lkSHeyg/bAsON37x+JdTdbGv44uNo1S8/0w30Nqhd/6HJnu+763CdtuOx+VXc60DGCL2PshlnM
AoIM3psO0BFwLdMZfEe3feqwHkyx9jzSc9cnfju29PBi5GS83ZWkUPSXwege9LJpx6emBUJ9xLDx
cOyt8p+5UBrcFuT8lU5UqzVsEsDLy5tvCZiphZBE1Yb8/EDU0PAnrp9As+DKOCy1bjKlW7afdUAV
s3J4nKp8UtEMRYHQ5o5B0PXERz13Ht88PxwfLn9GHFFJhzhfEHZVy5+UKJUIa1bIIT+KNmKKijMq
Dn1FWfzgIrz2YGG8cjZFxSYU2r3ZX6qrZrjLzV5xDmsvUpfE3sWkbLUEkTfg1u4lEJT2Zha2cIVN
CfiTi9AtDUL4Y4NOCeFAxh3upQsj9k0adh0JY3XSuzdbS0KtIO3wsRhAjb82eOqVtpm4MhOkmIwf
vunkR7VGYemOhwsVqDAMuLqyGKH1XYX84ngxn2hAqqCrEhN26aaV2lyrdiqsyEeNTxkckHDCUS8a
zxQUaC8T7s0fOEACPYSyy01qY+t6gar02+VY9v5RBcgpv5jFErk7ZBit8ec2tXQ3g2f4jCT6SwWe
f1Unn45Li+9TH68gC9O5B7NJUh7Tk9JsaoWoYbx3MI/6yjcqQs+T0FqNFL5/ZGaps2kNG05vub9Y
ySM9AmFXEkMdEAlPPpbsQN1/fUknWgeVW5W4TNPxK3Vl03ft8An4HTJkU0U4uhLLe9GvIyfIEqkr
RPD7mEtMNrUO+xgedegIdVdzKErPdtcaMMr3Oitg9Txg8yShOQbctkrhCG5myLuE/IUUzW5IIhcf
r+PIxRb6q8q0Plb8gBzOOE7Bk/AqRw38sfyHuTIwOvTsY/xeL2JezXGadaHuQpC8ycHfmKl/Fgo3
rU+9OCPRyWZJFtHQUJ0TSGj6BovrTHRcUutHZKSmn0kaaVfLE/U7JqEpJRJHmD7HIRTrLHcttr2K
HIlA8iO5SSzY55sV5AVFn7ERTaX5BseRM4lVMfoiN/gAS2HDhpzL8/hfQg34CwUVKpCmMff5DlVb
ActWrk9oeB1VwWvgvEqEoipzYwqguBtQc7Cb38i3o3NQMDNtioUf4XK0EIZBk0192ZddwM9l35OU
MoCDtH3F+3SCtFTFwtfkiq6aGa0w0P7RuLiZBjLpGIFR0thBZ0grTFR8QHTobGpTmcouSqOhQ61N
myymgxfAaUnDUy4fpN0+b1kxOFLESdd1s0FryRjt0M2x3iMCOSi9B38GcHdu1w+VHcgb4uEd7DSU
+Fsp+c48b6mhyCMYZ4/OljpZ+CiWrl3NbeW8nIaD498AsywLOG4ISBfPB6V8wQGMMd1nCIj4/5sU
vsRF0VIgLNk5xG90RSDgnUZjngcUGS31XZMOmNNXImiyTzdsDYDbuwY9zVd2Xv3ebbo6gjHV+tBs
3MTUWa3X2rlC4g8a2B/B//mZ9YnQSdjb+TioyHzXJFUI86N5kaciH7k/3FZqzX4nH5ZDiURy+e6P
tFA+4xsHyMqw309lTtAjSs6LvB5fpdkjekX39qkoHynLtTx374GxRzw5ilO2SgF9kFq0QgsIE7Y/
OIaOIpkf2F9qS4MSD5H3TP9Lts4T23Q8VFHeLHc+SkGzz8MJKgJ+r02CBeNHKKKpPhAEcZE3SwJS
LEvZYXc9C1lpU+zsswx8zCj8eQENc1in5oRAmPoqIoXJGEvF5n+mvxWvR3GgwFrw26gI9ZX6AQ9y
EOaTGkOlMX3nZ3XgRrKi6Z893zaepRV+Bhmk+RBG8HGV5MaxUfwjllPdf0aaLhiLKOF1DaKrp0SP
HW4q6UkgnaYSDx1Ej2z/Fn9ZTthfb0u2TX5pGT+HUFs8t7PVW/MvIVoDa+jg/yG747vtVO1GsIUl
7nZ5zotGELrqX+zwSBQ0oPPVGD6sN3oNnVlIFoYfjqr9WAoyL6yZpCWrOjjRDdxA6MfcrDGxj82k
h+p9lu/IOqD9KaswkLWidEuXaC8Pk5AuWeyyTe3QnN/TE72KutoqyTCnExNs5j4PbpXrD2hBo4Td
yIKWN6hIWUf3n2/+hQ0sAzCF3XNQK0unjiLre2/rTsakow+5gQZEhfpCYDC3Z4Vp76WOrsBh1pRZ
u5dip2Tl39pHxfUDCznNPBWNJuuu8bRu/nmtia+zzvde5Br0ATGUL5CTO8EDUefWHmpAzoFZmmgQ
AMfzmW44nNBJLf/xKTlcRVP75qUUjEKPkQW9S3iqmy5maahkjnXW4Vn9JKhSzMxFwxOfyOdRANTI
fpORQrsU6onsZ7VidM/b51C0z0N1KABEe0vaEhRSgdLyfGj6XaN5fiZcGnSyuR0McNdtsSxXya7P
cZbSZ2ou46z2Km6EPPB43sNUsi5jNZEG3dIDHFZugpB2tI2L5qfawjdglPixLkJOCcNyFYxqKwja
VLGeZqEK8h6FjfMc80ZKfhhRAzlpw3qYlz8tU+NI+0cC2CQ9VDvTg4kZQjV0U8Jgfo+MXQMvw9XS
a6tkV08OCph+ETiK1x+JpB+v/5HalDxPhSzpbTVvBSHv8KzbGT3RmFhmJRWvYpVuoro7j5hYjNKl
mUhhmK8kVioLrCAeCHXibEsLfBvKbu0mjit7i3YoXiwYqJJgXW0M/k+L1zQpmUjUR86wWogBVTy2
PRKlF3n/3nxnKSEni89iJBZvinf0VjoCnnnEDGflP+JttG2fuxjTOTOJJP4H6lxwnZpiu93VZUtP
yhhzk/qMHZ2FCqR1+sTepb3ES4U2Lx/u1UOeI6TQXFg+XGKXEEx/+ZK5KaXnp10RGWl8U4L/iZ1f
Owo5FutNAliTHktG/wM9eAHPWO/Hy1cBbAklL61gLLbzwuFYdFmZBuA/LXlvwwphzGrsRLfj5Far
vYHa/mTLl8Uif8iU78Mive8VF/RKOiZ2c3MzbWWQKM/CI2qBNd3RSxKAfoRbECW6iZcP9MmHiSly
Ya27wc4vKmTXQA8cMlkNCZA5959O5QUsk+bdWJpr9jDAiHe4Qtr1E+6TWV+FaCG/Op14TzJz6ukI
NTdXyYIUtLuV+ufNMOgvU4i4SLjf0VXPb+lzRDe9bbzQ7MDZGaofH4sfvaj/6lKXKcgHv8elmuBi
omcwxR365pG7JzsrlE209Tl9CL0tDBLqoO/o24uh+kVeojBnXUWJ1WS3DNMMLyS9+XQ972uDy6Y9
EWkZN9VEUa1d0NkFzE/Oyd4aiF9cqb8FAcnK39iRN3Y3hwfGwMo7OCiCYXqxiTQOq2S+bNgxgiG2
lkaaTSXp28uWPCEoKlgCaBD0dJWKeNkCEAn//7PoIdAlVZKOPln5wrqbFYcOjzLCOiC8/Dog0Rgh
KhilXArpw2g+7wy/zSayIA9QNG/u4N3YPV2nn8fPIjqTQdDQVLHOgHu7MwAg+jKa331YlSm9+YeK
ZGe6HJelwefn1Xr1taoY1k9aBe9GQhpUPDP7Ndxc7an2OLd2VL5qehV/ukZmSIJ1DjMBb9+DU4X0
Jn9Jkwo/oH+QDhRF1/o4jpp/OcLX7w355qTEDGL/b725D1z2eFpGCBR+va5nEGK+/+pIaLvHyA50
wZ0Zh/Jlh/iAs6+lx0e+6DQ6rBuIIN/7JaWsG7EskLSKwQppNWb5Ty6aRKbfDowDO4shqtUMKUtR
1YFoQu1Cg5ZfonecRC6njd8qkRj+CAltYW8wiNrR6D/AB3rhH/d1HoXL/I06AN8taK3BDCKf7Wc8
7hI0sUZrAQrPN8nYAFf6wBTOVPyYe2QFm66FHp9UBEhfjDZBr/Lt714A/KyKW77kI8VGmBmHvRbq
tpgmRlniWKeXnG0N5s/EuGw7zYJuWoq3c0ehLxVhn2EqRXJIM2d8tykIFj9SzT4/BPOkup9k1Ekl
w0DbRNEdbUnIT52mRrHlMMDB4d9W0NOs+mLqcqDapjUuEnYSKBPLZvqiBKoD8yPaeG40v07lqiJT
RqGHFgq+bt1pQwRdWLGoobCTIsTcXTdxYgZbqQca3JZAM7wArMD3BpYOVm+aeyINWR8PBP/QcNQL
a6RAR6a2pAMYOnzU1GiU7XOEIb5qCHzr0V7bbCgxs1QSS97SUGlY4XkRqGisz4SS7JcmhPx8zyRu
Awvc7HhGw8EkxZHjMyJmzulzurAL33M3gAWUdBBn20X49CB7UqgF7lDF8L3JADbIhZl914lY8ZSX
jV4vFJMcgyjiDDZE2T5nOgEr48QB6lmE2Pw+GM0j/Vz56fjn5IfyrJJydOGwmsUNQ53+Pv0m7AXD
24FBTNsVfqSfx/pn1YsS2fq1zL9WFwh1/2UKAJFtFCTJes/err37AyuDnGmlzQItMkHWt0dm5bAn
seXnvgaynD4ktIQqaUCqtxKM5/y1GBN3KW7Q+VRWB/7VhevunfFHhWrP3+nAi1gYKPUdU6Qw6wWO
C91UxnZssFoxz4Araezv1aoAGArPchZguNgKbiJ7ftL9CjsieSAocXs9QLvyPEl1HKDYPlVqGTWP
//hF+k7O/7NJbg7APYgUi912s5nzZv9wfm6rEip8VuZt2u4WdjJxt9o31UjKgoe5RY/aoI/PF3er
5zJgxJ4gGG+3s99vqD3CKGgcFhD6UsL+Ogvyg+UcZfjSTO8Jxk4of0OxoKW+2QpV/KvyLGjzcrQ5
mTmOasdjaTqpDyUVHW4NKtuq+djJo3yOHJkCb2Qi18HUGfd3tm1av1im/J3sIdz4CdM1qxRbQ+tZ
gBZzaSHkJum5igEkrR0r4KwFujCJ62Z0U+BANVlUkjgAYTS0uIKyQdsNIH+lvDY2IGDgzhH6hiq2
SOmoxIwumesW6k15bLSUVZWrp4g0slJ74HO8GoTfKy5SVGRikJxqvjk3c/8xY9q6/KlT3Wuw7noD
/8PSRkGsDXG3wVXYmNSHtxkZHMRUl5G/6awJ+nPHGEprLskkKFlrw1IjdVzsK/JuMVJMW9+fIBNj
sKDuO5LJOjTEbLeBKbWNnbFFtufxDCfqwVIAulWvEc3WEqDwTcIeBQvgTXOVXWHoe4li09AaaHMm
fZylwfN0p7gDmSdZGAFWX6fQmlKok0V+zlP2woZ49ayhISr9om7CDvH92KL++7sSK9WbuFOmWsnx
hRSbqoCWo+YKAprqlsgpvlpDdzetfu/NdLoLYbdvHD7ytyIBXCDX/ECR3XueEpAqhArnh0esVZF3
Jp+1VGwv+Gus1nT5VVX9/hgQCTuxMow0Hk+TsygKBQ4zlQcXPh/0+MZD1AsX9xdmeNkXUy9jyDnx
Dvf9Q0kD5hGw1puVi39Xl5RVIL7KPGCFSKl7q4xnKiBwix9lPRWeC6STnapXkesf6KFjVXoZYC8C
iNxl4TDPA6GzPJgIfqYniXVV+v7xoPxcH3DJm+CFDxYmiCgJqEb/i/vV5OrfygZhBIg/RmahVZb+
lf7LaiWjbb005SYLWA9EI3ZuQnYBJMi1IxxB1MOnvlwEcqY91PcOssn2V+vvXHBU5i9tf3CUIP2g
i7bF4y/oGo8zBIb35fTnPNNqykVdVJgOXW9nk3lp3NHtiF3295MKfKw8eOFSclodkgnOLcju4ViX
g5FLp+JxlBRwBAlMiNQ2dip6Ptc7NI4w8nP/vk+DWyGQie4J4oKCFksB2c/7wjKJO6reF7tSjCBK
lHDXVvrfwz6oRUIJtFeZtKD3JdHSc81Q1c2azn6TutL+zYQWQlWMbvG9Z9/Xo4ffaq0S599jNA8Y
3eQ6RiSHdslN/GIYnJXBGQmQCXOp3ZM+/ppVVaA8mAOFwdHiB2j8vmobrUgfeBLQRErmAKd8zdPC
ijfbLs1YF3EuQWcVsu4kOQuT9ClM+HD3K7kKcPd2xW1hUwm4owBctkAt/vCP9WHr5+PBQvl5xY7U
2SmpH34ocmi8EIgaxbvchTo7U5p8I8b9BvCyQI4BvYAz9NrTma6wmUXqCSTwNoIainkxloCcEKbH
GbM95ii94eBioDREJ2B31mwUrFFyNCozic/sVj+HotZCIyIde0bgVL3bZUUs2/tgUi2THLpvfHqi
eeDD1SWAJjhSS95B69NbBvEY/MfCFYh8LkR/zR+iwAJkkTqRG87cWTz9ZlbbVcAVCdT3SK0n9oXp
Yw97msNKK3kPRVhBNw7ToXHt7T/Gk4LR4haowLC+9pAdO9d/NyxA/d0net22zjHV0+GlzHHkUMri
ZtKHHGzXD1dPg1CqjKPdrlzKjf/CgmnJuBOR6Rxc4SnH6MN91CSFtWFO+fZEKpMpR+KiUP21FBHp
z8S+P1ajznX2+BKF3gGPfbeSYvl/idf7WnK9OiA9bJYP4yyM2idpQHCllFGNWv9Do4Q2z/nu6ZsG
lmtMZwsI5f4Kfab1Sj4zpJ8dywYGmCiWAzJ/Hybbu9jCvvG80GUg8MIz1KVGoOnFm/M3kU0R1A8q
HYhJdrWgDPIIk0W5gaGgJu29XopscLOHyVFB5uriiqUyiW15v7DCflxPS6vkean/pqnDnuqsetOe
Pr4KGREypmkINigPdbfDTFbyqgwBaf/vMcGBIdvNgzE2Xf7bHx0LgB6Qsw2fG7B9XmePEWc2IXD7
TPc7B9zdU4gASPW2jSJ+aTwiYhw5GnV/z+8Bhi58ypkeLotdTE2O6gCe7GWuSxUVt/66/tcOj9O+
VtFbwQCYVvmkpoW1tSp0Lheg6z6M/tFviCJyPfzzemQtKzuZ/Iz5NAsSDN85aMme6QIUgzLMOZls
2/KPclR0b40ePLo2X2ftEfNOq6nIiKKKRdgFgl0dRXkcgdCWJHMGpCsNcNmwL2caqO1q4qRAQ0kE
BgvDaPEGZIyJ18FDLu5qsdKWd0u9zmEHm8/t63oR2wLgLHg0fx2prbM1sRXcb4b1Wul7ZwsxREhS
x8kBzhwKY4Sg5SAA9Mggzj1cPAMQrk+joZcLmrgre6VGNRwxmR8AzjYwptMqJnK6D15rvjkOvK18
OkAap8/Vhr/KZg2cNRURX6Sbp12pduwZrHD370Eu7tfbgLgfSoq1DY07uR8IL6XsZR7fqH0m4ZGV
J8TQTRnlJh9rzjceL/HMJmQRoeLttoppfu28wHC4iu8DDSKO9l5YNU9BThfq36JucejAwxSdCoFO
spnjq4urFmj2YXdHs1VQwuKum4T1MLlk0Frn7jZk3QFOqi6xLnSwPpVZdCe7CZ7D1TewlzhbM1P7
cP8Tpu1JwaYjZTcceifLW/SGseTSlkh4cRUzsjJUwiSETdkhuGsjT9r5a417BiZCI4jzSamO0l9B
BJZ8GMGrTP5GMtZiWBJTRfSHf15yqKGuXieFGWTvVTLWDhw5z6doNRiLUTaA2hpcxuHoluDgWBzR
ntUNAmb4D+EuVa45Y2kIDkdrVUu6jRzxDJbIuqgNB7CytK1xmQ/94Pk25soatK7Tqxz8AxbAKLgC
iXrS2hAbT6qqfzDrpVAIoIa4BEAc2OKO+blBqSpAiQiwwmOoM44KuEOcnQrJ5YaOKQleam+KDyTk
1yxmrKs8U0EI5HaIGMD/zyimXe/VrNBwQYiGXSvLb9FqpiIwXBINAiGolXQx9b97Wals7Tks3kiY
egFYw9mBzI5gZuyMl/MhNtcunXJuhUkzWjW2V6e4kMIhlk676m0BCbRhFIcjXCVyUWNil02jG9Uw
UE4C0Vqa8F/B8FyAg53AmrTgZWatSgWhR26M1aMLN9j0P0BDRyyY/FOtSnO4C/wxWf+9uBovq+nH
+2zjDYTuHxdWwh7yP2uWarC2eru6jLaQRkjMbFinFodIs/f3+FXU52FspKcmvdZBfw6makGrimxZ
0uQcj1WQKYs6+TF0UfsjoB/nIkP/gSizBd+GTS/q0pDP0ogtfuLwDTMIn2c+dXzY+qPs4zcJmKYE
rMVo+Zk81jVHYArAtlJcIozfZZQNhyWEYzSr3dD2zT7jS9FeTO3ABui3HUrNNCGK/Yr0EDQ4P4+o
nvBvgXUAqYG5Zd6P2DPQWwKI3eSAFjihXDR7PGn/5dI2d6ZbL9b8TTNDcoUWLUZwULciB+2dOfuI
9QHvvn50jPlOHscCuAQ4q/aR/aW4U1mIABRtgljtzDM8eF/e2DV9xEjydl4ZkkV1BprNkFgZRbbP
w5g8owOE86tn3A+FLk2GLjoUtpqxI9dXf8S2/Oooo3QjUcJO99L9YDhyq8drJjoTuMspw3xCiuXw
PsN9yjfvM+z9JZoyztljvqNqcQZPDc9nXokyKZm+XyXKFsCWbL2ZQGJKj2QP51wecK+QzSqiRUjm
+Ss0ZSGliOwNHEu/s541wIPbsRoQZsfTP/YmPeprEXLm/WUas86bGfiDlE1iqIURR/oaqm4qw3kR
XUVP5elHbd5vdivW7BW/XxEX19/8d/C4gbZvgbzMIrLUtrfVu3D87I/netlegX9P6cbULT54O6S2
1OnEjAX5IxzPUo/i8ztJ0HN3ds6ENTE2SLxUouPr5y2npp+7W+ocPCWjnJdUioB2hEsueZqIxa6W
9zIu1sVNyf4qLOl+RhwgO0WxHthdTXXFuafQDE5eBJNDBnhbMBEdiB6t5emz/O6gHmPKzj0qQvGw
3lFxn/DODKHaFIUB1GnkZ+KRswvnP6sOaYmPkESmBcMY5V91+YYHKTrYvtslQ4Xa2NOltEpkNYXa
QVBNmgpH5ZGDHRMmN7rIzABdzHrm4bfoJC29zqKx9xZRJqqU47jHJl2+qfyopevv2Hwy1+3DZAOu
RMNupGXPTiBMz5/EjJWPWQL4RqQYnxjWDBTcilmWrJvV3VDnOlBN2M4fQfkTxkDav4zwZIG55oMc
+EytAKCnnMBgV6S3Hyc8HeTkfh56JagiYl8dOeUsML7iSH84JB5enl5nbi9uU8mBkE6bz7AqZPhf
SGnC4TGT31yMMZpruVzZDrnZwhjfs9yZgIP3SHFkibW+8K3yxqhfxKehu4cqTmvIIwSTvBfDE9KI
tD7WMbuISRtZwAd5Zl7eFIk4Y8GWVx/DrK144E6zQUnLvGgejjwF21p8UdLPydevQFVUUTWaz8dF
dUjJO5Q5scDqYDgL1FtFR+B2taUHVWmR7Uz72QUU6QqOrlRXgVVMSr9dO4+1ULoiR1qnKa4TOzLT
Lk0jYlBPthtE21j73DlvkqiwqkHFbKZoWzVTgGnolHsUmtcE1APr+ny8h2XvNg5sbF3SN8J69LXP
0eugD4rtXpT5oX+GDLtBzlLVGJEfMBTeULvaIy/nLAeYgdApVBwqhGWhUskptXPE50IH2yJ+IFU/
6ziBk9oWNAPFV9QZkNfgYmhEgyPLou8GMo0KGGSYY0VsknigNsfT9kpFO/IgNlXai6DnGdKUOdKy
OFFDdpC8R2tbXewOJJZLTfxH0O6TN6t6P1pmtDhkRPpfVNw+ntiHupU8OrrbjEUeEqT38iKKNSSg
IOcvQWzfXDF97az12abGz/WOOXBl78+R46j/hULGbQt+FHnr76pR0PZbIeK3vzg3IjHoVxrQDcAu
k9XYVuKGkw2eQa8WqLjH4V9jPHgzYg2sPPiNusG3rMcjVxbPnKh/BOgB6wazfKC+xp3F74so/4/V
EkUvzC/ACgLCRf5KSvN5padtHT8YR6XV5uJBAHQu1w+GylIR2dAYmv5QRrqQ6Mi+ZtB9oMgKnZ79
Y25lPm+Jqgw5bTqyEmbVkdXQLPW/0k31S90GjxaGiRlBADvTyYtbfu30iugUaH1PejUS2kl2JLNe
T86qguhDfaatJqlAIaXvYfjnSJTvXQ4dqCiMbBKiLaSCZRwMmDVILmfMwXeyC8VLZum16k8SCaaT
9zRen2N/MXYg85JMgeUUeJCeIKNnM4OCQ5rN2R4YcdyUxLXmQmWVnKvlcwGIeBbcvqRjRRHcswG8
u4IRgLwj1ptqZk240iOI9lYllErjEL24EipdSvaN1bdKrFzN96bqoBNFQIUD7KLrgLYDbB2Ae8Tg
2QNgipY8VH/poIU6r3oiUk32FSeIatbUJOWREsLNeoS/HT3DSjF9KcdM3mngFL1KtJjcK5ZLLe8I
jrxFz1sfd75/1PFDofwGYYn5OqF/NGWTO4s2gcejK/M3Fr6wZRAwfd3zA9y6inAiNgP5kCFMoyss
8vTDnJhEg7HfwXos1Akq8miMBaCQjo98AG5W13Qf4dcwDWH0RHpUylw3lrVfClDmgQf/dniPUgVp
czj8A2JTBwEybIinylwH98QlTzNTi5usX+Ynk0FgW0UCo73ELNEm93a8TJ9ZHgR2aFpYYH0EZkuw
IUY/xPEXcrVhc4iCQEZOR2W0WBvkSdiqO4RnyqpdE6QbuHax0I5ZQWHTFId0nGmD1xppuOfIw1f4
Sv05zR/Z355tJ4atFzlkPBKhpD1wkmfJ2toHyF3BOtTtB170F/z+ElbiZvDqJRA2ehoYkkDFWL6U
/6spSj4vrEpoQOpFp+BbvstQqAQPdGgE5myj5LALPGa/s/R6odrbEZYM9ZpMHrJH91HI3GClWTZr
xByIvyK+A1mgmomFmu2bhsQF4YVOitRob75Hj4WOb2b8p7SKKCucKYJpC6aBbalEas78dyzNWtzJ
xZIVu9IaOvlazp6GsMTOoJpD4mmYVc/DhAud6Z59Y/76zLSOsYtneVAEUy7SFiGu5Ibjs9ZR8IuP
srBZr0zVTHuDAfmofDHdxOl8YSRv7DxS6gjUIRIXMI9G2uE5QZj64okLqzdRWz/P3+tO6gEVerUU
VriHlI1Km6+b/Zc6/9US5LwJx/N43ylNaOlnL6e+1ZAhdn+Q/DIsbjgwgTjuqxi16VcXh4jdcxJv
iugWvFH5P1hRyFzlGgpKuGZduNJqckXsFADgSi9QO0xPRBTXS2KHF6tuYvGHbL1aWr5mB4Zay7hc
QjUgPUk2AzJt5EGbcHXe5a7iGqTd8P+2JEGEM1oOl54t7xcPR5ciN7Dj0InvMJE4x3wonxsUcCxW
5i/VcKKo0J8OQhNS7ooEmCXECM1Ti+lWrl1oyRNrk6NtuzPhEmfy7yKKmirmA8lmbINq0WW1QdrV
YTGZJLxk61zrolmzj/d098cD5IwBjzHdik2/H1uQj+gE7dP0N1WhB66yYFlixWcvhKnvrc6RZXHT
C+3EdXXhFj21yL8EEcg2VEfbl9Wlyd+McEQudctX3i8b0uVOpB7Ab7v+YGt9kW1Eqf9HUYvgwi4E
+jmF7tYUBn1YNMAxSw9LoFiZz9xrAV1PiPdHhV3fqIdiXeReHNdXtgcgRGZX1Y54dq8tXSPolbAj
DZDnoDsMsmHUeQvy4Q0RXSCIqbErUFJumPd2TCj3FniDQ+MIOPx/Of/xp+Mn8AynOIKDGE2zYbWz
ch0bhBJ5vBZSqMoHN+8cpTrRj+I2p1eQOued1ClcJqV/qIBzTO9uG8JjR111b0R++ZtyzqG2lTkt
KpwBKQePgm3YBvLjow5tD6fP5MfNLQSHJbuOeJ+ICx5FfRwXltdp+t5K8YWIgMSboFPHVmOGKoxq
mD/E7+vC1BvyYff7lbjBsr3/e+T7yBvLrhUAAVzplaL3+/ueJwdbd0XCVurN+bvEfI6dfBNKFMdq
GHxASmOvJluSIB8lz5DjXdaI7RJ+NlcTsSeqvTAjf3gU8pIkJSsV+jClyJi0lM7cAZn3KIRnhM4F
jOtiu1YyEoGIYH7lvkFrxwC/oy+ZiYsIb4iHQkl5vNwJtrYtbUldqZG3tKlCDmV2ULWNueIo0Lfr
Tp/Q3Gd9Hv/uKXdQVIYtSRKWssMZqI7+G0bHOH4hen7tApSCeOJr+xgVUO8ew31XHi9FaQrUYdzE
WfrBtsuvWb9XKoAnyFpFyE1JO/cYwNLxJu8TXT8z7OjX3z/QM4Ik4L7rNAUaPy8PGFV1WB2Hv47s
od4dcd63IdROFC+SqsGoizJcLbKC9HQPxqSb2v1tMS43goCQ0gGhHUZOJ2CundK2I/jsTZISsqiv
V52nvr4IWURvSHHJmJrIpy7piHJ6dFwr/UEJYWmRsgwC8bBYD6ipJd4kBM2TTuXyw6raXx1Hz2T2
6l2i7cY88GnqQp9m/r9S1I73o9uX2n7w1B7gOzqP1+DS6Kiqutrmbx0bhh2XSO+7K4upQam2l6s6
j+f260DPHvLU+krsoGC+vzuC0lW85TgpsQz2KmyZ8+/k5NLE0gG1VoFfQwPhoMEk+b6mPaI0V68t
qP/vSNjqTLbRCzsZjtEQUmPXK00oXnMtmcC+3rF3kaU2BV6B6d4QqL/so9ph8Rtek30KLoUhAjws
fRiaoowiiL2W4lRoCRGX5ZZGbpPAjO6Ng5+/HuZigLUbOBiP9IiqkNp2Z2BwrqPBM4g/Q3DJlUhQ
NQyuZ63FuyAdsmTqxv+NUErz1fqt9/Ds+KKtCABBuBqQ+DTMrUsXN1nenAYbQyi4IUTG50CfMJBp
GygOit9UzcS9bUvM2TxL0asLeXi31uGMJTbAQanvvEhrNBtamqJziE7oL4nE++M/W7bg823ijY6V
vIN0fBjUjOQXhMlb6KYb9SMG1n4EUri2SN0gMj5MwlVjlKXP3egJ/Bkn6L5mmAQa82Q0UfmXA0DY
Cij02gs8g5suhXRPJHBOuQvcTSxRfMm+XsHar8PhBxZ/LgclBx482uIKojOW2nBs+tWKC+pbDkdQ
Qk7xkdCGbXbIfqXbeXNE0aFvCMLEpTAJBXEsG3rzg8hgtlnirBt6NMcB34a0kcpPFlqCCn3KUir8
CZ9/yFU9oKhtRAwfEJ2OhqGqeoUKw0Q8tPvaZJTphdkGzkL1yWY9h3dtF+Rds1ZlpKMA4+8/eBV7
hMSJ1+yFXqp1RgY/3MsVv2IkmSf3G/F6vsgCo9RHFaCZkBPNrSPTKfiKB4uzAIivq74NMJ9rRYZc
9HYfwFdWvB3awQCrbJbGLHwldnNrW8fXXxxuZcOGKCMPML7Cp4Xdq0aInBJ7qGOo62pTcnTKdx0q
ABBPugmUrEJqTyiEZKtlueNZ399qyATtYzfLCz8AMl1FCJHWWdMxYYwuzeGI/ich8IQFOzwwR2Bg
P6O32CzjLXPAoeYy/cjTeOYJ5aajWx5LriXebIj6NWtv3xS1/WMocu4YT860ec4Q5euKa9NhocTK
3EXsnGn6z5Dg695zgMoM8dulgSW1+FLQiEwr98ltTb+GX+lx/ppmeT0vrmJK3TKqf7M913voglmM
4BjMuKu6Sute5/rPvVKj8Yud1rUai1ibg0HLyDctP1mXJpLR0uwHGapHqGfBXExhGePMVxR5D6RE
UcwY1leLfFfOfRjVzzbmubNxY4MxXV97y3Mznxi+5DKjRs/sjwKn5dt2FkOtCNNcnDdXKCdvqW5u
JfLW7khGGYkTAfoFud+LBIEE6kqZjddAzbYxMI89zHJntxrSgr5+Iq71bkMWEzwpQF8LUxktNtOU
d1pB3HJh5MhHwfR+hF5NISTazwHi5CsG/YMFS7CQIcnxgLmdXvs95epDgCgq4WM+haXb/2vGKRuu
h0D9TTcmEW4L6aRFH6jtHG1ZUVhc7YZb68XB0VC3SeR4JxLMcZjtg/j/oB1zckRChfQXhVGd95yn
iSZci4w7z50kkMS20bT45tSaCv1AQjme6K974g4pF2qNm1a32mCkclwNaddzON15RU4PpCtQ42IB
gJ0g50iPHe/7Ws+gEnHSkP5F6i4iPQ5u+C0QT8NDBJ2LyNux8v9wD5MILucS+ehf4zjuomjOyDDc
los90rafgB4Jhm6lzIq4z6+18QMmVE64ijsre2ejVr1oskzcKdC0X+tyx1fNSNlUjvsDeuupe+1F
D9Wi7oJIgkdwEY+Zn4MLuH0AbGVYhhJ33zxQE6Eog/DJp51YhLAMu857KffI2IDGWXofReCkQpJF
fa5gCaFnYz5327zB2jyIgbwZbbzjDpIt0zcTfuC+1cktvAbmSV/HXRkSsbKanvECeoNRMY1Iq1LL
2303g05j56u4Hw6dH/7sh0pOsYuobUTKLZgHugbj/GAI2eVi9NUFD+LR3NxD5dtNr8sJqsxuOEZa
IzipHOIyWKzO6quNKmIlMayoLniqEb0MgpKimrO2E/uMKXuhCxT/XMhhDLfa5xfiuCZO7WWB3kur
cHeubpD+F+84i1OHXSahq+XxGlqmD/o0SxzLy3yQ613FAVLLTx1p5Y9/+yGJfCStAxuDasL7jnSI
J/nnoDx+4MZGtMsAe07/tDr09eRBpcygXFWOX3QbSx2Oh9nywe+LNbfdKaJs5SN+9xBIJimAaz5E
4tm890iWipg8YGCAvul6dd6x9tjGTH1LVc+SI33Q1IO8i/Amfr+up0+vFaBuVt32ZweauInT3DBd
iYRO9gvuBZXLCbr2deb98HQmbr/FX22evpXIVgn5s/Sz+U/FQXorZ6UxaoWoxI8Zyw8B56tlh5nh
9MdyC/hdrMnmtCsFUP6LdkDdLG2SlPL4pVydAL+sef5Oi9/Pr52B3ZSfwZfP3wcM1tnMNe3GK1Xl
3w4X5MjA6/wt/YSRplfo8Znj+3kAAPTmtDzaB+84wx1LrmCeRf4VwI1zmA8007nyYlLw3B5fvIKn
c+6i148q61K84I7OmW4L4yd41IfldNyuLvpwBq5e3zvAN65RxD7tfogemz2Di5PpBnHuqBm1whjd
klc3Le73guIE0m44lZaPoM2ZX5CCxUXnLl/3Lb3iu/wHpfDZ6cfn1nQealBupeScg1PpBlxhnE04
xqr5qkHrpeB6HGJ23WLxs7BoXhkpQUst3qpxpOLsSvN/Z/7Y7Ir6yiyBwv4g1KOpcfPWpY19j872
fKhhu2+xX7YBbXTLoxOe0+0gWatwAsJ0h7Y7HeHlLq2yTs8ZG0MygvJ9q6H69JVkMW8QxXPbFkNE
03V/u6GrOgBHd9W28csCVimxyoCZYzkylTSo7ElqfczMrfsdcnpmlDrqBxNp1I8xwjq9vLu60LUF
3T8P72pHJynqqQ6egEXWz1RMptnpi+xpbrFuj8jKHeIfl+FZcxu0946jV3XcUUfFk/bq7+LpESJM
AyHAyetIyOX07sXsMLt9VsAeeANYB185+r+YJNAFsbTijrWFu6Lsqr7/uBg1D6cl50ze6PshZqeu
+cCMLNxzd2YrG4oHago70lFUbzmbydl1A2Mp5uGZ3CyiFAQwncMI8kOXVr5TIGXkpev/6SUNH4u2
CkN9+lItHwJGZYmuRL8k9B6KszvrhFpr46MXyCBeGNAsrBQwC4DBHwpIx5GNXzDvrBjUAagynYMl
UZqsQ8T9SyWyC9fcL5XLpYotfArTylUiMjxzaB9TZwg9rRAQiQE+pZ+quW6gUG/SyKy+nWlYhnfV
9y2XVJaaINYGFakOLJws+X+lsO+SO8ZkXbe+9/6Z+ZtOpT/JbAj2ailRraif6p5LS4QUbpGrs2kQ
lisDLZJ06vfJrEayUiHKE7RmBub5pOzo64qVvI2bxf9gIFQrw9MHge3j/8Oj+BtyHcjoIfynowJv
DLcxz+AP6ehH0j5Dh6fSEQilSGgrlKwBHco5ugIqRFABgZ2uCD7p/QZmyiJjvuAaWPbTdtEbr1AH
wd38R5+eTsqt6LOsT94ZV+SSJqXchj7fcFENW7gobHcWMV3RfhbwD/E6LQcU3+StyeQfEIbtAPfo
UOAkslj00CPGmMLC/VE6HDKyKLUxGYJrvDxy1ERT+wXC1lhNZS1ZvYpw9hn9Dw0m4OZWXY8rXz4s
i3D5oYkl7zKTp8HAuwMu6+g/bNbzsDeRg2ag5Teou+L7e5oVPfKUI/ZQ8Yb///KVhSl9N220z1v2
7JCigLpfFJ3gWAaRfSKChJYLaoDP8tEFO0xw0whrXYK6E07huQpALsDx25F8eZe2BFyBiIGyfWIQ
4AxC+WhZTdrROuXbzk7yu+eqxnXcKg0HSolV8XQtlDelFwcYY+cuiKU96KnqI08uZ5zofc4jGwYF
hr5DneMbDZUb28YDSBGnG7iRVZfKEBBe+MjcVDSTsRK/QG+gUWEB1B5n+zBuYM4Hj+XJXJRajh/L
U4+RsERe+lfv52H0eWU1AZFU4P6xokwNiIOQPVnlIb6Nz9EGh+m9flzuoCqxPejv/S+iMtGvREZn
jVeXImVU4QVleQAGhLj/+AdLiN5BEp5MTM+783vdrMLKJ4aOTgNZ0odiiyvqfY2tXvaSpIpcXqFk
fo++7wRVr0UJbX5Tic8z7ywxQkz4wyvQQWSAnLnTD6Wl3ZFfsTqBi2bxgu39zjolMDDYyYqhuGDC
CD5w0iotlbnRynUrVQjrN79DMHpJ4kSy6aB9ba0CWVqIj7Q9Ub1+vJGTf69Xvf7OWMvaN2UnJr+8
YKyQ1jUJMwXA5xKYgRRGCn/8LcYcekE2fLdNspHFWP3sXKKVIYXSMKil/7VeA3syHzYRWpGV+Tnb
AH6dItQ/EaBsMlOdVvq+0saADB8HHakjG9saeckYnB1qid9OE0vvcUTBnVdzffzkxtBv4memtxpA
SQtBxuSWBScat9PRe4uNZXGfz+B+iDzjBq57G2ygPZLKNDk76gux4JCxcXEHGXTi6+EpUgpmCZSF
fWkea6gU1ZAw3VcdI2RSk9UkKXCF0epXQqzIjCTTU2T4v2cFkbHXOqCYhjbfSaYZYKnyDPp//now
w9UGPisgV0UZGg5LV+Gr+H7Xod/NcsN29CpdqZgBdJYtMI1Pq+CUNpD0CJTa9W1gqx6Tm9R3K4PU
cPt/STODgGQEQJtjVOlmdLtHN5XT8RGj8r0wjmd/Imj4z0nh41KqDcI4fW1GetVE/hC2BRbZ6u5Y
lX3S2ks0RzF/hUGcF7xOUlIKnPxBhD2ZiQ4wB5TiNub7WTfajsRD8It7f8iauGTvVmsrFa2BWBmB
lpKmzd10hY6SsgNgpaFh33T6H2ZvXa9FRdCOh8UzZhprtcyl8zAZKDC/iyl4iVE2rku/j7XH7TdA
FT/7mWAnbg05NQgPHRl9I+Q/vE+Piq1fCmSLoZEgv1wp6eB7Syek5KE6HFpa6fA61t36DUVo2Eqn
1aWXkzN6U3EfcG1cN8OPiy1EjOZsrFuRxstAWu+0jFkCgX/Gls8drg8NjjpGwMu11xqiXo/3dDEy
SfmMQfgXaMD1BsLe4xYXUQVFeYbrEqorvxcreYXoi9UsoxyQNg/1CurFbOIHPcrQGZpl4C71er5g
lHEEWUqHH3Sx+R70uZiwwH0MKszrk5ZR9Ftgc8DEbV53BNKvKTG7hq/67seJoj8zrKy3weFHXKu/
W6Yw8Gh15UqkZUdGjyD2vJetoHb0qmYwjMwyplYuDj+KXuoU2NxkYjmNUy3ErWEOKZZlnAqJT5bP
Y1OerQKwskj/d1xNCQjrr9gdopNriLFglZT7z4NtU8HKPf9hEMBal6I+dXnuA62QVCscHgNZLj8X
EWJfUdBzaoOavNXdmRx4oj46gW+a9YT696S6WV4e1yBA2fB6dzNz07S0a4nHTJk2t3+VzOAS56C3
NTJLRmYMSWUJJbT5MKVFZ+cY3xFRB9Y2P/YuqkwF3Uluy22NEUG6VBw/UmgFNLIRPdGZoySaBJjB
vGMuGxtoeLNvRFiaDKVMUcBCO5Mm2BXRQ9jq+FhyvjFTteusjhYEgsDH+ZfxmhKEiwKaKC0v+ZsW
vFXtRioNZxLbMGXUJ/Hgowg4Gk+UmUcCnuUOA2DfatRjt3Si6vzLrBDBY41NvGPVoJbL3D5U/Lci
WYxZd/D8q7B2G6xhMpWNjQKSBMlOPGHpAGvfCgT9j5Acg/yubaDg61MYLYSKttmp5gP/wukAOa2w
EXNQrACLCBcDw1cpxqsOGzMRym+iyN9PJJ0sVhaAkmYPE5dt7Ayg9or55fq951ixLNwcnr0DELCn
wyus6KNLaLA84NdadAkkmO8Nohepcj1vivGze4s6o0NI/Zt9jvhnbA/r21/O2XJLQJU0TFu8MgCI
Yv3d1TV9suOKciPrYUXxiCqT0sHJnHg8t1IDw9ChyB1f6m9aGBFvBC7Xi7LV2IV9HkBk248oAQxR
i0CiDZPw48rhOEDjOT5jIAdePm6IrLni6lvzJgTKMtPs2X9N2KogAoYf8DN7D58joo/EJen/n/4E
ZC4IBeZq/PDMA07IEEhINsnNXS5OhS2Jv+qh6STerB1acT9PKyC/XcSLR1GMMK2mtm342WnUz/AS
JmvgFDtF6biunFVA1Vor9b5dmD9dQltkmU7qXLehVbjEUeiiBLMpuKNxhVIjNqwDOpL+td93Ip+7
A3fYkg3F50IbS1KdppI9hGKIb2XxPGG5Uf6H4ytEJ4IglUzHaWNo+vK5h/9Da53hZrbIqNlwPoae
wrMNLOOkKipXsIRe4CWKVOfWXFVuaXZMvU5AiRn8hJAhtDimg+leqJ6BXt9i+BWF8cqNRekOXaBA
kvK4gU8BjbXauDxFeFsWzWr82JDZUo6gM0sZCVqsU/ACbn1J1yoUYGVhMZBw5++gFtKgL+o/qcrW
V+F28ymrtCWieXQ/cALNnzeq5QHNkCUR6TKncqmLVd67xJtGI27pNTFuZpFpnNG39RimzLwkPm1j
ZIU9KTe8tzodjq4ZHTGkVa/nKpO/5AyT4HqsFYIa+B1jDCBJGKYKU8PVaLuPbbDHGNwIi+ojgnJt
QlmeL8yv1caTGl0GNpXyVJC4C3zUOgHL3hEsLwhPGJLdRBjYj4/8eoTSeDHTEVvDzsGG7/k8N6jf
W+/Zzp0bfli2azW4YionTj5cLGjy+ZUfoXpONejLNHLLnqmpjxs72RHCUbchHICfjxrT0jjTlFO3
Al0mLb2dtAKLLwQF0Xl9FjK+GJIvpf+8aMUyZjvTr3zQD24fVYBE/+xxqGUCTUk1IVizJgwdfOht
PTWG2F2FejNZi4FPT+jhdnIL5+b4XcKZktPaD+HGVXDmN6TM0cqBQTzXxeoekI+Ne9sbJCvP153n
0Ki4XTpUZEAk3uxaDuVBJmRiWnF8rG/sjtfeq0XirfFo5pMF3QZeQKx7uCs2Bx2g4aPLvUFcXXG2
sHfnnfm9eatpIYzlJsqIOGyPym4FTl4NxaPe0+T8DDzgrP0Zy9C931kopk0Kz/B/Y1Ww0uTyw1/Z
/ILsfGjL178ds6Y1qFdB/dJfO8w4sgXYi9aVwz+cRCUHM/i0U2C0uTasXx2Q8RPdeAiyw2GWiZzE
GVel6E619EeAixx13jfVL0ZXKWEn8ifuger0NskcmarwV0HnX7kopNr24X/Ri+QTAMP6uIeu5sKq
l/PFXIpvqCPn1j2vJt1uVwDNZ8hMLRfiYeLnWfr8da2yBX7Ru9ph6KynpW0nwQvDVP1mcSX4Jw1B
6Cq2m4wvhYuFcxAJsnCYi2JKm4UILmxosBUW97d7zaWtzpf7eG1W/h1sczv1Nh6/s0Row6XhD/pY
fJtJHO2rfq7sATect7Rx9k91D8ZMitBrmNivtKZETaZR+IxUBfCjCH075HKw9/vaURdJYFAaTFBj
JXMO9Bo/kRFve1qB110JhFClnl/Q2GSjf5olt7Jd23C6NjFu49rN/+awCY/Oa+N7JoftHzwqs9Gz
HA0fFxFa++W+6UGYwZlUDnN/R2EGyQRQyGAM5usWKF7dyxwHQRmI0godwYFjoognL+LQliTnwWPh
OKMDMNOmt3eoN7KMymnkGoxdo93Qt3Fqj6XsoFFSO+qCGb+nQecoPd28DSbVxPvsjyB/u/hdQs+E
r9KTb7soZ3wEv67Lw+1yIda+nebVXOhvDHVMmTGDkeWQhgE5gpiKanjd1EQbfJz7TSLx9R3RBV04
Mgezr9Mt8bkVW6Op/EIBiztQvPDgjh8T5QTQiQeU97t+s28cKEs8YMNpnQltUL9zyzQo+ZB+X/uY
Ighz5hfmKUl9Oe4pl9wUo7aZGd5wwjA8rjNgjxb49tzVjFz7ebI/QZ8csq447QO21H+/SUx5jcNs
IaU8WAykn2NvhibZPao8SwaNO+mTk0SUM27QvI7bxiOMPyslp1kf7mTqZg39lKZsubdVBlU6T2e8
DkJIKkH2Cou7CSlH43+bF2gCe8i0Mutid149wynUy8Pyr3+Ky0KNEOyasbCdQJCW7bPRZqaqNOOO
nbXUHt9u9ojZIEq+1I7yNfz+0NvRSfox+/9vbqepjDnhL5/ZgBKbqgH7yL5qakwwkdUEikyFQBat
AkXG5S4YX81f4cwMwEp+D6mTjnqTuLsHFNZy2UmbvFft1ttAkRzwd+W7NuC4zCWe7iQuyrjYssbB
d9JE1/XuwPDVsY4o5HI1dyLGOCpddNLw0vTjtxyt1/KXU5mALGlpzy5NrmDtIHPxtpLgKBcdV1l6
alI1f5XfXraZ6ej9uqxcggdlEz67tAunf4tetZ0118F3yzYyaK66OXW3VmpBPc9SX/LkiK/B/j7c
y7C7XUxcl+QvAo4DioEzequAStfXULhvVs34NUQnC9L3FIEat3nvKZeWutQCxLkw+MntDz+jrZWJ
faD/t4OagwiHw8+36rbx3CrREyq4dM92WxjmCdyIpZ6s+YrScWDmWmGABKoQ0ln6+v0L+HyKGsxE
9oq6ih9j8qjue5QCHX2QXGbs9GGQrm3Ke4aNBiecWPxDxnRyjQl1F74m8XOsv3DWZAKvuJr8T1+S
Pe/0lnYZv5k8JI+yPiCTV7+quSxXx8drDwakb/upU5PcEX3QgCufyB4pzbBv6kizLZ/h0zM/rjgN
9oeHn7OirH5cRI63WEUmIu7H4Cg2Wbh9L8kJNXn1qMo9JsN7QMo3ov9WXWL7IR+sNRPScdaq27zj
hKsBD5CXXrjk4dzkh2j4rWzHa8WwouswVek2c+GgKOFihKJhG72w5aGkkuJFfzcnTtioUMShf71b
6QVwLLjdlsxJN0xBqA1of2q71SDSIBmFHrmRmAdWIh7R4m0dT9pWESnP6Ala1Czv1nNMs383gO96
GsYfNGhgCEawwGzd8AEhDFD7ZptYvTE9MzmFr730G8nmmq4VOoBfi++qSCvwwifMoM77WLcxSrrM
qD546uxq8keybUf90MlIRw0Clj8wqe/dVwKydkJV7ncoqh1kKUKnebzqGu+XbDqezw6ddK6wgNQD
mgAScFLgL+bTCw72jq32lWcmqjQwpFumSwZZ0FXgzgglLQfERkZOoZEPQYc3ldIMIhV05q3kV9Uv
XZAW3doDfAVhkucDa/oIRbBqgeB/K/r4B35nV4B3nyu1YdPKxehLDOXRQdrCTU2M/EwRbkpwPV7e
MdWlAg9vqVuR9o8klWfYhsji2M2rp6BGsi5fSc26INiWhXmTvuqjZGP7zJicGFo/Rll/rUnjttbY
cCO8VhfPZUeTXD9bAk8nqvekSS6d+HSQuUZLY7hixH3QYVEpXIh9+T/sY1ZHGhpLBMt1gKj3hXsI
qED+rN9MD22Y7qKvMO9C3Ym7YDy3Qjnxh6gdrx8dnjazIchdYM+aPsgO1N+RpYBn4Jg15oF2MGh1
KfuYe2TZ28O6QafkWDqqSDHhF6ujKdP5YC9nDOXV1WPckMdwGxSIF1kWX+3ph3mWC0NXKYslOlVU
cnRgX9I1rj3v25TWnp/IpH6tt5l+28Z8Vd1Hp5bHc+ZyDeqws8aEQVEkU0awlliccIf1S15dCJQh
16VWp4zfPTFwMGjAeHf/jSjUGRwmIwESrfyjYy11W2ki5mQx/srzGV115zJh8gIGGEIYLTZL+x7o
TFPxpTRSg/alrPuUqLPVOsIxVPiVWxh8c266FkwhPKTc133aa5zPcgvqrGGiO4ZdQSWuGHSiBi3b
g7O9qQfXbFGK2VbudA+vRICfQV/n9h+FbbVDPnnMnil+pQZCYeP10GDWOkkjCDtMbfra7KBZ40u6
60i97sLKVg5WsXIQl6Dp8awv+Z2UiZj9UH1uaVNpkoIl4ey7qfsnmaZaoVXpmkz6Wqor7pvF5uzk
/lyMVSAKjPPVrNS/ylpkQvsvzhew6Efg7fgs54CKq6IScvEcCi+D4fKjZzRHQUs9JzaDKZdLBM2f
zf2eO8wd0YVXHaYwFvr5v5hltvCff1fCdmdK0BHAv75smYXOOBxDHCd48lgGOUYGJz5Ebs+LykhE
hmE7/HC+Hx26tDmPLRky1BbLaT4/GQCPH7P72cwwpV+NPAi+x4c1L028OYD8lQRy4QEDPEwWISfB
3pQ97EY8r0UEiY3rgYH5EQuKZ6PVmzHXf6gy9Bcdpgr8lt3bLFv3Tp6PVGLYvqrc6kdE7kmdYoQ2
Y8PJlbWx8QhYWfQcjw3YVO/vKVp9Fb0VqfBRMWY/Z3N1fUWqB1GAivC7YEZS6TPqAORP8S1HBkcS
mHWtIELiO4qigRDAhBLT0cWjhdhUWClrEsv196tE0M0v29mk4fZ0Lu4cFqSBjLroiETZKFt+v35/
LFivmTP8oS7rkDswbBdH0Hsqu0v1UIkwuhNibRQq21wAGq++q1Er4YiSzDV08hkTbAeQvBTa/DvN
BjCCbN3LvM8yxJiZhapVKeOYH3GRL1RWd15DroKzRQEO0Bwhh9AnaozdLrSZie5Q/UNXS3q071P7
cxy0YSOciuPrKq3W8U676oFXKGx25ERTyH2O4nosVqNWbB/+Wnl9MAJ63EP72C1pEkqsAlaamjXR
etZG2fK9c++d7I9ECEnB4go/mshLcZ9wiM9negUCUyYEHUv1V6AXLzzi/GDIgp2uUE9k9HQXNweB
QOgLUV2z0Z0mwRoNdivqFm4TM2z1qRaAmoTiDADpxKK7GLayiml9OJ/940VTP7QAYlTEvjCtaNXz
f0KpwXlzmVZbtigEW0/roLhQmhRn41LQkqzdjLqaYzy5kkm5QmdqXAk2w5wsBqZ7FJhCQQ6KunGd
jrYgxXMtBjw+MxpC8gruD9dnZ+G4MKzWlUumbgkOKhq1jk/FdroBHs/KhpqdkhpBlR2bx3ZY9KJh
giMpbJkqAylQm9EHvYmkv6ucQW+aJgvT8hV57vKz2XCta13Whh0Dn759nJIAmYbj8NUW+xC9Pmzq
pQbCrsX6ZEMPuOSXc0nAXjrBf+lGzBBKqpEvmh3qszVMmMWeADchkCNCrY9n3lkO5DbDvs3XfV99
PUcNLgPqBHCFj9TRUqMxBe8Kft6MZsar771SVIUiVMj8OJTYx+VKsbAhod87YcAlQbwnXynXs2XJ
AzmWnx8PSk0EC6Mkb3nayANZV7wvo143UOdEZp7NLWX6Hm9DV8jUScFnwhjB9j7K+pqPTjsIUMSo
LI8FpSqTiWWDCQBDWdbavG2yR3CIr1E5KZ54SB2nXN0e7pw6PvxEmm4z81pG51BODN8Eu+ZAtJS1
boU/YT3sazJ4VNIq0yi1fBdpBYcse/pIGC1oawY2q8qcPRXIGFoiY25DLg65LapKWdfAe1nip5xX
PDxLhQ9rYZdVIVnFYYPZBSy0yUdy2eI2Bccq+vNFI6SRj4w93oQlg2eyeHn81b97gHsbQzSLhQc9
izBSfOymxtrlH0CEzJhJIA4AOQ4aKM/ppc3ntWFDZKjBFupOTPr1rG3bPFMip0OaJgaDOrX+8Jep
emglgrIBGyoACOy1QmkPkJL8upGQqTSMeFAG4wJYKnBiHCRH4jEcILLslk+SJrC5FqBhvli1kU3L
nnPx/b2mbr7QKMWQCKeJXSHL8FfqqDx6U1TsKHMZ4CD44/6af8qaS3e+F1MmpFb2RF+CDUGVzFfS
uR6Kvy6Y5O3R01ZVr0aoKxZX1YsM93d7T3UrD+uOpgmqOJBTzUYARB6PvrXvCT7L3I0KM/ZOoa1Q
CCAkU5AzEf6QH5Cd3RPv/j9+4GaEZOtsBrONjji9DIiCubLNNuVr4no+2YIdHPAhr0VT3GqjvyFM
O30QP1tq/2HXnAsaLQDPtQCZKJAyE2e5n8LXQzIE7qU0W34Jk46VM8FnvbS6Ikn++Ob7S51yuKIR
52tTmia1HC3vqezD2ksF9m/TUu4zkkqXmNIt3kOtunsl6acK173esf2aSG2w3Oa8QBdQY15/AsX6
CoVTF2zvkDrhFsNp3Loovwj+GgTqHQ7b17Xnl8gqBIVqn5djsj360ltekz9cb5otLvUTqlzCrnoZ
635zlseR3o+qD1GmCQMbOiSdxqb04Q0hckPj7T78a9T1YkihzDgus97o6kMh7VmIO7So0EQH3aXt
uOj8laOfKEbz6gXumcVRncnuofB95kHfGghr5YrakPWIx3HlcA3oDNXa+uNvl2/Qsu8iznaQzODP
LVNlX/RSGwG68r9KEGQsjiA8Di6wjWuLE9f67tjTlq5fJYexWPgi5lUnw6sUgI9Xu0WsYxx+JKps
AEPrzBkk2Ra5WCVwuHvEaHTEvEvU4+YJvXyC5005bA0tm5BvhsTJo9VNAcR+hPRzkVoowNc7W8UN
eCn/qM2xuZr5AWiv4j2MKDiEHC/a1xvSszrTkkBNnkwyfwKHhKBMzRy9AfQEf14laULMUTB3VFLS
sFncizdVHXY8bv3Bnw+EqMd9Q6zol1sJfy4RmahXS6QiyRh2ZVnGHcM+iKVlR8wQLBSkFUkUaSFu
47txA48yCymV+22rCY/h0M8fQz5QAypxY5KOo7NTQiFDX6A1TYyzVPJZdbTkiPlgC15js9Hd+lc6
yUzmVi6Cn3WEsPi1XYvS2lrUVpAPxLSQr4RzBorpbcItk8prKMEYtS6kOM4lS+e/peqCtYc+YNAS
RTMyQjuC/YVR11UIsSm35TyCgndmssd5DgxefUksa40WO14am3vLN/1+GuEHdUDQCizFy0zNk3C6
ZXS3t5TL2KI4G6GWk++anbMN/W2+QdVPwYuZVTI8cOZ+RkfvaF0jaxYcmseYknF/zynyTJg6nMRL
hono8RjLu1hgDqQQMbC6RCTF7IbhkfGsVkXVga0ab9z2czeBjwNTnfel5mr6QEn3m6v39G2pidpG
mF2eUfcQEM5hMuP9iRp2plT0T9/jAS/qeFRmQHw1eya0Ktp6JfFe4c1S8GE/xx/wNckOnN/7IHiA
0Y3NQwBl9JUTOWzN7bvUvufUOQGArVq8bBszMG9HWm9Z1BKDM8HR1G9DLdgyVS/gbgbygqpGxCIF
j23jN6IzNkkqFdi/exeXx1xYyjfKrrCh9RAXuRo4LJe88QQNWFf/YSICk0rACO317ApgqvP5BTtW
vZ4xTKieqhSg02tljz0JgNEmLRMFItfQ3LPL5u2dxC1yEMt4DASRVq/ckCK2DOujHLGnybkUhURo
iC5PF7t/zYxuWykrHoigKE4TcV50yuqD1ffz3QyyzZrrpkVqWX7jWZf3cqwvN3asgWXHsCAuyA2t
T8I7Tvd2NF3krAQAp85FDpj27COGCBjJFYKkz8c71LpRFTcO7T6mLkzm6+86LuJUat1ksuGNuaWI
2Z1fxyhBhmXnmtzHpjlB6fnsjBEePiYhf0PeIpuitZPouQ0Hez3pRT8oHRk82TIDitZwiqym67ak
/o7ndegSkxcLYdphYkEGAUnhB2r8vzcrhQNtnVbGFWIjddBMn0kHhm7rSc5EG3+eKhX+jD0gGJ39
Npz8iDFt9E2JJ6m054oNBhDFzc51fbDsNretqzso0lgXE55c1GX92Jw2aXUeuLhkF2rSJ9CMO9a3
AF619usW7JPd3Wt6Dh75eSBuUpZPhTPLoGawDyHArJOHajCrDStD4TvGqspOBxoZ4Tu0F8WV2r+c
rFABe4pL4zgUZobH+Wfrf0gW2Ao3VjPFtYVJ3TOCvgu9arHfon6cDDFjQwYRBSYjFkPun0LXvUcG
+Fg02IryUewAyNVrWVwa560X5umQaDY+WUWZgvFKwzA5lxfCcByIfXVqTVmmjFoEjcDxEMIj9Qpj
TlEqHN+afHzVcr2VJui3Lg9uxfAHY4I/Q+qlsQZJW9vak3o8tLXF12AxgVw77aSm0A1WYG+VFspB
f5QFTRLABdCkF37b5RKA/rAum6tKc5BL+KBuP06owW5EDWXUcrfEm9emUzo/utiZW3txzZgpa7jE
KNqoJNWGQEtAbuRhLK1h9Q8/EX2KsCcdfUyXw1DgU+wc4CZl5DzOGHZlhG/xtZiHkPVet0P5E9HH
Pob2FqFW9+iV0cpteRv5IuLmUrwI5zyXPT187+m+pYKF++qTQ93C2cw51hCMJgj5vw0GpbdjdQw6
zhAA0HMiuh6CAwgvLY17mzb9zVhacBLf8EAQ8hLkl81gmGQhuJHfbVrUA18rZ7BCDnoWNU6lTou1
EI4tFj5s5FUmmO3f1PtVwcbAIun+I0HHphIWBRW6VN0/bakattW36Zp6vVrlBksPeh3RjKErwWfS
ZwMDWf3kL4rh134fOhWZtLepIH/5xz8yHJignxTYIGiwJmTrUeiw2ywJaqvx4Ul4VnGZ2YfNAKw/
BsazLdZCgw+clhn3Xc20W9xbrNMS8LLE4svYhfek+xKTrP1krj0+RILQNPHEzMeDvx2PD32Nd2pE
ctZj6Dp+VtuNNOQ1iMQOb5wTAbReu5C5jPTgPxpH26XvCZc0OExvbqw2WflbOx1Q0HhmxGc8FPHp
xSXJlU8xbmP3MB8uWJJ2P+cI1lpQwAgaQFMUORZpmDZL0AxaoWUKHRxnr+tArC3VHGg8SyPf1HXb
3JyPDIGInW3I1Nlhro3lzpyISRpHIep6FKRQz64QYyD4KN/5oblFUTEvmfZo4aJ2dMSszBxLXkVW
MtKMAYRafwyP8Tjb9tI/F/A2UeAG2pFgneyfi88maHy0My6gVgiOFlXFlanKGqMXJb/tGhO6WNgo
Q5zRmWEVVMU+nR5oIflPOljmMU6zjrCVPtjaj6Lf+4h6aiEzrGarlXuF5WILjKJa6DxD/EbHgEkv
HU3x1JzuhNuTwUast5/JVkkE0V+DeX8ogHizQUs6zBXUS+3y1b6wkgD2aePLBPEv2i+d+Un90w8T
GlnFLkyELBh3mjNPFaM8e0GmQftEh2OJB7x0vHe9IYlQlh0QtAJWW8txRWOJ88RIyNMJoBtpXWVM
6X/JC+j4/06/TRgtXXH/WUmLhImQGJ9Y4PRRy+yBxQZBYjvaHiFVKgifn7sdb6Rf6K0XtSV1ljZT
xzvntDy2Z4EfMWkTMo1M1ZpSNeKFgdqR4ZtTMmyA32NMjMeUXakCXWZwTNjzQCmwaRIMCnuD0iPh
BRsqX6N3S8bFqWzX/NsJF+zCfZLPSxKuEmAwM4rjsxNqtRtjF1nnI847cAlGIj5hoO7biBWNnTSM
tdmfF5mjr6u+9Qu83PCN6a7AOl9CYgDGrwYo9cx0z8UG0wyyAFjZa12ZFIPVT7CCQZ+VAWgZJQeh
b8tdh1o7GDD2kuyS4uLZmdYXG/5Q7NfIjSKT3AjrY6ePf6xEfgEFLi1MbuXeX9PgTS7U5wEFYFzP
tNU4cp4fZdeZVbE41HaoOH6bXXbHhux6JP8n1lMCFMZfIuKhrs9MOVURAbSW4DW0YPBtHingWD4k
X8XcXmnguU54pVsJKBTzD4f7hyh/JDGfCH6zfmGNdMv8ByMVtwTe6LveNui2OCgk5IqmDrpkY2Jk
yW3KERc/2VxgMwV6kxbOr3yUHNxD9hhpChusGkhPEnD6Xu6q9FP8P9sj53jbVtrXdLJdaCCdi10k
9Pl99+X6MC0bcAE/sqLO6UolvcorMenrmbHjXGXNKu6+CUSOU65BgwW3Jy2V9DbrF/1zkekGUxKO
lJ31TyEQrt+fAuTa09U+g/My/plZuL8vGsbteRAqyn8JJk9Z2tWGh5ISNq3RiEXkZbdvzclTIOXu
aI8uAnset2rRPzUAraw+5KAXLqsPEqLchiplpO6EVvg2M1zFVR5QedeRYzRKIQRa3EccC0BZ6YSj
ifXeMtjt5H56WJLso51DpBtgAWZ8W7XLiJ5+cO+THHALUNhbA6eCOw5/Av5MB3V/3+p+Ai5AdAM8
p1fSuSCoz84cwpQG3xy7zxD6fMvLSVYfWNYQkrcYxUOHNmAPh2xuWs5bAvuS+145K+N/UX6BTMCO
pHfldJYy3GzlAWUj4KIXDIDWrTooWgrRuL+MWsrnV8K9ab3tlbQHUj+CiTBMI8wj+na3gaW9DaxW
dznXqC1OU4g8Bl5d6BEIukzTX5ODiYwcOLWrJhF1jIIoGP5XUXEfIB5Qu/CyZKFSzYMiRSH2Ut8k
bJCqqYvr35QpC4+hbZrc66hrxXkHUzAn/1BhGkd+xTvieZF4kZYkoWYXvuZBNITaxo7VI7vA3dsd
pK0m5ZYe7IFB3YVW3eLhEhQrePBRocu3CuWfgYJpu7SeyL08VNLMe6mHclv6YQbfQQ7nfQWMn3Fw
PLwij2nDYjr7yZ2ZBfqZXrtugCFoDbeYajvSL0h7DZ3zw7GTz0XpQ5OK7TI3rqMqussc9k6Nspks
DNpAUnXLB8pM46KCpkfovVM5iAsb0dUEf9LEAmbh/zi6Sz47ZpIJRMn0KV+PZ1O48WRLy7IPWxfD
ITd4UO7X28FAZLyIFpG8hXv42YBYAOg448LF6TP/SW3Q6VKyoFJ4zdwT23xmJGTjrbpvV3TJi5Z+
LwvctaKrb0zV46j52pmGTC0FN/ZqUnc2FEnNKYyjmT+rlxIKLP07wSVZ+kdWFpYw6+i2sYZoG5GE
71ZLqyTRW5mG+PRuExBweWNDjqh3HCPWFCoudyIb/UPt6in/bpFhBmDs/OyeQ61+GY0+Pndfw3A9
Xezy5Ot9uJHdTbAUvfmyu2ykith9c7Qe+Jp5hpEIcWx8+QKAz2jCBXNxBpArpTMQZTs7wGFzOffp
cbGyQ+NsT3BmbTzYiAe7abo42ovEIez2M8mqyLdYo1W5gRNf2SztMmSj1KSIJB1pYJceDlgiGzJ5
9wu9grjHgTbqK0/Hg1eBm0lwvWEkQoVLr0orzivolYs+ed1Zyf8yML2nQ0irlTonxBZRPyY9r6gz
i+0eXOUEr2kU4GyKD/uFxHEhU/mun5c0GHzGTegN9iMXfGokcXKVg01LjENWLknlCx5nS5we/4NM
u3oMHV9fmwu0PS/eN0BLLolSfqsh33TcbzPqGnf/PKewkU/HAf5MOOYuuk/ojKio28R1G59W+3+H
74D4vlu1paHzdqQO+inbRKzLDPg4m+CbPl0e7AuGNcVUd+JGlSZ59wQ6vuxuvfeKGblCwzwkCoaS
VZ09USJFRONecxrhGq77vqwtvcjBfLqX+o2Juh0dYFXAhMFs6nGVmZQupXJTDdXLSGYlpTee6gF/
tFqBx8i2K/zUFvFWyO6ECJbkp8nOx67Gy7ZqO6AVj4I8A41cSvpifhqlTCDBXrszHbiD6aFasqn7
2eFut+EpuWUVZb1g3/WNUY38V0rHd7AhwfYGqcCSi8jmoU1x6YIUTBtCZM7ng0cn/l5rk4sFSIwu
G9VPShitqDew+nx0zn5mSgVKYjbzcn9I2SWh3jinNss/+8Ak1hX4WUnOvYGprnhH8vAN/LWZmT8l
v63txkIuwjN0bg87SBm8pfgei9fLoGWeKymRO14VcW/Amtxljs/wa8CieKMEUY/CtXD8QvU865Qm
GnVkLQ+xMWvTbN8bEQKAPMBWnJj0Xf8Il/53OoMQX9xpADWcE+RvlZJzIoLb/4O6SDNEIk4EVzqh
duaQ1U2Fj6ztFmoZ5S6Y632ma4wl63kwT2ayw6nQ3yRgJeDRYYcwVstawxcG87mSa8/nhRRdzI6v
lJKE8wSFUjeMT4pqG9sVCVYtpv5w9v+LDAaHCFNiSpBL7oIeLEo9Wie4Z9QbY9N9e+AKs9zhMXcj
9/IQ2dPUQF7EkKCE6OBOT0HIDRTahGil121f7aqQbLXXYaOP9Apoc7+mz94NL4dOKzbviCEx4UF+
NAwTaHf2DibaK3Si9rLoSuFxoIMGHPKLtAizj/UeCFD7eSNGOd7bVWWlc8BdzOsfTDFIAAybReHZ
ORjbjvC/efLKDcfUynRPv55UVIbSaw48+uo91l/HZuwcvt64f2jgTXOjiInuKp4p1X+/9NCq32uf
lCnpIuucjlOJak4IEwNe83LQd+BOtAzvOyjBHXKFomHztwgVxFueQqsUWnrOmyvRarH/fylXuy/b
AiSbHw62rjkOMXRcLiXJQmMUmLm9WO2A9mp+pK5S9HAikbnUI2GgyS+Hruv9etiejMxWPYwodKF7
45bz/EDjjfTmZJszlmLsD83FIoW4SFNiQbRYLssSJhfG4Kbyx/r2jsXxqBCOUHHMVY239D5YBWm6
BL++EvzfLezFxwN/9Ae0GQUdhALLAxbXVJdekyoirYiWS7M/4zxToqAa0JJtMmmd2c8CwX1obb/S
zwelRwH2evISryZfxnCC+GE5ySyzhrnF4lqCLKwId2k7yGIq/Z+GxU68EuKXdJaOgZys2bpk/tGS
35gMd4OHIERB8amFKRRi1utg3JjhBQ4WWQgakfP+tvyZ7+io7Q99OyqjT/dUzFMhuR++0mTwGDf2
ivUDHyoi/60991F+ZnkdzKwrSSV4ACFZmZY/PNvvsB7n1iupxFlPDAq02O8e4PSPXoVKTOJrDBr3
dFryynp4UdP4LmALrUfa9GyMTSE2ObbXF9Wra5ExrBvRypA3VAWqxi3Zhfi4Kvi8L5CDzDx8IL/y
vDlb423AJcLkiw9wj5qsSQOD9YQP8i2NhbZWLsjp47le4IOddGvODWXRnBPP91IH3hb+AtVzaUnk
cGTfJrDGUZ59tU/e/yg/vIQbn3BTG8Gbr8UwohJIO7w2GTQTdwMpz65HyrMiFIVoDOiOioHoPI/B
Bvd6C4zYNT7aPV0RMoKphECTBfrGUx8ifHZ6UdnF36bQ/2t5bFAKgIIYvfIskzyqiU5Z5+FAJ61/
URW/x8MAqacSqDJAeAP9e4mEWYK+50Ekk7VaK7TZTc+1ITPe7XkEC3sbDNleGSSSphbk6qy6JPsa
fGqXRm968VM1YSfMlqWyzJLNRUNJZFK/Iu82V/HKzoTOBfUlRichLXeAWlC6LxTwb8asGXFljlSs
aeiStO4QHC6O0HVFkNDeknYIAjTLa4CQLvXDfATSKNXHqB1m2vE0phmITYu5Zm+Hy6Y3zL9FNzTw
imdix0sGHVry/6QHQ6v63tESxOcp2Q9TSuD+UaS8zhqaAfwmvB67DE0DOkbZ4NvmJ09BdYMiSCI1
Clu8aY2P7tjd0QSkPXnGBbyRjt17hD9HE0JMKfUMExd/BC2I8GrYeat2ehHkbya5uSwhBvsr+Lhq
uxUgHJmAZ7xzMjqFNhnm50KddoZg49RifwHqXBh4fZCxAzvc5qvnuYg7r+UKySznC6Citm1N33hr
50G3k2KK+qc17XUDrYUOzGmpLGugI7EDXq/2VSNFDmcVGu4Wf3qeQC8Wnl9h/ZZPJgVmhimcHIta
M+n3pDKFGRhthrCkKneBzPPU4K/IBeTvcqivAZK9mOsxpQDCHwgedC1yCBnWHMgyJAZwY1I1Sbmm
UOGv2tHfB6IC5CCQLOosaAj3C3AxmO5lZi5ktdux1ExcalK/MzStyEGpb8zM8e/g7b0KASJg/O5z
53bKoMiHHpZnc63a74hBS67VKTMXlZ9ShZ0UvBYradWsm35+whU1R8SkHKsBsfKkmq6G3Cy7nnZh
/p6tToNHb0QBvd36b/4y5Sujn8LHAKC6M/6XQqaOP+d05DkE7cg0iiJy3ScTzAvhA2vOaMEkl1sM
CHIqXO1NfVXF7OEA2HiW4BllOWc3mNoifgXeGjYSi2Y5Cg0JgeMNOWsXR4ml7oRv+5iBaFVPxwXB
ynHd5MXC81xcY+qU9hisfo2muMmr+3lAQ7FJvtMS/DEGcHkJtHKKL+nr7DX4fLax6vYBaxjKrmZy
bSXiLcJgNFDQXYug830GcRgcv+CrXoQizQSNwJfV+4N2r8JmEHf1QJC2EKqLk7vJxP5q3OeknGf+
sMYSlACc6bzC2EUljdg6rxg6w2SlMCbXlBBnEVctkgL4D8hYCjQ/97vuH67t/EUFPjgowh/cB1P0
lKAApiqTteGh0F4UJ43XR+4J123T9elN2Yut7uI2MEXWe644Mc7KW02QjaQyL6Sy+xdLQMqUQgG8
JnvItlhLyZnQcbkPqE4s91ZxPYEkLxZ+mP4aozEyhIE+C6IE7R2w3J8H5mplyp+9aQcBz7H1oGv3
WL7k55XuM1L5KNwQJoJAkg7J+4PLmEqF7FoO12dP3wPXyLP72N1Pg6iICpzV9uzkF5hClY513kO9
s5kN+ZKFHOwQhsVKs0vmU85M4uEM3MlrIVCAu4AqCMsZ7TZ9YHQv6AfPsfDyiKfbRZzrCM6wcdXC
mrYLyyRHD4XcP6yeqRsq/6jBYCK1DNxpDwO8n8fdT+0lFuztNpUX3t5/qlRewkNQR+t73xoB12LI
7TT9GT6EaWzHrr2Hv6do7PjxnGfFQKauQ5MoYE55/nnw15qnDNzcruVeS7MqDqi0xXqFqrXIE3Yw
AckoBOGCDfChP/UAbBrDHVX42EYH58Hfy78UnUeU5kYOOcZwWtP81IKBzUU1xO7l1ml4GMqvCQON
1vEheo0jJqSj0LmAQzDi9nygPu39EbmkrbqqC6wZWd8vSkPjJl2GuHBXGSGgXUtXzvytshsxjuL7
TXRVCjvGqHNTsn3x5dh7FJfJflvhsXdpglYzIILVenZDQnPtYEqUALv1/24SRCDMxukJv8y1t/Gg
er6Pk+knA1CBzRbqnGxkMGkoeb3nWRBFIJtzFgoOn0sNc+UdY4Y4bDP+YgIW9H2AYCBtBdKZCekq
A3kbYMBkzSNmf+mQPWXlxQZsB4XECipHuB0fUAqOltpAEwq3i9uf4prJDbcZG9VtDpkYPfpg3FQ5
nwnK0cLDfjWqO06FWXOfcCrrnWem/rIjRHZeUDn6Pq7VIMneVjNGihraUZziMOJeR7wcwKZ0dfhx
Pg4lIb2LgeifQ08mZh4TxBOgnaIivKA+9F8O8bdLBeqCAcUSIhp27uaPc2Yw7XHOwxWXNswqIdk/
KIkkSQBeZ0yOJfAqnWNvRlGZy449CxQ8QMikbilAlhNixU3dIckx1TwnHV7RRskfqH+zR8vWOM6z
dRHnOfLfg1cYoSPKkRW25sTmk1aiH9g15SUqWfaNvJh46R6WGd683Hx8NQeH+SntnF7bIocE8zlj
98eP0n55lehnMvWg9qwX4ZuWtQY9W1fkTx7eYiN1tbH+Y1pPI4cdNucjH9KCBFe4TK2EXIj/dm+K
yvqDRBJB9qQFqN5hcCvFst5Ofcsi9HKr6Dce7WGkN5Rsg4tAhAM+WfVqS4Rpef1sACCsApWaa4Ny
F4El73wSEfutfmvM6ufXyBrvc9Bammbjbf3NSG72ozONNDVVdfiEv56rl8f8r64PfogCF+VHH8O9
R53yBzH/k2u1EiCT7mufIcLpIIgDGNl//jPWxJMIpt7UuG6l+29PWG8EAst/mSIkog63WCdICg4g
pJvAXmzC8MhiI3SnBElaSYKdVMBd3HrCKXWHF4+nUrdE3VUHQh76PAEst05Xz/Cr1AN4yRE71FBm
slQs1YuHrv18akL/j2bcOEj1xEY+3Atc+xxPzyVtfka1EsgJEKbhgC8lcg7raIDDA71mbbRFCbM6
c7xJNmBp6SsCZe71OZR0M0usuH3ToxD3RoE0I9oVLC+49ucgHulS39Moc7DWzC4enrLakMuBpDXi
8un2brirSsZlH2Hl7BUFjUSPmPt5f6PgukoDhzJ4gZ14GXmCEWH8cIzUPZDAi4fkhIctpH3khKh4
fop0BrtoVCn1NHZLqYNLmeDpioqAe8cKllXKD5KrbplG/wPfILz/OYoB6bwrzwesfKAybdkbdZ5G
nEgOtVmXh4tCD61ukCrhjw9J7Vf5AvYTnTsx+di4mZG4o1LspUdXdiHkdfTyVBCTZQsQ1TnZxzRg
sf/yaJG6yotOuzAWtvZSlswjNWVhTFQ955GYBNcxaU9ttNLG3BdcqOFtz7ogzJlURAy/XF7XGboA
bVJpUx9epsg2UKmDiR1nb2BliOcrqe8a7LKx4TdmreNO3OCgGi3/FrQ/OyotVmO7i0lAqWNKNGVW
wGEAoNW4j6XO17IhQLX+iQPqSLMSXz9+szxI888EVSm4c/WT/moU7tGuSv0UVpgvJqhst4tWD07f
Uf70rVretBi2CwfUTOQoMQk06BJcfSjpTrVU8RGo2mYcy+i49u0l92ihE1ZkBTosLhIovElqmqkC
4dzfy/dfUzOtHaTfirQ64zfPzJ1qMsUu8Zou33En0frqqfWIu6/TiYzy7qYiUegwV24uqtnaug7N
Z3NLc+3fdAyZsTgh4wxwJsnlcFJ5kvHvNhpccokKfcMayToiyMhFDtrUK33fSLqER9DnRStVfT8T
b9sEtlg1+o6mH5ooRYGUACyGmz7ZFE+o0239eubUT8+4RPjklyV55vz8ybV8MWis580KgRSStx9y
iaZd30wW/EH+wSJugwnd07GpbUvAj84Asbs7hC7q9iBEJ4n0/+XApxQGbV7nq6WaZAbDWv+Go4HX
lRb7+dxKpWVikUE56AcB0N6D6y3so9pbd/qxRqHot98eoeDwrusUecUFOz3eFKnxyS+u0N+rxbUA
FDGkcyRFl07zd9iOHCXsf5hrd3Hve59LEZja6TCUFqma8s+uxIh3S0gyDLAbsf0VgBsojX6NQFQ7
iQGovJz4IbMBn+jcKE7t3GZUuBjtoRNdK83KBnq0IuFYq23i2vl3NNIjg0G3W1CogkfdwnL4bylV
k2TbsUFko68AU+C9mXicBGtJcHQdZscilRXOVOX93H7KslHciSvHwXopaNEmJiroI2UtCIU7lg4x
XWq70eYHsCFpBpT5MUZjNum5OkI9umRbJoLJNbYz7ztr0I7aS+vu1jj7Cj5XPip3AdlD8CNryRKr
bT1QNFI9tSSN1sBCgRkNvmnp4m9GEAmCXsZaB4/Q3qaM8Q+lTs7Y4v5+l0M5SQsRioTkr1maqSsp
bRKqyHNJydNWf5agSB+PPrdZLMAZRyPlBMLj88+XogThACx/w6nv8YGMxbG9I2Yyq54TIzNfPTbw
tz3NJwaz3xLRYjoZauOImeFCW4Ch06kGJlTB9SBjPfmIQAH6cf+syYVEwTqswqjs5T57xp6FjuGl
EoCqTNfPj/g2WWHe1wxDoZLPi5yJikya9ZMhCAULSKiFh6lBIpfQZgkPcVnBQ9P/+TTBXt9bS/5k
RXda1qbK/JW+76n6diEAzBiOnnemZ0O67vWaDpcntLet4+fAKOsXeRFL8pmsBjTqmIatPGYzv5pg
Pa1Rh6//LwgqhIgl1qHQ3ZAX+EsjZ2MSLl50Kk24j0yPgPIEdFs4leDonKIjDR74Hp2ijIDVZ4Bp
F8C3DBLx2No46gAetj7r7rsiSzWzgNqMzblZTN3hvFNfD4vepk7YYB1FSEJdEFnXC6+fuvEBxSMq
2CtOq+V/OVML+P3H0F5qz/LmwcBnbU+gVkWOiTPUmJUF3/hvDFQkSog6n0nEAi+ROe4uu2HPlb9Q
VtpHwbcHtpfi4P1DVwkjE3/wbeHtEDVb0nVnJXWObo9UYLCfUleWzhGZRn5ZNWiiQpG8mXvK7BVc
op2SykHOFvo6eWXJe6K8U/nWhSccbuA+ilxn8AWDJPfhQZlig7qt9q464SRKcTK+ZuTuPHwVo2gN
hrWqR2TASrlWQpTHRK6LGILyLwCeSTl/8oLnpGhjRwDzF5Ndtxu5um3YePEwJzujVvlvdcxBkBIi
jOBcy3HrOCdCeeerOMlrhZ0FRZuC49z2LIP4UtIgcE9n5Ggr49oSg34ixR8zKg1BN5URwSca95ad
CPubLHd9BgNnfXUeWsrDfgaL6oWe0Arx8CCI+cvkS3b0FfW0d1S+XBf5zldnC2rq63KRm5vmGls+
aKd12S31jEPW1zyRp/ZpXsXsUSnPW7cs4/IN5VfEgE54522RLvtVNVUgik2R2WxxIQuVh0aMsvpV
SGhTDAhEK6YzCTwviJrAEva1sFo6WusUYEbl75FFb0sxUSB31BCCKn4EUwfZPvW7e+f9UPH3L0uh
h4bIJ+6i1rCQ2guGCikiq+/Sw5+mlVjiozLANmsqyCE3VWIVlazDN9ji6zilblGbayWpXa6iBE1z
7VYgbGraGyjlSRRVTU3sbAM59bxiLcZuctjWHt138JKwpJjTNQKxu8aCWpGR29RVAWs+JVGATe0P
hsqqPJhlkw2lkSRT6WwOhiVEvXcmdFiNKh1dE6LOQrDMp094RSJCfJNmDLj9kbFOrQBrIb3gOhBt
v7RjYjiUDgiytpfahDi0W2rvJXtaUcJXTarBumpWsrXdNAd8+fD3clJ/5DpE/FiQ4KWa+bXWTasV
kpecLxizQFFM9PpJf0+X/6Fbv41hdFFI5o2FrJN2myrG4l/U7dDSlRZau2zaRI68FkNHbCmsrSDp
vNlt+iAbs9h/7p8rpZteutovkWHiwEavM8EEfYPjeYe+/He1nGViXfg0koa89VXqkujGvo/PHUKr
Yo3Hu7JwSBTEty7+15/yklx3rofMvrYAmL7qEi3HiMDtF/AZhQCKUSNUEq1rM5q5+7yfB/aG32bY
EcR3B7GXAvIRyhKHHRvOX2JkH5U/oc1u7W10uqmOk1SeWtjuPykZF/6fnkaomiiv+dR9FbFIS6jZ
DF6rXdQMwnyHpyruIlo3N1G65oJHm116gImiTJn70xkgB2/0Sl0c0lD00iDKpMjybJ45pz06+rFF
grwYaMqL4w/3n0/g2t4z50V7rZXuvcc1divALIqAxtzSHVx8RDX/nxzHFf9ECszHQtxTYX15jKDv
SFKAghE/a2vgToBfq0i7XA4oQZO24GcNDcUXtLnutQTks0zVbBrP05q73ujXwicuqiPUmkD90stR
VtBUQt3dhNAMDXNGxnDCJIrKwL8F1ifBhhION0D7EDRAFLght9Vo4aUrWLUcYAv23pxMUUWd6pWC
UEd5yZBGjB3l1fWW85PfvEyDPvx03h65pvLvJkaP169rvGljeDnwNtT4vkVDkxFgAB1Bza3h8alJ
2jZmSKBC3tHqL4/zHN5KihI9QdHJCJWARG6Jc/ZpHJIim9wRzC/lrM7gQY/oPuxL6qWezCLbyF33
7pDEfaJ30D2bDUc1CCpj6qt+Z8AA52TldE5yVcfJQ2MLTiBNctrU/ZMZ/IBRuTfMU8gKd4C6KcgA
vpXdqEe52b+9GinPmeAl5T0UOSsVJZlZGCUY+j/oifh38BmKcnY4ErSYHJmG3Sh/IXl0wfCgvHPe
6WTacqmGtxUDQATyDRDX6M+TN9ePl8FLn7lipt33KW4RwUpAj9CUC2QNMrTkHHGjrjoVY9dUZZta
Q+sfSVf/rSL0SmGyClEsAnt/Za4Au2ClW2MVoWKxvSMjQBwFRKkEqkfeAuXiF1ePh3ufTPEqF98K
g9r6xcoNfZQBDd6j0OW/1lNRjCMQkFd4SLG9eV9sF9rCHmzR4spMwDx9Pbcyxx3Ib0/QuW6eKJuV
dJIGXSsjzBgkkxuhZV1+w01BwJbZhsF0NUYSBowENZq+PZpsZdGQYVJDzPsGlPgYC2BohiFBfksv
bL2WxVkTkR5/jl35zbeUfmtTaswPH+2A2cR6QzssCGA/OFv5guY7HHFtzEWzMkVVWYttJB3omzPT
wubH0Al4iKcydpGuNdeV0qT7F42VNOdwMjqKlIozeBdlwzwgaBj3xdieVwT+SbQARzvm6G/KBmdi
uHmM4J5qQ2IGQIVH4v+61THEbPc2dDTnWwyJzi9OLBBxR8AaoLrNKbanoq2KvFjBsOx1xsQ6W49c
FSCF4axLd8D0oPWLXHxqrtjQk/FXTjW6CMMAFf6yS1l/ZOsf6druVuF8wnEioKtIUBAEK1Ndzvcf
zZIffg4XCM3CV33f09zpPy4fUQDeSOrfnUouXcohoK9a+G5tC8TGB1rfHrsKrPLkSQ9YKOQOYVCe
PXYQBQAHFDoTeVgO8EpUd19JzekGQfnkkvqlib/eg2kS42X1YIRNMOgWoGSVy2vOyauRiXX+jqll
jxC/C3ZoS2L6YWg31NbS8xku7tHeWTfo0fg+ik6MQe6KK+CSQ8txa7x65Pn3+7HQVcOYyF7cEEoW
nsui775FwXamv5XFk7oBza74InXOA2QPNtDluRgtnMQ57KpSFs6iV9NrvlhQHml2TK2pb3GyIDoJ
WLnJUM1tUJOlYPQqhz7MVxVgl20weoEJPBZ7mQDFWP5gQ50Qoarp6LQsJ4EtpdiudavehVDzvnG2
Jlhnk9BNzvpMxm9D5HDb878xUYytGxcj7LHh4PWUlvazjvcG38EXZ5cihxplQaLeo3Gxfbzw/Hvt
kXVw4qmbOSX5IBUcJmpovJAeBRYpLr/ya37nvEqilAtYeNjYFPITKf+x4194C6kW5zxxxbJEGWRI
4Mvs/AckTwEhUBjv1MCk76u6oD/9eAJZY2kcQtfZzIzShzyDXDY0AGovKjFxWqjaGjqCngON1b3w
Y/64X6edWGrwMWNdDKiTn8bsS4jc4nVOqGbjag3puw1/EA6RD7KYGSdnHpvbeXWQSDy+4T0XiBHZ
1djrrsWOLSxdxwsVHfg/+VDqTeNhKjg8VXrHA6juWEf2ZDWf26xoFLRCAvJ6W6g8zXSxNVZfY1hr
YYFvdLhP1eQyxMPxdFRFQu8PNbJ5ya49BiOUEzEtFMUWKOMvjDou+YHTcm5+9UahVamY/Bx/PFUs
sylJQgV7oCjhvtQgIVgS0L7MVr1sjOLrZSWrsOvRYE4CG5owCAnEd76s8iBgrQ8JDPcd7f8JXWCz
eJ60BIbl3XQqiCV0nsbrFGUl5Q490Ygl87NuWE+s5Oell0zcDJm9fpenHGekArV4fae0XngTPYG/
ewGXfORMXOxsgjg3ghxTg2whubkxQ8T/V8/V0kKCleZeXGdPdZppF9PNEZfcMpJiHa/rNVYIsXjP
azLzrqB21enPeOJDNk/tBFGyLxN9D6kbDuwNnm7Qw0ZXEHcMKz8vo4iRfxznkjAEMLO330kOIUOo
DvFLXL0V9o1g1TdHLNPOMu5NiO8ILLzr2AkwJySw4T3DhY2XEN8pCo6n0DxNjMJ5DSi1cJPEPh65
81Fsb2mFzByjZThif4X8RJTv5I8O+n0bN7xsdJ6bpoCI0d1USd9qidGvEQ78w1pG3fw6nB7s18hY
w0bsO4MQOFBNtgL2e4ztJhQ23FISIqLDjwIS/51jfn94svp1AljerjPRoZHu70/g37jm45Td5AmH
Qpza47UYegCWbfv/XeCRhllILCtUDh6htuPsS7NtbW9P61GDMDXueAHDWQcowRfzeMY8CmOrxFU9
p+UhLI5XXerreoZZSTXmdjDMGG86yKyYgbTYBsFsMnBEHQCI8k6lrF0PSF7dF+WZxjyJuDN5+8gr
EMNVJ18Gn5vXkOhRRaV9CRI1ZBK2a5OMIxPBkRqUV1Q59vVUG28eolc8E9wIXFmpVLxeeW/mYFLA
8bQAmqYdFBngRESDKUH1qPT9TmtdBGQNpKhJszvBYdljNkKezszE3LLHlY263hGk983u//F2nE0T
n7CraDDSeQvuQ2oNQMmfXb0VGrM0Kfk+BLDJ0PNzRXfYksn4CdJo5EndaG1CnLpZrbOAWnQ+cVhW
6f/oSr0Yqw0/KI8hJ64mCuEXW3eMkrkyooDMNmELXYP3kSe3OI2oh2KwvlQlTJBHIST9u7vj05Y3
5+t4iso26K4iAxL2Dp2mqgWhhCPEx3fgfz2wtgt34yhYFAJDzvPr8cTTfqHpVDIEtGAEOrYSu4oU
K6jXSoUzodtG3nd2loD/kNFong5falm/O2iurlpXRkii+odXsa/UbGfqOBaorQIQYX3DrgU6RqU3
G52zfINkP2NQCXWItIBsLVp9GbgitPn/FuOgy9hq59t0JBo4hEf5Cac/YrcAA98gAycRQY6ZKS/2
Vu7YaQFVvGa50ZHwszAPbcYdrrbTiH8T1Z5oSeAuRMcTNkEWqmXblZ5+7jNRlU9jcqw9+tJV0PsC
khOUbAb59raqrO5i+bVTLYgD6x+i0sAPedGfE9F3c08d1rEXtDKEGGMIZBFLU2ABCSwAeNqNOYCz
bXTophaGP9lNjF9oyOmM9PTFIfdVsxkyZxTTb+BOJaCaZ5sKxnJxfSL2HXEoFdARt77HTIdX1WtL
Waf+SkZWzvWhrJhVWnj4oXebcDizrZYuKF+UQrdX+ZGk8LEePKfbZfXRn1Zo8FrFZoHtYjPuzphX
RT+2ghV7WrV58XRcmjPYNNkUzjjWsiuojBDOGgASfCo7UalHmTdvaw5FO99vaI08iJNVtpMawieQ
sDcJR07l02Z00B7rTRyEINsZ3AygvzxYMRHlft57WVpZKBFWcVa1shuHuMnQjxpf9363RoMO1Hpd
cQ87uFVQE7I0IlfjuxTuCIOgotBQPESN5a37+/3qxQNhVQicoM+Va0OV79O4aOVJJWeSYVjqRz4F
Us8lOTe2tiV1K4XtZfA3uGPi102W/DA3B1ocnxvCEU5hmdz5K2boTklTa3bNgEp4faUU9t1AQxyd
EIeAVSRnbmoc1IoXcVLX8qMchMcx7ZtnDxQuD2Qa0tBkIoD/N7E2+5bHRcUjoXLSdhk0jl23u1cs
Fuj60vaoCzxWD/x5uztHqqkeQs/PU7YWPgneoXHMMw3cFq/9emiVnwObwOG79TZD5a7hM5pbmJv4
e1nl049EvzAvXR50Ku/Ca2UXosVxMe9nDPZlwj08ewCtHyg3Ier1ocgC0jLh0gmIpHb6elzcQV6/
he9+UJ16Xj3lE/z/Hr5mbwrk96wtLfmU5pbuIJz+AHBm7W7eSH2jjW/GYC0KFGbys6xOb+v11gsa
MBZyhULAPfhh588dMSaBFSX/EXX1qGUaQPYLv/WXoacXJcRVARbJJ8W+svyLt2ov9h3YTy+OGE32
CWmTCT8g41XL9gnzFeCiy3/QzGboWfpRVyCgvP3+IyEnDR/+d3SwriFKPaojUtGZldNZ6e22/yFN
MqmsPdEnLyc4sR5H2mVOfRwoK72nYmoAuO8AOxlHoUGqHFiRNkt/czUKgCMpnxK8L3w5cjs3ky26
NmU2SBSeU6FJl/sS4Dk9R6rPT6UneV6k4JsBslY9vezkzDYLri2FDT+VYw2cxTO/i7kGsqi6V5gk
+hwPyo3oL0k4n3vac2lWRXnHdOOBbICE99x0yjAhRPWsY863S7bctAU21KqdM0qPTCCvBOBcviZw
2kIJ/aJVYZe5O2l9qr2TnGpuhY93lHzBhMHrPuZkQfqiERV6OSaYKaaLzN25Jd09qFTELbSbHU9/
t/+/y65KpSBM7SGnadWR5hBP0cdTjpv+7gdxl/bIvD7Gg9/Z89aHPLsSPVTW3pwM+62jhjIHQh+i
qf6eNZjZjMGFK1i5XU0IR5vKPGhRwnwCQvC66fuquOtS0RujPfQFuCvFtLEZCUJuRKZ7IBOBc0SK
lCTVzhoZdQ8mgOzSW+l0xrLu79SWurHtPA9O+q6heFI58XDNgZ9scTgfjv2NmqR9lOnlKpnAuS7k
Ap4F4sLN9V8bQdsMc6aUy9GrMCk8rQKC09hMdRO2RMPKcEorO2jFOI9z9Sg8E63MEtdlh+/4D5uR
8oRwDn6UEQRMQGMqq9UCQOm+MMB6l9+Df80Em4Dd2ksuBXoWIV3qJ5zEihe+hiO7WToYcj+z6R+j
UT3eQBoB+5hBZICZdD9rFQSNQcFNqTbCvf33TSTd0f/m/tqr/kEz0GhWSGaZZhn4f0aSXo/I2wOH
TX43mi+ddduUkkNqtkzBUKpem/ZK6yalgEv2zUZDBMn3+T6c0u6/1600zLwAzxGo+H91IqPlp+Sm
MF7V8Y7NZeMBEfbk2RcH4TW9AksBYCEO8b/+dKu+4tgE3DmXgGA1SU3Cf5MsK9zugtGKal6SP3DR
DKwqzWBYeBQ9APXzmC50TcdUHwUETLBvi43wx1s9zQfoyZ3XeX3MMxwom0DfUIUncfk1gHftac86
03g/cw1D+hmC0iXXQghjxc2FpXZ9PZMUAEY4t/HzdbXdVJ7GQLowBqJtKj5rPuwNbYOLQCsKCQ//
094uUIbwRSAwuSsJ5TYjeheLD2jJhenwsRrvE34QF4bggJbaJTI8zzTHgRd+hSksSCRmlSNfB/V7
xfHkw2r3cX9BYgr58lu0mI+Tp3yaIstLUQ9YHQggYma7rWrXQzEKNkr8wMzUlv8HvuQdF2hZaPaH
IPW3pVUlV/DtWBJZ7Cs9K+CIeMkgEjTBegVNS17oBxbqFaZC4vSNOPHFbeeik28wyQ1Ff+Z4rdMt
1y0iyem/DJO6Ql3HLiMxRv5sx0l0Abcu9kxv4nw1H9Ml8sQa46s69VcstB/r8izmbLUbqxHvbtoB
yGWkeZBT0Y2oiNJyNFG/6T26L7OGNWWk2zUEewIwjsGgB2DGZb8j5sMWt6+OuSvZU5pxi3ck9cJL
nljDiyeH/ktZ3LKb25JBRQMbURwfvn+D7p5tDAqfjqDVoa0mGzfNESUET9cX6r86Zz8WQqnYkHIv
IteWtPlUd+AJTG3ZOUfwBLL+AVbdG+gsC96RURuoE7IKC3YgtC6ypZHa11iglIliz92zzC8EXfYz
+7NfFSncvsGYUYSguhVlMDML6Ubc1MzHKh1D5weImsIk1E2tr8AXlJyM9JpCizVT+esVWbLjzDRv
mO9uUn7ykxET06tK8l2JfWwauwGsdYIi/KqwtCGv6iY0qWup+wY6DJIjjf/jp112r90TYXLzz1sv
ymaxX6CJgKaF0CBrilXfLIUdklE8P/dukeSj6X8FAxNLaiCoNV2i++dRFv2Va/1A3qyBZealt0YM
aL8VFiK9tHLlCYym5wjrb9l+LrC0gAxeUzE/w8OgoREjLHLDnQdDyBtGghrlLlFpzAgtQJm+q71S
+PXQ3RYpZuT2WZFfPwgRorpXmdjyJiVAkcqoG9dfr/DhKnAHxAvbiqfP0ioEvv/y/JeOO5uPzFZo
gR5WSmn38/H1XlLYQtfjUwgWRQR02DZLK4ad9wU6/MylWE2KjA8cZN5lVhpNzmqoo8tfstjWFapb
SiTUk3QsOAMj8omJBIEstDZ6L1w1Oes+jmmxAbo6MQZusE4fU9V4ZQ6CXVRW430sFoZs865WhKxr
FV0WnOIv+ndrMInasgkbWZ7gGZqelSg4bcQ8KZUhrGUdBo6HS1U4lpek7IK1f3k0UmGfdCq5dKEw
MLju5fVVh3g/oHIPbpGe9ZjXXCJrTXTn8yh0BssvKoHqWYPLPjnwnvWV5VgnGohQOF0jL0yBvIoX
oe1ch144NK2C7GHVT4UwMgZWr5g2CeaJhafEqkFe1nudo5gUOs5FqPoUEFOQSPmt9wk97ijNqUKT
nZDVRS47lUzWCcLG17mo4l+6VJSx0zIA1+DEJsWeECNuqjXjOI4BQfqAkyiKAyzNrSWTrZmJSbMi
gT0rR8p78fF9jpzkL3BeOe3NbsZiQW0iXmW3rh6Iktnyfta51DXlrrQrn2y1DMFThjooMf3Kg5tZ
T9Ts2TBtdOixTm9DBrI2P4CQINn9cH/13S1mlsrEJ/DCg+uMw+5BoHQG6qaNxnIOUiPcqHLHJk8z
Qy+584gXqCDhkV9jGx/8TgQqK2Vxu2c29L7ZZW0YGu7a47+Z/CJ56/KBaOD+L3cjDfS0iwmvUMAI
2zv6M2LYIyiIhimQ8m1aMcZLPgblGvFne4Cua5cdnElerkPptIuicu+VzpDY1GVK2zpcdz+ROQNg
pcaJ6fhIl7OKWLhlQOG0en3DPsGhHpA7qU+o0YFK0sb4xDSpTRkEbjTRiRfxEkCko8jBPg9Ha7RW
4wWtXpiRmClbdazNe1F2keUHe6WOw2rOkgA6AeHSU8sNNlEQTm4FIZVf2O75FE3jJUhLDbvDXHW0
AXpv+dx8UY1VGDnb0JRoKO9kLdQmdOKlCb0D2KriAlWVOYfbFIrTYfoF7eoUm3L/r0ETOg3aAwBV
0R0HGU5FRWyHXqQCVd/MahxiWWvQiko0Bb7fQBJ8bPTkzLtEuQ2CCfR5+p+hkXOBRjqhw5fyOwZ2
eQaMpgKLsL2XXelqPkfJ8qLEZEZLud0Psi4gXFvRAM8YxHm1iajRQ/6zenJ7SBR3biCWR91R3uFE
A4JYCsjdZfykUhZMnAXr4xfQz9vD82BLxRFa3CrTzJYzAvlz3vyyk0XFVQ5Omjz7/9ywlCtuKSmG
yoInPbOghG8054qCieZ0Scz5HrYXvS/o+jLLxr+LCVV8Kc721v2KTYhr0JjY8+MBtgDAvOt2CQw4
Uci/S+MOrJh7J8e775RY/bVw+7bOlHdMBZpyxxORHZdzpPxY2+5/zNPlRASCc6N9ltxydhdGn/7y
PvZrq2Et5CXF+W4jXAIdC916RWiEJo7eU1z+6J2kbrAZnbnmGrp58gOcbOv7yEASqVEpuIWNm5Ct
8Uc9/afjNpEC0Vmml4MAJw3DzrSQCe5XGfms6r6qO8uQTddRfL5fmRBIeRUb11bjWwlRGra3hWIt
oLkiGDDCY73ZToARoVLeShAWyO/bn1gMqcBKP98JdKaNhqzlDWPs31KEibuAmEf/ls/TslYJTe9m
OWKDYHXBVXkf3wRwefBsjLLYmz0PMLptSq7V45u784hVQz6ydAX+WXC4KgB2vdwGHmjg99WHn3XD
SprW/M/u/vF61HHmIRpayOyOrjZDswOydwQsRXRGx4Is9GrIzG/XiQ9kf630SNZfYK2Frz0Rc8X/
G57fLuqeNvg0bBtIqXm2H3M1E65lxefmt/4KaALRT4FoOX77ikpbV9DBFMboFF8hESPThSm0+Vxv
s9RDsMd47y1XBPGDLdQKIbENijjv+lSyWBZb9NMHgh5rgTKfTWq6TBPi3K4zPMPBsrkne2l5Psgi
qt3TTPS7omML/p3MjbV3kmuoWIg5yyLzUVl8a7muTHNM+Ephdz17anNWW9SEJe4TaCcjMczccRDa
Shd3Qyr5bzBbmkNVIzul0EVq1QPSrlAp4mfFYjlbZ4ujmT3mWvShwTdV8WpW7oNa6muIcSohFbnT
qQf5ABTN4YPUA7POk+e+1o+/+9xO4c4xIXjuYVNI3+3CSsTIR2u5aFVTvODNaa6wHa2fEIiBK+/1
xjQCvFKuuFK3JDcRYxgHmmy11EcJ9VJpJ8AAx9cTQxIZibxU62ial1UAq62NgRyeCginwtD3fbwy
l/ELrcWd4dLhKv9QOuKaM8XcpAQ3Wc8sUP5M/wMXyrsDrs1Qlyc2WBUB2eS98oNxMTaDQDVRyGAh
5iop7omhctIjNkPwKACjKmf1689LAoE8d/DXdSfHOrxhOWs7tlD8aCc613TNnTVwbmiiayrezCsI
w6sdM1o5gpJkgpJdLHRKxlXKDUZHkxjutVG5JU7oy+9FYQ4vSrDjNrML/BnUwsaKRGiWjcQqRARF
1VHBbVusrr+9x2gZsFfbZ84LIGsdSvOru4vbs+nwzvDAGLouMLBrN1O4b6v2EBFLxX9pLKuCn60F
pcsLQ0a64RNyu2oPxXE516y73bS+A1sxId5sItxBSLdRPOlIXR6kQIk0yByAlz650Zjd3qOqNFTd
ZkHK7Cde27n47oKv6RtXR4KWGD/0LKL1qKDPF1qFFeSp7+dcyGdIvzvJcgHMCJyFexdNtcg70w9b
WpzITeqANFkklnhsBneXzPcb3BrI9JHv7gJk2ZTLLWNO7P8wPAPV//Lsg0kiKMIPhe6rqV5beIAl
rQkqMJQYBbB/vt7iNNW9UhcqoHVgoJElvLkH/LRS8VvLMP4iJ6HcH/puV2mFtSE1vXh3J481m/MW
bi1QnLx5fwWYKYe3DCR4qzMxIJ81O+WK9Ul7WyheCdWQw6nhuz38DJJmQl9AZGd6R4afkXh+jn2C
nDsm7rggu+7LghSGKLbpdlPnfBaySRbyRr76feZQg8RRmHzwwGYvFtmU2a6ez8nIzBOY2+4PwTP/
4mjbSM0bFZriJPg8dfSzunNGZsq98EBTCxdVHwKDeNrhuABip3wWMOA62RYVW/pczRoqX/DDSpbu
Tv/VqvCRYwPz3QRE++uPyVFes35z53WE7n2a8vfsJHKuuODXrUkoJEG4hpRUc/46sqNULkPVxpl4
bwOFsk5g/Y4nT4BU4ArSiUzOgRUV1X1Bq3LKT2+C9UNaRCLXSe03UJdwk011ja4A/WEBWLg4+XBD
0nPfvi+uM+aKtQDcsF8mW8Aecr+LBaE9B0Om9EHdu/KWgngZIzXfQoqGjbGPgAxhMNsxwPiM8vcL
bHHntIgE2WiObvjnHW8hNwdDy5Hd/Eptw2mqVB5PuqXaHk2G3lF//wR71OhIjL/Qy0ZlKhhYyCdG
Smq1L5DS33JldIUNhx1IwsN+ChGMXd9oD0CmXfwbPnwPIRfdDX8ufS/gg8G3YI6dMFeMSacR2aSP
fETHstFmjBc5T3ILGbBFbIl3UiXhPRDPWXFD4pvJ0BMdEFX21n5vhFrJBCUQEPFgEgPnqbuE0YpN
g56if8FBS65tLr9FpE4P0OMkf3OMm4RxCnIyoVZmFvSh9EeVvezPp0x0V2/74TXFViFM3LITrSIT
w0ISWOV+FXsVQMAnX0VXZLDws/07A8P84J7PACe9HQM56+P4vR9AhTqXLhRWeNgsG8bozbVIy/no
KeD1z+Bkz3NWzQofn+Eq+g1aJGQ40BoLS+wqQXVdV0nMYia+H/+zkCqYGHAimEre8Twukqx/YOcY
eBY8gs6a3HghwKw4JHlahsbs7swMW3T93/lsszfRVrVXXdvAcTaCsQiOnQu32LYVrdi8fIzBCdsR
unoaOZtwzSYb44gyt/QW41R57tC1nK2B78+BTkKFa2wz++zLhSqvdx/jLo+uxMrSEDZ5hEcy/vOL
2fx9XZrZvwtKZXnInUOCCD0/xnag5oz/ZDta1YngosW1kyAxaYZu7Lq2MEi33WXnC2r0x8dSDcQA
Xz/DvG942PQJv1ltztySUhdabr68wbW4yNw1N+f0HuQcYo/l6VxqV8Zksj1tFSkl6Tl0yiFvGFHi
/CqYRdRHS3c5/YJ0qbyKIHeu9uoEObosOg+5iXP6ItLfGYFHLf3XyPObwCo+W9jfYKlk4wHY/mrx
x4wtH5cA8mW08w6txDhDo29/WN8uaWrV8I7Ce+siW68YJXxAPDjh0KkC53aRWvpuarOh/+lYLSKD
NbpsMX/8mYX8s57dy0ope5QgMfedTqBYsVl1QM0EN2l1PIW3JlnEzlLMZo0CMI2jR4Mf5lBprNxl
MrfOXONMBbSufcXA9NOHqvU5O4fMIqQduK5YPo01BkPs+o44+S83iuLoObgOOnpESQXqPSVcmbXT
NTmGfVgzE3Np3gritWWA20eQhDyywjD0GTeiECfGRg9GYvOfbCEmcE/uf7HeNnj6YxQfqiZtJKbp
vFpuY7gd/FEhysT3YsbrsPJ2qbPfY9SbGj+rKKIx+HqjJICqlJMew48yHZ5anlFgHt9K6Qygp3JA
hoEXTQk2MDUriJRPMmXdwtZVb2fqC86bwnnlEWGSAVJ/OKeVjKZ0GzGZ9l66F59ZazvwDGJKIf4q
x0nVhFLp4D53tbjTuEaICFwibsE/wmEfoFHKhbaZa8VOp+pMS2M9S33og2h49WTNkntHqpeo3F5W
sg4q6txQCBshZbb1mgI/90l+hkopEafLb+9GuqjxK2yv9mWX1Npw9K7ADW55wal9uaptkd4SnMBZ
8R4gQzLWiPbAsRC2aSdppF+AMsrPdGzSUy1VMzxjIykpX90PrwE2fAgOXVnd/vd4XjxEmtZSCHT3
CZqhnmxmhCuA4OAZm+A+m6CfhBLNDdf4+OC46Py0VsmU36HYwQKJgGQOkC+NXwjDfJzvEZ4WaDTq
+2Y9z07xTugF9uiybRIMAaZsJdKRYGpHgEqEptkPefdejqJyhuyQZ8NpjhMdnPkdDIrK8hGkkQ+O
HvPH3cJBWJiP3bKfFzWaeFmpQjUHFfggyV2ixCNGDkJArq1FylIbI8wS0CHuaHtq4Oc3p+Updohy
GT9vZwqEpGQDsWG/9nobJDyHDNaAKSZean8aFjeYAJyfG/HEr7v+A3hrA30qgjFBjgsC370aYjtA
ZCKZiaYYEsud+Hc3Et33W0cVoJG3j7Qv+pWKYVHUyU8zK/l9H3x6PyEBkOegdUHiJVPGa+azPI/X
1p89ZsCfCDlr1G9tn5ZGf+jAtEQe0aMEx+amn+gtDyXdSWj/DsvvbFNeeDLqe64AqT551TSUb8gM
vet4ryfbBd5w7jvccR1hC+dnoaWPVPRYwfLtrxP09Mw3Twf2/PQfap7QyH+yl90JV9xupmg7fPdc
mGTLDImF4nUd2oWhevJDzxUXxSvnatD+BT8ipLMb6ruUuvQ5IrUzEqUfnGblOHYITdXh/LxRxchV
JCAXKE8aSLJkL+pNig6y2ifhqBE5U3KISUbeyCyMlK6WCaixK2iuNXT94b+uQFDs7wqTiVfPttJf
gnHOWWD3EKNtAOpLEd0EJIYCQS64Mt1xdmbyiTAdT7rVVW+fDbmn8/rBtRdgpJA8EvgGqkjky8QR
5ObdHJI5vYCqZt2UGmm7KOQzF0kbusYySItCcMMWDKnS7DqFBHUNe1UmddX1KjHDEDfJPPTtQ85o
jE35gE0qOh8eUepMJTMdWPQcxaEM/4LTZaumi2TRGwG7vP/vE8qWQ5hX4XlL+S1wDfiYZBHa1qaT
7KGPpjMDPs9vYM8veWJqHWOolNjT7xe5LRwHuOWAb6knmqO+kCp/K4So3C2y7RBynhwHtISe5syL
j+l/JnRMAbvF+QUkK+2uNfVGu0Nn9ChjrkdgIyP6ImLutNnX3e9+BM1xJaOdVgG6XekBvJun9UqP
r2P4pt5tvCNhwJzT6K23PAyDAHuWpVQL05UUR5mXSpaZoJxyfTyrQosPa5vmlY8QMUFkuUafR+tc
qIPQbuh398ISb8YvjhUXKFWE7R3Vzogze3vPGwVk2eEJPD0LBa9hh7AYRC2tA52524uFoBuQmWoy
ChrM0USNpO/OepqLrG/45A6KOI9Nmbmvv8ydeY/fkiMlBk/FVVMWEZtrjYUVX9FZ974XRvg/Rnce
sGMVRw0jN2NxENQrjqDAeM5mZy5v4MLErOFNqzK6lU4G6+aUNKA0POhFTWw7DwVCc/xcRgn8BxhV
Tsp2GDgOrCUuVOmBfvsex7D5Z5G0CsYeSYCteyjPw5O/bV8IoTja8i06wGJRlO0+Et9LNgEAjrCX
/xbuMZzLuAUOfnJW6tTg5MWROrnbjiBJfjE+QgEgTR4Es5qBliIUmIP3+MIr1rq7PO/+C0/e3FXB
GWj8Qa9ex9FEFmst7vxiSd0rLXkU7LCulXwY1siTfW2p1UgYWsRzGVsrYCitCPkDwsYiwtxAUPzJ
J3vtplvIey+Nu4DJm7KpwMPujcaxUVGYb5r7K8FrF35SDWukNvjE5s5MW2Bza0QtZlrJvw1UHy8q
dw/Qs3H3KkD8vjzzVGVJXWfo5yE6V/sxZOjBL1pnyE4UbYFGF21QR3L3vNXd69rd9iIaKGUPdbtV
DBNWNnpGiLje/GK43qsWN2rqf1nnHeeKHR4RjLntVY6vWXl065thnIthnca844F+EVLljps1jrQE
5Y50XRFPvMaT7VKXD4MwG6LG/5BjvC8h9RmrshHgRSq5RcLV2eVW+AbrKqRtOX/Gil00kjj4i5z4
oF64ve0wfqpzqjual0YlSapLyEwMy9XZIIxjdbOHkZXtACyuDjOaTxBhm75hbRoZCRBAYffhpwUy
9of5HFI1VkN8go906pFHXNqF4ZbpaLD1AaZ2iXuUUTlitgoaJ4/FNQOpS00jODRC+B0R9SeH56oX
S5QN/Ld+UL3TBjqtZzEKydoC3Ue7IqmgwL1iowHhSvA++GjEHdfJG/hWYnvqSYoWQ1nI9OlUb1Fj
Zho6axW3sMqRg9rUZRDkzILdIRGujcX2OwSMHaeYTcsufDWCHjkvRO9Jxogg7dU5QOvnrcajpi70
E2dwH0ijh3Nr/w0z+m4SaSiPi+tGXJUrOGdVjWNNHuAj18pXFxM1cuSftbnvLTyv4R1eMR1VnnCw
eQclm+NX3IXCwyZIigM2nl6POhQ+rOvNUnpGCHoGJ4I9mB1QByGK0YEh2XUcbkoBZGHtSbcFcDPa
R7yaQNIOmidEPW4IcKq8UDSxfRPv0pM2EyI8O0fKQkNPns9RL/Dp+GJaOmY7p76fN4fpFQD2PxHp
/T4BAr1h/WmD6nXUDkGD5cMPHAl45qUYsXJrwjBJCcwIgMd+IGCetZY9vcUvNrpwogcys6FJpVqT
S+tvLD6J8KpsX3f8YVb135WwSWP3iWMaI+Dq3ADaOlh/kPgY0xysLYVdTuMv+USHNThnswSuKl13
iPf3+fGC2L7N3+J0EZ/ICg7GHh4OKqe59M3Pxv7bDCSJ8b4CJLeBIgjfH9w3Hb90pLADYvgpkdGm
s+9CXSGOtw1i6zM13XYTelXybjo4vYRt31pmNOsCnyuDbPFA9cnU1a2A2X2ET+GugDqVIdRUqejx
pbw2ArlebQwHf98v/DkVcCFw/cakcFD9OggaQ6eE3ZXIgCjp/PdAeOEyIq50qEzT1NeYiUDu10gh
1EOqTCUhapWkekVm3lCR1o4lBrU08wkYws0kYyVZ02WZhu9/WUqZ86+e4iDzdPJ53uFH2m6KOsjo
1kUMEzXxQAxDpOFx5ADoU4TPyxoubCpDitdzcyAskGQ9PnDfFjarKii83QtRGoi1MQiG/ZNO3Fkw
lZZxfFSds3HhV7q+VGLOM7tqVzQYKWbzKjpAecMk/FUGBzEnN0bqnnlgi92uqNqhXdYZn94phwWj
DqdfTb/xh9eDI4+U2iDuv/jrgqmw1O8L+nBAfaa85EX3BxEsLXt6coagFwpMj3ypwdNnPSjFl2dC
7K8guh5Qwkhx4+gY8fkkmh/lojPIxywszvU8rMbFdOjaSC5u8PVmARY/Bkup6c9hLwZ6oxMvao/3
Xq0gAmfVX6x5SK6F3VK3fy74xmAYiBWiKB2tSXOsRx4lq0xRYiCU+6EBNqjxE51Ot5gtXShb9R3H
b1CNHiiibGGo11UnG20p3ofBs5xrYkCKEAgQBNKrd+cboH1mSAcKvWI/fnidLPURf0KL4x2tOhvx
P7LZtKG4aprdlShhM2qzABs/Nj1NTGoGp4cHIgIjinSsRSnRhxoAxHDVszinFGAHoW1wdU20NGO2
wPgYzL5pTUnyyYbkqQ+C3A4SfxC3SvYJ+QfEyjNGNMv4mqyprBcK449ocSaZsITwKHPpN/cOK8s+
Mi2N9DsQUkjprfPyUxY9h0Bn9TAOEQT07CbW5eQEMhuHocHZBmXu9JHuO4hCXJ5xouP1YkQBWzKy
C49OFGCuiQ88tEfHv/6s8puK6baXOQOhJHwTPlsFrAKJS10lNz/c91a9ckyiNJjeQ0Kk3ihweFiU
mCLPtEGeaOpAk2b72+vkRKOywZKpsqE9BGkT2zXTBsP6IO3RmS/ioFep+THJMtfH1jRO7ZSq3+OM
5Qmj27GanY6QyhwR8TVw/S1xWaZbJsZ0jBrb/wFNYWZDXapRAbxvf5fwg0MN9ELbz8BgpiHw9m2k
7TP7/uFNVTTGkq43hbrgyAEUkmPd8NFf2sdISdgu/QYmsXjuk54AvSe6yHGmvd662iHerSMfySOB
CsTkqPxbaZhKL7NyJOIJLsE/1eYetMPiPg6Yq1645ZVa6Pc6nemh8sO8Aa4okmB/eHT2NU9wmGMx
D9ZYUKrEESboo5UvOVKYQHBfBZwMiPeDBQzOf74YWEK9PUSFFXhRQMMhaG8SbJesmftfB99tEhxQ
+DJ472AAjgNsdOTjs8zTHIKMlWT8HlCvrGoUTTG8xD5RptIa1LYjfzqVn5TXtChMnA2qnSA/b/OC
CvBNvgflzSCrkRY/PartkP28n6KBDAqynB/XSxO8XTjwcqlT7P9zikWUwMMBJ0f2xhYLFgrrNv2l
FpNopNrzZn5YdXHawuXYeOndXV3ZSpJl97EvHuzJGPcvLw3YDNvRqBJvTmJbcxQpKxBMq7fafEFe
Cb9aAOgnQLWvglwouCoR6wjiuMvkghRCeFyXOwvJIsGrbFTtgsjnzjrMtuf0z/JKVMXQrfEZtQEu
d9u2jIX6ThYgn1eR2tpsp09xtPr2AjDSaMt20CuDcTLBf8EC2qEnmS+0UGJmB/o/M7YjUI4eZTl+
fQFJ8ZTxv95+zctf1LOfdzU5tELcp6PXgbN3E0dvpkmYOGL5+XzJqJQ7qxLL5iOLVEpyBUII5gBX
i/t2Z8CqArzMMGrxM9UqsLguyDI3eF8y9LRRtbD4rBSnodvglgDM8Ty0+mKHw2IIrSQ5uaQOMRhU
6nn7gEjMK2a7dsI7+FQcpVP9AYE9iYA3TJY5eX3MXuoddbFAN4v37hVHxeCM8sEs1WuSDYk0icLK
zcMO/wI6TiwDoCMDaeonzkcjeFYv095GJ3YGTZ3QgL2B6xHpIH8fJA7r5wZAaKlxQknN7/XPpytF
Orw3YCXn7UHEH3wycRhsu9u1KaHY+RMseSKv6s/9IbdtTQx9gyJyt321+PxLCCxHDx5xixm6G4sh
kgPKOJgjQ7s9DTiWimRSx/dMSjEYOgCOMJeJcZ5iGM8B0vlDfihd8GO7Q+cacIWkaMx3+YqGQSmV
wCmyXH6abbX5nEQ8FsT+PHdYaLfa0mMQbS+Y/KT0hl25ugJgXuWjSAnoBUymu05WOMZupj2aVC0W
E/If5ndYNAnD7+yhKcPpzP2lap4y8+INh5hMNw+Co5OHVmyQLlz2AhB2/ZVFfVsnbpKpi7A9/z4e
KwmBUXo+83O1ArCfjpzISZnwSB+ciu085QF24ozJBytdIZsGPOxsAqX2suf8KSHNawaFgW8HoMXl
HWVyfwNXaWx+SQVKavfqFKYLMR31LK2CzPIfHnnMlcIh6asKTw7LBucbOkh/2x+D7wnRj7LXtU/e
HXOR2Qe8QaH2DKDG4sYQBtsdhDda6WJ1R71blZ7w8ctlK2Mkh+XZEJyKBlU69n/WplQRgVTRNDMV
KfpWA8/CUIl7wXAqt+xUarvpevhvPVr1Dkk48UVBh/sxXdDz/MV0YzanlQmHI83jzXIg3xpT7/BT
Q95ofR6hMqhX0l5RXsZ8Ynpo3qtwb2ap8F/r1Cj+ptdsFxcZeGKJ2u7S0uYDIz8DJKvEZ4DJHdVz
Feb3B9MkVPMg1XOJxrYOLxe4hvg0SSkhr03stzwOY/Hs2W0+/XkyFl02RZVd6soODFWxkD1oktOT
72m7C9gfoR13FpDNZMwzU59DPsnNOcZgNCgWcysJi8RC+v9t6t8TN3vunbnCsN5MDVDmVMHpJanW
aRAX4XF93Eh93SPtTE97pqHP2EmFzSmj1OteiKDMev7cDUGa7UafBvio9vELO0eLpDwWT0VcjBZc
+vmowFX3Vsb/OYBobK0MEZ6DUqTO9ngzwVtjrW7FzfGrirEVXaQCOK3/SXr2Lhh7JsyTpXX0f1v7
dZNhzfW0yu3dI0k0mTr/vhiEMt+Pa+HIBQr02wZXgNkhGQZQN86EJD6Dc9ywfycuJLo5SLYSzwQi
qlYO5nQPtVtjMvQ5HesQbHfs4rXgnXmhi/p2fp+qm7FxLbD0n6B9gPK3wuJ+ArNwqX9yl6HYQrb7
imjbVldepwNVpboR5fIrwpSutgaXZ9GzvpTUSw7s1FTxktzcscvTYdmC6xaARPBE2bVSPvfVmAau
SluZ2p3XpCtOmynJuH6mm2So46gRAkPRWVofWr6+jFQPqYwe6LaGompCKJccYfQaObiS6Yp8zR8t
tZ5q6Ic7mo1yR1/KEXEtqCSo0wmicsJr1t9+csq9ASFy3P6fGhDJ5SXloE7ojpME7rKB10tzkNei
ZJW42EzFqB5k2j998HdqiDR1DnQNYFKSJNqAoS0b4oSUiNewLdtZhZjNtvN0Ih5GG+idr0mTXm37
R3+gw+9W/aAUtG5jcHIbtfN2XfQK0dwXzo2BSpHtfXbraIpP2HqFAGbVodq6cW1OpNUpm67QGVxF
TFjHiLA7vmHKy8Cp6DMtMQnYBRKVrig5ZuYJu44DcP1VXCK46i3JxqYP8eoVdiwA6vbaenKhveEK
oKC2PIopt+ktnxWysxDCE3Vd1XbYe5XDkYkUyXY/sTjh2/X52yi9nh+CIhIqqDZGEuPg9NQ1V6Gs
ZnnOPfN00Dm74FwAkUA69UNLDHKUpqaBDdIlWgKOoQTTuBEkbRiuvSVNN3gEJq02yCKJCwINP6G3
WM8yK3yWCDCL6p7X78wrU4xo4sz170EFN/B61icMt/10tZPmNoNGfyInCV+uQfGlWwxLfZBTGnsy
PULEt6DjkPz8lZiGk+3SxPHuUxF7qHJZmWylg9VtBcXtbzlOiAxc+yDOXZH7g4EKXVCKcmkkm1kA
QxmlWJJIrXxqGy1gu8kofznAy0POyt721ljvEJ+YxQhvwNkpou3Na6M3hcspFKSjyUvab6loPA1v
pI4hHLl/1Db87tyFvTRJGNmPVkkYhgryhJat5E+ShFVt4CEz+wHt660nuqcZ0fLgsfW3qe3w2vhT
EkfDp52QR9h47rAtRhGJM2UUsAWPExBG/3z9s7A8eV1FMbhGy0g2QnQbLQV46nteIhE3mN4ZSb8V
pnwKVxsjuNcvmTRsbxDC1MzOV6n3wdefPJfNbrU3efgOoPVjv3PEiCYHOEG0g5zGLS++H/EahSV7
i6UyMiIYpnD/WIUubEd+Y3i7DVzkiIRVN5aMvViebOLMSNOQx6rF7XYHsEST+QWVIyLLUF2wHUf8
IjoV5B76B79/cRMlJBgeTQFe/C3TGB8MIxd0LRFy6YXPK8sDMoz7xcTvmuDfvdTcBP8e1srbhQXS
UKsdHlgHAvtdjoARZOkCRFXi5QYoeprVeBgdYwBIs1EjFrRAIabYoNARo6C+35mGSQO/RLnh3fXJ
AN228aJQ+qgqcG7EDl+pXkU2SmygiXasybK9CXHDvskVcee7oI9kIpBQNOh7W/79IFJiqAC9fypf
3GSPAL5m3b1bIs451p8QOFgn0zB1o1iL/XKwHuVLAtIMccq8F50oWd6l1C1oaDzdWLzPPLNJ1128
NSzxJIvjhidwZbKCRtbHyG4Dxfpw9ukprUuKN9xho+CqQgwIiKN1mGxZMhF+igVthtY8xbhrnPQB
Mn79/SdwPJLFFkJRwDuFRPQZeJIUN8gv7cL2Oc7Vux90n7DeRi7/ePzlzR9wuIqLE9YjuK+Mbj2F
sqnUGyBdIkhk+1rS8L1CjCtrjbrhyFc50WQT6naH097fALAaV+ol/hn7T6auaT1hnLQTUtECVuqc
f56crp+lcQJs4cmJkKXObcGnQaOHdQDXM1mwHkFdmTjDkgW2mCsb3N1enYe3ObhNPFiJr5UbNBzS
/m/zLq+Tbv29n9e/bMGUEen2Nma+edajH6gypiEXb8/DF0U2G7bIj0z0rLOQBYEOdlSE9qZ2CJhZ
uM6Y9+KkpIA8nk05tPXWHBpUPL+IUC1b1PFw8bq0iS0A6fd+ONZhOMQVYWocAjfH+/kcZhpseDAD
8iQH/tbKkxinumLOwSWhpvalDkl38sOgf1kfgHC3fAvvZwIxDl7r9UdoKHqiyCf/FpCTn7lFxQ7/
HXpzWKLYyKujoFa7qNCGo/fK/4fdVRvLXS+3xyNMDVdd5xWnnLfFkUPMiQUXjQWWaW26s9+f/PFC
Z0S/fxM/dvbnoap85l/g/DU3q+8ZrxfKfPDmNM+8G9cibJ5HB0ZGC0oSIvKJxWrZQGDTjJjJrei0
nxeMxRJVSdy+TYDAxUuwvHWNIQ64lEWxB8qJ4uFVajHKfE9IPioWCZYFMiVmdyzEs/NNQT/XVX29
KSC8I+CyLvY+DlNvY8o64IRgcuYpMTm37IfZN2rEcTgUEQcSI/QfTZ6wJ5JpX8quoNuRRXJWBkBO
rGTbXNRONmS7a0MaT2+hqPu8IYtwiy0kfJlk0ibXlWAI0uu+L5Td8u5vB+9a8MhlhwMdM2SRWaJ6
BwtlcBmqtX58lZDZ7ZVlIdbLi3RA1/jJXY0fAo+sbHwrVSlTdvYm9/ixtdQEfWmYgB6WuZEZnPbM
rgNDDHYkxgvo+wq/YSWi8YtAmyrChLwDACTn2V4OdJNIrFfnrc3dNDs9abo2ET9PPl+whneFGxy4
/0pIjXsnFVP1Wl0CaGofxp391c8I86Skji3Vzf4qtp+1Bzb20GBr6WkUfPrxhI5xnyPOUqddaRRP
gaP16moS7PEaqWEIlqtRddxV6/ss9gIT3EHiamXacQkvSINVGGfmKIhLlTRLrcFdJmXOHnnwJBjN
JVTezV5br0CfQM+Uz7AZCMUueWe+Dx8Q6+yPlkuEkDWIufmdX1GaaH4pNhOFzB++/JvfCwvJ6OQ/
Wg48BFEzTcdHt+X1j/WlqRijzWeHpHfsdUDVlPtWq1U4GNvvMKx3UI3S6N0FsSWL413lj+Av7v4j
xBq4scGo/hniFl1zTeVNtPXz8ozKwc3W8Ji2Xm1gSKe8tRMtAfrNHOLh137s4+oKKo2cD9m58bNQ
BnXlLzEZupSZnwOIxdiiKaiIb5zb8Fs4kyoTsL0lQCqHOUYs2GLIzpGJoU6VdOX/RN2WjzbtlCbY
bNmCFEIomsNTWbXLcArX5GUqhMtb4OgGkycxcnTkkYhISc5Ng6BwL6Df0Mld7NPXVFAC2F720Mpm
djARKSc/la/+wRpHPwmbWAbVFLW0UHBCc726AiObt7ImUN/kzN8eZf9cAbqNeccivAY9ntuqWCrY
6+pgEnxcbJvX86bucf7wxre4hVuemhY/8gGqAqt8R3t9RI2ubgvgFxcNFBcJvrIgXFKYXFV3atBp
V1nH8b2n9GE1oP/o9NBlTDzcaTPyGqg3zfGs96O6uQdXUtx4N5dTX0911/llVrsYGSmjoFecwf+W
U0C3PF7LIvSj3VdGhjEneYViaAwwIisC697L19bhEcOkE54HMN5gTIXcBHFcglijutLrnW6J+i4Y
GSP1RDUBsCc3Ay/5fCtizWUgu1Drj6XGnAIJk3Cjqng6BMr4esesZrFGeWWWov8C+0uHmNT3/mTl
gkpH+/RbcjmD54RjeQuZj+DjJudpK5GvJX71UctX/5fag3KSasS0LzqTIpl73oFWdox/ihGo8j6j
/5FYEiXB/6c8HU2c1cPkjou8NIVzjrNYBKDemrBZd/l4/UN6Zc6Quex1YGGS6nqYj8t11Fq8qDk6
kkY2j7kuaV6g7CtaRCRsUe6fDHfRMMGyx/ojj0JodhMgFwMRNDDHUpfIwXpifNK27oil1A4ozQyG
4vqUnBXRfTkkym458uOgTiidATsBngRLCORxPydVtcHIQuAxxYsKs/Awb0WqKbIZpBvCz8D8ZKeW
EKGVE/iywIFInb6Cb1HwgImE0zc/JUBPT/IsUiIl64qGeq7j/LgUI6QgxO/v4Ep6lRav3AF3S//E
8SEC4/gtT5eyrayQnBOnXZYgP2reuF1zXZaGWzXejaMj4roiSPi+ljOx3nXGKckKEbDetMnNXQ7I
M42aYx/Szaj6yNFG/kDkLdZNrqBrDQpHlQlWzepTyAOR8jp30eLJ5VdW+FhhbFDhr+yKv9wy4Euk
SOIuZsdV/p/SIgBPECurBdgNhiFLwATvFOlggr/CjOlp0Engek7dwUiT44iclSD9Rn1ztdXsi6X6
FWE9bMizYpifL8ubO51krMsA2H8nQZ5F6rSMo6ITXaiY1LlpkY/6hNypEEnVeipOot2hvKLgKWX9
CyK+588+XBsCY54fMOoQkKGc81zwwuxgoksulyEV5QmTZTi199sPsrycZsggRpV8PNlkCF6yjR/M
hEMBwMZER00xU+VuMSH8Wv/ERxTTaqnMrnt1Jc64kby61jy9fczuj0uoFMfRI46SU/3LEzeZ/P2G
8pfc1oBxo2woV+CfF5jULWWwdLhcYwrJUsb0qVcK6Qv+wZ3KIoxvQG6pbffHKVYUJEWGwBoBzNJ4
WjLvaOerjczr48SOj+srtUofVuKXaVbP3zh9VAc13SykyVQQmXE9fl6hMomxOAR8kO5gRYMRwPwB
J9b8n6um0Tmct3yMklXodo5nk5M+FFeOXixA2QHS59kOoXh6DfselzTiqI3nJJK8cpWS4dYCHEPW
bfma2bQUSfGFNbp+T/vAnzuuSeLgcWla2+8d6xQqtiQ2D10vzym1OquBueglv6yMnoDOmYN45fN7
pGrsRXu1kEUGRNEUT+rY80I6hK/qif6lORq3NZ5eAu7xF4ciEfxMNKrCsgCc7PBPBffMXfwYtIog
qGEDCYFh1JqUJglqkzgfHeVvpcuRNX0c2aJmSlVUTX+XVZ89IquhX28ysUPPw2u4hIpOuxCYaXor
k15Nw6vz1fEuZq96WilnhQVmg4EIzlVYzAf5moDBZCum1UbKR4HUdbIyP6rhkGjU5scEEGuTfwFr
EYYUoQhoZHBVAheoJT2PJVid29wYI/01GYh8BYjiCcA7vU7+Lo/yrXI2EELzp7ik8hLl+DH4E+kv
A9X1ve5o/VdjQnJojcMevJnc6IB1RFwaRD0/KvPtBGe0AJ/XuGCCkhqAs3yg7F79Ldzx59BPMTfD
AxA1ZKCPeLnszMpfjBt1XodZSkvu7DLBQeGcxDh0pFE88mXjCZwiRlNsFCs27u/+wMagh5kOv9L0
qmMNJ8dTy0Ud4X17U2zL9jC7mAuuutjddy2X4kSibJ+1H6fOKstGQfWLOwLE/vmRPgjKNMfXO6kW
VTqxy3iYOF726Vd0Y917h0mbi+b4WRsS52qsXdmJI+RyOgGZSC0+/nSe44piB+jFR5n+b8KvOeR2
pP24A8ul0kkDndg2xeflr4N15TvaYO/LtjLcuNyNgBBdTLCzzAIm+62IX/MDDjcfnkxK1fjx7ndi
3vLwXXegFMuV5zoxU7fBwxWEeknz/rkoG/2YwTv1oZksUzVihbPA9n1QOK6AxTPG7rWLBSbAo3IS
tn3+lyUJuz18OD8q1dGi+bsC280sSsLT1qbFxeDscf8eVZmKLixZtst50X+DM6TCxYma4Nuixdvg
tvPA7pmfS9H4bmxILBiQwkkjwwZ+1zU16yiphTKzFoeY0n9SDGdmJq7FlTBAhjWWfRnq1dSXEawB
URVl2YFTzOiDJRSNPgdljr0kzwiWD3PkGu64XVCokbRXtGJiWgRSCAYaOqq+r5l5oq50OJXRJK64
iUkCOaEWocq6W4bIQXhYvlyYw6QnvTIemxP3OcnqxPCpLcoLY8+cmmwPkLqRWNBeiM42CpqKXxOF
g8JpmZ2xwLJsCMkxsnzOR5jRpvLCelLIACuEliu9wxHuQpJgKqjDvdnGtE+SgeTrvkQqVo2v7qqw
bb3ZVEQlmgD4LrQkuZmwGfV6fsgQ6IDhZBN1vFuQDgyBD8xX5oYCXHH08GOf99JjuBUWc1lJ3NQk
k8nXC4KNhBm5Li66RDCB4ilRkGmPXM0LNDjSRL5MGx3eESMYdVcCjX1wa8YmTACY8CqGYabLNi5I
KFvT66aCVNHlAr1dj026HSzrBbeREh7oS+GKzN0jO7NQpGQzUHa394tXhqiwaVpQTYtg0tM79nBZ
MxXjTOLwQLggs3vv12dI3wuXvCx0U3B9sWdjUYU4OHRU5I4uHl3k5VLRPMeWh7nJ4Wf6yH8zUuWe
Qm7FN6edlWYkfDGqNjh3kCO0C0KfayPekHSDY8JntEAGdCGoXn7feXilLyODKPEJUun8QzBQhVYL
5VGUgKoov8FcKR37ERemVF1lT7YNv4ssDkfrKtjlHD4NWhGCX6pvfbGoNg6gzJ8Ofueqi0HL+DPD
pQ2ZtqaKpxIfZArTsht7eFAVemx7PPchj62gORWR+jfm1KgiT9UBFa4WPiryXnz7KW8cKvpTzXT2
4m21qh6heyffVH99LHfsaYTf90JInFiFugshc8X0AxKKQCA5i+6JBNUQ21lm+rzruC0PRku7W7DX
Xu4EK6V73G6+uSnNWqew5zKyxYDpDSfWn0H5513zhUQPQcodMv92RJGwwsHNf3PJL8K/AHzvDYU+
ntpg/tIRO7PtGAVJimFdzcc5O4w4PsQKGz8xXJhRm0xihleDeye+9BiHzgufsMgNZV140V8lbcLM
cYApWvpN8+/UIVExXuHnbHW7GzyJTvSNw+mEYq4NhzaESBj32RKQvYj68VtKGFQWlPZZ8bpkhcyI
VCI1O8Q5VnPrOMAe8kXgsQp3iT4ElhUaj/PlsPJxGrkDovkGOO8ygiu3324p4sllGyKz/+h6ikUU
Bets+AI6Pg5az0MEGw1DcSWaiJSBJFMqkGkiF5TuWoukfEiINSO9ifQ2CJYk+EmrnMcwCXR5kkZ1
NDyFLTt/IhCJbCh84WMhzAoS8DtFzLjHc5dp+tSkhr2Y91w1bkzV2giU0sBXIJLFPHp6niownKcK
elkL/d6bBoefdXb2WCAVJQBeCfr59KDfbDF9TTlhtAjBOG1s4KO6hww+r5wZmienxl0y935YqEyp
U6G1L2SkX5UpMeMlFIe06p89Cpy5/YpqSeNlolhk0VbXu9khOeN9ZVBFwEwW9eADJcj0yKaw2zyK
bnvSvD2KsYrL5S4YBwsIQ8RrRPqCII9wzsNkwtHFQVoLSpv6gA9jzD1a5oglyekHQHvfWC5vOfUR
eOVFL5MrE0WvrEw7+Fcw47V5LVlwv11/6FVC4A8TrhL2F07JiOg9m7PNBoHHGhyThn9oKzA0ISks
LkJ27gswUs+oy7VxKZWp7dAD9ATJErpKPGlvW18RGtiT1cgKfbvg/eNS4PxIyGN6Eg4FkbL3fzEu
XzhzNow/yWlj+VHsinQ7csEoOrWbL2vUEbbbDG2c4mjRfi0YBi7z8OxH4Uo0hGHG/mKGSjCzjLvB
a0CdviSov4Bih4OpZGF+yyZWGFdvvV4cP7QH5z6GNIDBSEQvQYs1acNyAPUX24jN/n4yGo9kRmw6
oCrlywDPe2hwzHgSBq4X+9hp8z6oa56lBsPROAE/LYtmqfJUFAKChC+lqioqT5Cvs9Nettzg80tK
VJvAeT8zBLpeghAJwOE4U4OFK3PgyUWElIRqAFE8RurcwTtyE5DBUFYD5zhgvXJh+fZ96swv+aWo
YhhFBkO6xiYb9B1yZ2sOLrfGSRx+/X0RoMDfsOB7+8S84AOzj6ne1Jd88GW/SwF0q65l9GrIFJzn
3OtxrP05EQxfKnO/Q9JQOtR8ImN0ojwnWKA/auX1//uvuaeXTAlxQ906z56jBlAdME4g4NQcdzqy
O45FPdlSBIBy+D8cr0GMOUgUQOEtLcE5txRL9IcohYZwBLCBz5TY8Chluz5Kdz8NQnUrYAGEWYw1
ABD+Hs0V+XWfUvcdFRlu04ezAG/JyE6c6Lkaft7YWe9AvxMd8TJF20vrweViBTkOsxCQHtkuIfYw
I9upVmPMmvtCgqEAVjE5po69wjcwZLjKr4GA/sRmco78h9EtSbjolL6V9txFoCgyXoNyVBC4+X6F
QM3nPGCSbFq8aRFzRLegk+sUNtOGrvUMMPjyrimqdqS4czdeEOqk9N/B+R8TbXsIMDdVR6mfsv/a
t+ofQCRooZXC8Teri0pSahu/8+0Dfd/7HHX5wDjiE8iNisTHhX/WgwX7eopqukY6iORAtbxr3abg
HWBCfI2wpHeZh3CqLo57VS3Z1rkGyspKrqhlmeyB0TjqyxMOTPAq+rR8i0NuJouiCOqlh2fC8a++
tySASKH04zwLOv7qqm57XjXtEPwg8jy9pS0Cx61qAs+fHP5eKTBcN/gQ++F3Fpl/47Eoy7CUbcd+
oxq8yL66+lUL4eTTc/daWHkL8RRwUA391FpirmHSQ6xl6b03z7YqTv5EYyuXj5O+x3nWRjf3khpI
UJcgleC4nSgvY+DOWUgUS+4IrI1Dp33rjaa6tsn+I6yzti5Gf24VCuf5iFqP/lwF1GcUjgT8ninh
wUCnI7cYV3RNzsC+4lkwmoLl2/0FqO7Awdfz+g9YCCO45d3pa6aRRcs048eCZBebtYUpneDc60Bx
DTHOSgDXkazT3x2joRpbGjMqC/nb/UKs490XbaYEwWusvz7WNC1qFYYUAt1RlVuZobF4dcw1dO83
TTllHwFvubmDCJvLJwmIaaLia8aXyXdvHZt+ZnD/suKuH/IgMt2R5ySLp77rwUpQvIcOveq3t3yw
1xDgyDg6MUcLsoPS+4Ox5SRXz4g4OKOuqRHAEkXviblzTu78VNcQkXpEV9hfKfIxvRuxjAdDs3qG
tXq/zeD3Uz0sgXdUc9Q7+LoIFqsg/gInSMi96RW7T0uBjkeVTGC6bRDL3KkUgO3ljpLH7YkSU47x
VyPtWDFy0Tt6bgk9xEdVFEFXYab5OruDCysV4o/FbpKoVDzPpfWdij2X3Yl4UkbJbhvv/ejXbHhL
bKVFAItwP08r2s5c0oh/1DD/J7a8dFPxG6X8fCWoTaMWlluSj9p2mKUJ4HzOBvdOnwJAxSrHBHLP
UldIL7gHV1Sfpj1lek6rDF9lfyT7gVs0ssVIiq2OJ+qkuvh22DVnnX/WoXlgm48BXWNO2DUTvQc1
mN7VTtpBqQdkMfcWdTJRqpD5Hy1vN2rG2vtUsaRzSKsJAZQL4a2GNircQ1QREv/EffHiH47pHlhQ
2JS2IuVjrrCSVZpChAVorBpvKsaFYCDMPjhyLSXNWCYeAxeglACBZKsXfM/zbztSufSn0A6OiGA5
qAdMAksuym5o+kCF2zKiDWxJhEYm3JpNp3nd3v/Q+r/+SXB7o4rMsUz8yyKAgejAGzbw+pl3JWSw
UtmFYv1OGb+wDvSqpamPKBun0+4wL5x5CAuFr292eW4fQFX37StUos3FV9226Un6BNJK/Arnm+mv
ofFwQtvJY6vle8xFpxosSanKm7Nck4vHiCWv/MWQXBgusb5T/6NuKkwVYcRnwL6FRluflXNJgt+S
IZtIt+iqKtWLhhJz6l8BOT2QbnkD50XoeUi1aPfUnHjWsNFerTdV6sfwA3kmxUctVjUGJvPADgyr
/bvKiGdeRimGOz0/SUCCPYIkbjyNj2lSXhq8YMKX+DmdOraVfomYcA0YjmGojT4rLF8gizv2lYj2
XYXPcbrkRpUQBHtsquIyuLUhIb37N9iNHuaNy8f2KxxJ6icV52pY+Gs9GVd15erove/WiZldzxjL
801FdN3xRC7sPkUO2djFBbbdpKhGQI02p8SQiVWP7Uhs67TLyUM0WbQVbT0HV+vMJG1RqWfbCCnI
KWlZD1Ivyovniw5QixCKdydprnFQXdJ+56SC2882l06p8ddkKS08GZ48TYh1wouKwrfvv9TASGOj
7rXkjjMqrRIXp3LHMTH1lw5OGg5H0anA+mj1ZdNOBlDzjnaxWcPsIy3I+FgPkMfDwPEjF4hMcpZt
1FEj8ypOTvnAlp69JeYV65w7cy/rTVWzqFhUa9Da3HZ9V7SSJvwoTzd53DMwtzLyBJri4s3wgijX
NCLTvyKFkJ5VtpRq8/cY6EqZxO7GwnNvNOsXGIrnGmXG+qczrhH1YFfbJ5wwAsPvWt5WVHkGa+JT
Gp7UiFHx0nKtya+8X9y+sPkn/8HU3SSePUgJffDsnpAb6NfA6BIygNdwNPzMx7WzX3XKS4R6TD80
YB9FeCDIQKd46z6hW2QjAnBJrG/wNdjqx8IXQNUL6VUgmQ9h2eHY4e0ZALJQXl6mDmxiXxqeFfhr
qH4elWoClO9kzVfOijjURPuu3MOZl4t77/j9mPrAaO3beZxgJ7ziP63pZGq6TZgtc7bJnJTqjOcu
LUgKtrcTZ+eevbDaesmlMFjE5JLCmtR2LNXXMCF19UU9mMGkHH+ejZigLRKytw/HkvB+b5cBiHhB
wTC7OJVGbo6Y+L/ACdN326DLzR8f+++C8It3hFGOt7o0LK9hN22Kke3ZPMQikKsVIvkONvT6xqLO
GgvE5lGeqE4A5c+TeVRrPUgm1IxGOn62CVMBrPfc4rC58TZgmYR9pCiNZzfP3ytzuCJcOPRVHCbO
vO0LiwMC+fzWIGp+K5SnStcyusC3vtmtjyQi1QKtH4FDkZ1kO60u9cuNMhxZXUXEAePpGUFtsJHc
uILtQl1xeGJHDyKjZeWBQoTuauVjnTfVKty3pXJPWOUrWU6geayckoRU7OqapCfAmmTmXfyKweay
BJsBdo1Ls3r+hnnge3lUEwsa4LTRDvAtWaxaznlUYOWftE5C9MvjT4qHI9sFeSn5PcKJEUT3fz2J
OfmRzjSL5nFO/3KmUaqWl6pqnYWL4/OZUbF5FjIdQnz2kWHgcFqxJvApq7/A8tFcnD1UPn4BiljI
NuLc+Pj5Abtk4kcgr78j/M7lLM9KmiB6sYJcL1c5xqjdgxeJVTRXHRChJc1TUwr8CmPOIIGBt83L
nHZlIoiY5vbghh8HulEkihH0osE3q4hcosSS/Cc+v6JUjJ4/XtICp2KFN/qVbpWgXNn6DUh7G1ug
Dg0NVbslelF5yzcqz3feP8YbJ2Yp5y+eMH1I4T/Z7FppZPqy6M0YPeYONMtlCV61PAt4MQPkURcH
rfSNS+2zEdK0WtXy/cXlIWmIAmd4iQnvQVDYmwJm6e5OCtCTfrbOG7T0C8fnIghuZkVM0Eq4/dNu
V/lUwKfvVWPgOCelNiBTHLtTog+/uK+8doE0DcRsZtpHmKZCWh+MqWVR6iuub0ch47plCfRSsPw1
TJhRu91BDmuA+u9KXzZCfkRV9PZfEZVqQn4MMnID+slKCErLJ9pgs7Gl863MkF6poWalFwjGx9No
sEmRgCUEPfYiJkpLQwrgT/P3fPctGC1MOonHBCx0764BlDisMT8vqnUZbl/OBIk2sMaBvecyBxi6
EfdDUdOHCAVkKYUefH6r0Ic/hgtgqpwLeyQ0ZDGi82xFIZzke0xn4XwMKpiGnZNNsqMUw8uRHKQ3
JVzWw96GVz5pYgjzt8BL+aRhb1Hp8Po/ifVYzdpv36/E88HicMDexixuv0QoTp+HHpfrhJb1/pYu
US6f7D6iSzg4B2zOTuVaUb9QNvS8L4wvADUIDgQq0c1nqPxvJKDW9YEp7vjrmNe4HI5ePI495N2l
lu0/2K5M++HmLRJGhrk/WuvCyPIBz9j3R/AcErj+OrOH8vEL57TR5L6LzM9Zx9s8Qd+R/GOhmKvM
4VQVKU2j4jY7SFxVnHW+5DVF0Uy4BY6I0fhsVaPqT0tSGZsdeK7XDa116Y70WVGg8ctVr5zVysed
D4k9Vd69lVMj+IM5lHEpFYxFOSVM6dThi/a1Tk6zxt2jXphHdusWrxydKWsj6Kr2vo/Ko2V+uj15
G7vIfOBlEjIiPnNILw1Swgzyothuqe/U7kqkbWS0CtlbVGGF726lRHIcRIgTTaw8hyqZJzo8Ju3I
197sX2AE+yV1VTh4gJ6BoyAlQKueTYX6u4CePEAa8ObxKZpKlrnNBhGmb7M650VVwbJ7InHd4nxN
oVLad5UaOaanWiSF9eyGXeooDLE7iRC/cD6I6PkntpLAPtKGjuBl3sKsIpvWOAIVGz7eSwlwqJFY
iPOiVivJL0W/9B+QJoqYEYb81nGp0zko7YBg5piLgpMoc2G5xDNdXD4VIxdkFTlC8HWf9jvZJh3a
6+g4goMuo9gdj9CLmbmvcJyLlYA7o72ZegEGr4Xhyw3s4C5wEO9/VOopIXsJDAak52qSJ3+1LEe+
IsynPJrolFXlirqnIxjmDQPOB45MrSSiJATbau4aO0b9DYBVa3OaeSzS4yFPIhA+13aEWmi+Mb2y
zMWXjJGmpT9sJovnZolNcnC4byCuzb329C5Pflqf0eMGjPOU3Hfl0tB1wdm4Yzby7fKrfRBXGlaL
awCluu8rfBNYmyKJwVr0uk6CflyMYO/yzESVrkn8rUpvdfaC2BPmTttXINpFXJMw0QQNMeCQEVKd
g93DR14hNA8uKgOC6VP9qQQCq/EA0FPb7wegkS2Iq/6hWYk5hFq/Oz9BKbilCPNjcSU+ulAQG4yi
X7MdA0pLdenR+yI2Ac70VYGeimy7b7iab0nwI6U+5qsJreE/MCf5NP8s1Hzc861Xzt14tU+ut//O
eV9muh7j3YU4DeZ46+SkCmseemBHxZEtNn7ZZiLK+1J34wfmi3YY79jeQaUR5wcyL2yuRe3iV//4
RP9mQkpG9XWOa6Wu4tBAD8gCpu1OJpjU3GaO9mk0mkQ+wqVX+BO4KlHKsOCxQ4F6kfywYiUbgiDi
cV3pT38cBg5H2vdU8wv9anxDOmlctTsV137JFNXbDB3Ghmy7SKzYiIv/XywD9oYP4o/Om1VK10y5
7TFLqJCB5fMiipH7vVW887UKp+wgbElvSRkQcpK6ta3v4kAsymd9eIZ0rB3IqvjhE1DLc5tBwvit
ln6+qCZ9WgnIrPmv5MOaEX869aT4SywEWHgd1gGinOW+1MJP4A9/Q0Ak/6s9B6z2H5XTNd7+h7YW
LppocDR1Ph67ZIWnt8d182Uw8PW3mYHxGYFUCBlJNMoeHfpCPK48+Y3qxIq/ttMXOB1j0c/VAfUK
MHJMaZxF55oQX5ScnqVq3HeDF/9f3PiIGZIVn736Avb4Mt1Qs0TMwJsErRxS8GWNosBIgjSLHm4t
mJivUuSWmcUSmV/gClHC7Osq0qblgTB1L01J0n/GBMmgB1r7VUziIFqvMFMZyAaNu1S8lSnv6jYv
TLZSgImJkVsjugEypvlGkWUumEFzlJ91YKhwSBrey+7EslSte5mfAT0R0jWMRSwwQOQzKe/LU3K2
a5+cmkFOCIAKvirh625KnD2Sd2jLNKQ9LxAZTA+fU2QjFBjfMOOohbsIw13S0LmRWaywIn4cKEPL
dH+EE1Mzwq/IdYMXtYKKoY+bOVY8QhSDkG0slYvsh29rcmkOYtTZIgAvDZLZwRxJtjClakpvjEqp
sO6k8Pd562QWwixzK7/M+Qr5R2igSOhQ0Nfps3hYomA1BgQkBy23HMixOMwNVmlFJx1gmcyhZ98y
wUvhY/lJ7wCv3q6BaWTj//AN4kHIIRI/74MUKV/C7Oak02pRgCZN09RP3UYW6VRQ6URR71+VFNo9
d0E4zYwpU14RoSueRU0zmeuFNxEYHMMr17jMOZa5GEpRK5Mu/J71mUyYDQsGftU42HSfA81xsxlx
MDubKpntYqDGhmZisoTq67S21U6mshj09XHghH3JU9q/lYLe3vkY8hF8BQtBXkK9RZqASNTgvQ6N
S0h6Xi2iNUrOVG/tywJFRVv89Nnqh7f9Jcd54KeiGSRYxFZDjTMPJ5DqWDyWomLO+fnxt/MWRtux
9Fk15c+kJoukKbIC5eyfct0gnua6g3SSxP2NJxMc/smyhfxIfokP3D8Xv7ayPuJX+OA7NNLN9WOc
ctdFqGY+25+/7+uNaob6z9h+b+2FKgOXb0VGqecaDewNRFf3fpV/O1JFbRuvaXOakXQLIGoI4/gk
TRKAOk3nFoEk+RYXvf3sduAC6B+h+yxvMvSZ2w71kk21rZoRkxcZRoIy1TNuho/nRy7PymeyYiwC
KuPNDZYPcnRphvApWkeGWrGb6+TMkfHe0qKfs+u4EuaqpGmuO68hfsApvjrmLLmzpnDE6rQm2VwS
MHT8atkXwHr8WWueDJWFfrGzLohnjMAJoodzyrCyQXeJqeqYH4m9Ry7p6qwjYrafnsDyGNCSYnnp
Fm+sBQ5YuPq5PyYagNRtgBgTthBEmuHvxierNLU9YrrvrMT0bzIeufUhHkBDIOE8nAtBH3AFM3m+
yHjEl3AogvEQmLiBPfPWK4yn9eQWgIlm8lvBtTaq1GEroxiAe39nxoWROSaIHEef9ejqL40fmMsb
ktHYFad24yRogaZY1jraKcZtDXi9k3JjdqTx4g5inwcRcpa2cAHTMohbDOArtY8QZ3Mg9ly2vXq7
/ODuZI1zACRxGScGtEWdGTEQzBywvR3ShY+pMCesMrm4eKvtRXk6KF/XsDrVOsP8ri9hu4KID0Gf
I2exp/GbcPlvWU5+uLznuI2kBpOPXuGIzfE0RN7l0v5rsB9elV0p1fk7hBqRbIwaZ5EAKDtZBlLW
9/aE8OO3CmAsJY1j4dJ5JmBGnGkx9Bqj56+T16lbCoKjgYhP5aDjxtR/dgwy9HnLeDFeszMhga+N
iwZWHsFlgrAJ0URdF0NEqxQ4PRfPiNjUB3W1Puph9PH74xAu+iOf1tjTn8IquPz3i7HDU1sj8Vfv
7V6vjWuhtsvu6tg0/aXO5/DFyEutEwFiNB+PuC00Xr2e6+3c2ObRvUSBrFGh1Dxe02Ai/M7HRfZp
WNEo4ERX8xhH3rzL/WfEpWuiyoU5QfPzODKWOQx6kO+dRpMLTNo9JNveqp9k7WeIMvKLEERw/ORV
wQ7nl/0ONFldFHroe3nzFWUjweMAlwHaccDuQVJgTwVuBAIp05gVjWv8vzwnfx7XsXN6H1Vg7oek
V2U4njubXEjW9lN4TiaAqAmJ8JagF7oQB8PHGpleWFyAMT5FU6lrtdelPQvSY1fOjU2xfNCDIzjn
BrCwjAB6QpTb2Ebtuj0SmzYY+QIQmqyfZmDjUYMQicDpLEcUihFCWIa/fUp+mFH8AK8zsVFd7r6D
DuBybtDpp0z79rOjh2gdlP669XTSlmprlM88ungDELIAyREO8VzVCqAfM/LBpmyO/cybyeaYsuaM
of23OoVVjv31/kXQOG961pkLxLMK4hRL5Q/+9uiUjTKXmdOv+tPXhKtYu4ohc8MG9EjhAfp7zy7E
gv94b9B9KLw2IrOo0Xgrv97nT2UJn2NQDqRDm6G/VVqCMviGjZr90w8mMq1HsVhjQ9sRlDb+jphR
UEX4Wg2GtpIGOrSeCS7HT7ORGoDFlyGk0OVEf/m5vPKBsdHPjubuLlrz/CZxyDkWIR2WBZyROTXZ
fF1EhF7Esar1urlWy/+nZhBT0im4RLKL6hsW46gEV4RdCMlInrYjB6+1he0FSa7f5lL+aB74h+Uk
/c8vHRd+/Ykl/JNpfNhvvgTE2JN6lcBAu08B9hg8PQ86qwXsBJo9gLGre9or8JU+rIfvR3nlPM2G
L77vf7h3TTENd1Ld0v4bZsNMSVbE5rcV0clf5unAQPAxsim0/3yZt2V4t+Y2ie+tcBgSyn2P+mxZ
Gl7fMC1FWhluAYUoN+Iikj0VK5Ghw9PEb6L+EIf7fS2ZrrfzRd1qaHT2YZmItjGiMdmb1Jaa1s2d
aapTHUr5RdatcRRyYoRu4vbKY31DxTXkNAlkUG53HM/ixnHY6+1gHuutD23p/Tf2VlW5dazLqnWy
4Bli60SmUAIdj+KtL/BxDA8TESRvz3WAvvt9HmpQQT8fNjvKbj3MN84fxid9M6eKneR8V5+PgPiE
FiWi0NQnl9nswfrV1fevAlISDh3dCB/knCkFwxa6AEkTyykLlAdxVkgNDzDiPgcbthlu53dC27wn
Sw+//aega1/TE6Cm+W/fkP9YpQtKXEc0EuSqQ3qYhCXtak+1ma15wlOR6WVPrebvXp3loWi2Rqq+
6kjPSsNhhUtDpAUTkPPJvqs8QBH2fhdtciecT0vLtEmGuSkqjH/LdA1zLrtLbroaLvWAR5tH9+mN
2GDDYw5kphlnc45dNH8tJ2u2YQnBI2Okx4BjEjE7JQDaCUTMPp6JDspqXu0T6xiRuFeMBberSitc
6hKZ6HYoq+mx7x5v+B2ujN4rCjKERmj4W5R4rXpfhHV0AVFsQhhXNleVO2bXoKpbuyI5GwUZEO3H
HDXsznt97yBPIRrjy7PJeJ2nhtVENB4i6D6ATKriFZjxZenKhI86QcI1RNaV166ozUipqqBR7YmU
zo0xWlBSpkRqa9t4xsDL/C11rdzyE3CtjiwsyFPCEmTV5Tn45xgdSaGnHtdPAuePmfQSnXtZr2bW
CqCS5cx0+eT97KJgT3IA1rUKGXZ4lKgvlFnbm+DB4uYvafwZOqjG6iDYtyPAOsGBhssSEBXOnJlj
9bFHzWO2AGFM3/lSeutW9z51K1jKKoy1rQj3IeBi+AGf5FQym0RhgjeWN63LiI7tVfN4HcR+LpCZ
b5s70aCB0QbLvlK5ewjvELaKIg1jZiYFDFaETBt4DVhp2kxYUUupjMI4G8+DdemsDGD+dHvZq/DH
6Duu/Eurkawb88TCCZFJvsdEegbbtCeER/qUHzCNGA8Ja7DPqDyLAMtxWS5SomShW+OIxTmqcWeY
Cc8X93VEnSPJ92BMnqaHstScgHfiXJUDGwI7NWe5t+EP5bAl9XbVfzu8Q0EN9Aijrg7StYp5KHAL
uSR7oLg+0vxTfKMNhnPF+CgNPHIYyCBtS2idP0f/iz0X6IHPVnRofMKLUhQPJJWZRAdbODUXUtHb
U4TopfJ59tkKKD321Npq5VRyyP06Mda4ov1gATzLXgeWKk8XkfcP2HyfK56O8dgeawSLvNJxyy15
C1MaWgtVeR+/f3EKbFV9R8OULxAFYevoj3SCU6gglkxD2QEJDx531Sv93KGFnNEz7xoiwKnzIsyh
DdlEl6ZpMl4moT5tbufrtvaPPp3q7PEXYUGu5QzElPTjliyuj1IqAcIUR2FnAlQTVOK77ehDEuus
4nM1Ngk+gVa/2UJn8kpzysVBuKYpPmfXms2iE+UJ1HgAvCMUVq0jrFW6mpjRV8+gqOAjtkhZnmIi
JLY9kZCZ+rGuQtHHQwPLJneXuX5Wh35Eq45966lD2lqvAyxtAYwh5shJe3hxa2X/K1T1uGrPtRbg
5jKthMs+2si0G6SOtC8docwjFDaoW09M5KE0cb27VIj0mhFgpc/1qhGU4rwIfjTVN8szDqSHt5nY
SqB6onuSWwFGXqabaY4Ka1F5vGVCj0sM0bkoP1N85Y66kJHBJsH68yS3XoFejtYLKyoxaTJNsUAb
hUnaQL0QTyLbwY9ftbi5Urthm/GIld90kkD4fkabKAq05TrQh686IqzDGnyPTBcesv9WCZ3YP+nK
lpfUooetEwmfSohNBfW/LYi3SJ/McwVQstUwt0w6+HaHTirztLFLc5kubajHQFw6BKir1cvToygV
2FtUACngjQ4JJ3tnbUyaXF12JXYJ7QTODHkEz8SHxftrFN0y821slXWGoFUlxxyGHDOv7kREYnp6
9SqPiEGP03yBwX4pjEf4Uu8vq4l9m0gHxW6SL6FGdrDwTPKLsHx4+/pigZdpca2DRw+383aHTFYI
yX1cJdofMPyE+JzvJ1Y2/MJBVjBCdu7XqYW7xteiG+BKcES8OXvTA+lm9/Rm0PunHjrlGJUH1IJi
TqaiZ/6lFlczZeHioFI5dvdIFewVd54m8xz27WVpI3VLhpTCNZutCSBoikrJHB80BmptSWerP4ms
wV0jMaPOS34gqyyhkkvk/WinFWywG5WbE5ApjHMzT8m7G3mj/b3UawLJM+ascc+oVbLN4MPwO9/W
2ylYvj2MyO2UKv2e5R2A5nR28pb14tdV7+yCKUz3thQCHDXJ3Z3X9+QKyyhOPEa1GTuFNGslvKXJ
d3ntdEP0K/BfyAscJImgwXIKyRmYKLrv+XmvyhYQVZasCaiAScTmU/quO/k752LEoB0o4Nog1XqB
AiOesyZMfUe+UwbCHUfKgWOyL2UVbnHLCkhmoEdqKWAhK9QBxpjg3lB4IQNwsV8xuMlo/yl6hivE
A0UZS6zbslm3goYEnJw+qTUMqABAqoM9sOxgUtBDVSApT4lw7GU6pUdrAEfc/hWOsrGm3F4Is/EZ
hw+Yh2cep79KJVCrx7uUycLWTQHFzYdGi4bmbJBpVZzeGuqggZY6so4sWk0NFh5hLLs1dqgzwjtY
Wa1vMYTRKXOvjcGtSxS/HspoN0xzxX6Xqq1h/gJ+Vj7ogkUQ58hwMxh/YZ+1f9Pj1NPftHq02t1n
4zWMMSytRlcPhs37DDWpRf92P4CsIbsy++Qlw2oImdOIr2v21NEHJ+Bt4H5P4+W6J9TFiKdPVonJ
z3/3AndhlTcKGm0trtC7GrxFlXSEI4/7D+A+CHU7WkYcTmbn9Lb/iFZikyL7KZKAkhc4vqa9XbLq
68W9s8uPFBe+YwIQldvw5UIBj1BA0IW+0Z+teZqOlXczaU6tR+kln5yycPfoFlhricjsH9dBZQ5Q
gDxQ2IQZr4WpE49oXsOFohFa5WgCnPJvC+6t7HPBmTMwRjp3VI8ped4qcJ/Lyj+wr1ZJog1a4Zaa
/m1V3fV+4yggt5NHY5BkitU0RWsJnp4CW+6b9hqjmHZNezrfEghqVg7/2nWQJ31oGPRvbZDolU8/
gHDa62gruSGqD3/mIr7vrJ1rKgCElJ3pKMIadmapta+gsXuPtfP3kDYQ1BukRif6DLhAJ5H3BCO5
sza5rUd7TM5CExj7LhAzVeu1W5l96yz72L6tTf8fYbOHc1SajQkkUkimw2rY8vk/ym9bBCzERTA3
CZB2mAf4VqBryPqEcGEDr7NisCA8a0FLs3L7J0vh4BJ4MFzZiCyIE9Xccb1wFah6HjcyyCdhlQYY
DWiW+CfEwD8jSp6tLNaVj0ghSGQoypu7btZa75Yi5sl654gvhwgUoHC+izQZiqTh3MOXzAbI/IAZ
mhO+haygKXbF4u8ZXrl9lzyWHbf5tlTyverupYXpUgLvh1jhai3IUw2notFHgSKFJnMZx22+kAls
xAph9GkSwtzWGiFmpnmai13JmeSqx8DeQlvdfn+9jzXh4RQS6YSqb0vdkz2buSuA/mPUdUvfBmKL
T5RGhgGCU4nlpHbUQn3R4BPWHzUE7pQMN6cJ1XnIE3/iJPvcEjs0NuUH/3OdBF8lo3sktQ470YXw
Pu8b3ex2Ml8TkfjlmdoefXJQI/p0ysmzToUpAv8/oFXunOHp+Ajdh1nQ90hxDQIGdRUbEaMN7SQ9
14jVAoF+jPpVRX/Zutv+aZE3iITeV29IJi0YS/vKPBteEgkigVvlo+2p7dLRWWo+wnsGgcnbztgO
ux0gKroXE8eSgGXFf3yCgHat+Lqg52GBV5PVA40l+c2Ij8+izNHna+7bjczYlx/al2xNBfrIbCBz
+cKdmNFcYOpwkIRajKHO18upfOevc1dByA1uzoYaoM5ZHBLV8omAIKk5I77nxEddyF0XAkTh0g0P
0z2l5sfVCdd4SDBROCCgaMR6onR0hyqs0rXNd07U2uLZ4+blwXUhDEXqWqyDEQ+xaT0V2BsEPzhn
VfsvwnxDv6xjXuSvPi9j5cyg2v+N+Bcj56LpnqgD3XEr9MRJeTQQ8E7nXd6FkszsdWZ1fMz1ub/I
5pVS187nH/7sVxOEAuo7oXNj2bozIK9VxU+O+Fh/aZHKG62Mbcm/K5WYimi/d7uLZ5h+o7/4dcj/
Fmdkc32064AFVDhKJeBM9zmiz9V0gFhor4I+rASbPxPBvp9XyIy9sE9ABgo0rtKcEj7DcOKh+GML
lFKiMwkdFZqTN+WgfHGLv1bg0e9lNcflARBEYeSzkpYJBXq8rU9cB0vNvXWXvkAfo+mlgDGuY9Le
BuItno4TbrRo7l3KY+whkPsyAbZ0HIugu8zBowxJ41eGCQo8bDTIbGWceORwgsVQjqjmswEz1Elm
g38HkiNF0ojJd2LbHviwepymUgFW0JRnDm+lSW0HDr1ZZJB1BQFSevH94QrHFIftkdCALEMCfUOF
ocDkjEvQshYxxfHhXfyIPLIEt75z7QBR6UWOrJfuLcEbtROqsLY1Q+SEckQ42ZW+Rybh8GXufmqI
3CPuHfLtERtzaXETtRi5Ls6sYmjrajrBq1AsLSZXh6vkpNiRCeQdJqgoxc6PsX4OAMJ2m93c2nII
PSjAo1I9LIXA3de29/xX5kNNr6mYowhNm1cNE2DFVcPrMx7rGviOCax7wQNpzOcWYMPX5kT9Z4c/
OMAgpuk0LzM7sPdAMIf35g1uSSIzSwKYVCHyZBujuyk0fxLOG4C4HGKuu8dcIDqI9PyQAkySsHkB
gwEyBigRbLsM5ZY0DKsKIluowdTE8dyTRQXEqYR1HoQ5MpaVL0Iq04VAef31vkuY2rDQvTp1ujFV
xIt24IApsGvJiuqqSFryDnjv+iCOTZKJbnwsJ9HB+yBHHUoklXRyEz1v7TLGboHkClualhHPBoto
h/0MDNT2wk1IeY4gpyNqPrYueAUIIzUGWiZ7zI8NVpqUSg/Y8ZCeKVhbzxEKwaPbaxndoSHYkvti
T7VuGm82993U9D6zfaB4TTQRRV/8/FKNcjRaAWkwF2X+bWHJ3PwZDvZMK9xN3OvHMe6lfuS0TFAB
TqpgkxIbYx6+OcoVWwXL6VPDKvAlkZvjV71G7XdrKuaIad4uV/GoR0iau22QXHnBSlWCvUQoWWS9
VPPGnXUiWi5/rwVx/fAZD2HpA5RRY4xtJo8TFea8qLcfb96VtuUw/mmNpjkqy+vWJLoYWh5ax5ib
3hUIrdNbrfmsQqcCaT46AowYhD+SKZlzupWof+1jCngmjYh32h8HogTlCCYIHbvFpc6aHzjNc60u
HasAk4oGylfYOo91it4yXdwo+V2WQW5koTqw7a1qASf9qydXUrVI7wRNZxHRi/gdqDVFKL+3lK9L
vGH7xbtUjCb62Qu2oBDYVkDJc6VPgbF6cTpVziRo22pqpoFkYvQrJVE4h5X3KbOgKaoGD2H+yyYd
t9bZ/NuhakevCYlSWgdhA54jpWzkuaGhoF9GJOnN7tMQPX6fp6j62ZjIiZx4n29SFkelJGDngeo/
NdNr9nIZgYpzOHiHEM81V9G3gIqBb2HIEHElvSOzr8wdzQBzlCsksAMQuRWnlt0cg7LNDpufgDS6
rQtLLstevxHlKE6uX37Bor9UBCmGHC80Q7UjBiA2b8wUesiUXiAJPlve1XEPyuqUUdnYxAlsL/vD
F8brd1LLpapGqVEEe1sLN84NjMz8EriwAAiMK3IHodwM1sDWCmg5Us/9ETOvauLfqaQzQZBCRCgu
eO5Nue4U9TeZEDIybjTIp83E/UEJZqDcwYRSURpmoIXMcZNSuJWNIR0VNZC8QdrIdRGmGEZfq+kr
JZOsFEpy8kd+dBLTqOIHdkLtjKU4pv4Vpm8a86OykA0TgIVbtaUQbvPWFFL9MZkR0Yv4BpZkJ5vW
1V4qZqHdMZ0DVxs6CnORiC0F/N3lXhRReYZ2c4gRCW92gq0rBWtxz5NXG28i1svXokw9uxR31+qs
wpX9unBykpoCHdmIxSLCJnYJIBOr9n1mJufbP7RD4mSLjJ/ckKh9Splg9Jx2f2LYFRd8dDIAR1p0
D96dxY31U+QWO/XCE4bct7vpZw/DNkzhLI9S816AatYQfd8CpEbU6jRK3JiDyj4/2mztsugBSurx
IWC4K6BhyI85qgM6kDx8DLigKwsk1MoFS6Fns1PFXmBb+A9traM4wgxxY1F230qjjVvQ7ITPu1xf
U0bIFx2EFf4Y6uoH9AYuzMTVQPkBwS1JnX/zrl/F4e0lMGySrrZvc/q5lkTyce2hvQGK8zRhdqXT
8M5BlGFnDzvf14n00MOtHVMSAX9CmitBJ6Y6Stdnjp68Bfjl22W97U5bodBE0IZLHAqgvhO4OPj3
G7Y2WotzVF4vldMdkus+cBKiiqOqmX7bgLd/SseoD0gQSgyZpdz9ds3rTzEVsq/pM9WUYIfCnkpT
fsVTyUByKUEXu9nwCiugQ6ZXMW9thj+KR76xC9Kh6I3+5NrGsHdNnINMiuLQYP1na4EEPjwtrlvy
1RvR6rezFw+LD7T3uw4vjgamzDHEE4g5GOZ8YQLkwPQXE6TilF4BTfDwcOvt9yc6hehiT1Mg//Nn
Hu2OFjE4BbMu78gPpdvZm5Lw23svQ9K6O6srbe9mfLFyhOfJRHbni0+wmZz9SS+C8OBvSAs1HDQ7
8fFkAGCYT31fG+8zJth0I6SFZvSjQwDk99IjuZVi8OtuxqQ0vDRnTcLNeBJXTlVpHrzio89NoZ6m
b5gljfAX4WSwyzdoluMdB7KKK85BhvZBXvMZZB9DIoyj/b2YSv1VVpz+8sidIkCeu+WI2gPqLxM1
PWyd2HxQGuSKF2J6w0k25VeNPPIyzQQhjxCmRxsg83i8rVkBnacOzBnfRivFAMSiEBycScM4inE+
2IMcpiMft5ciabhQaU92RdMz1pVDJDC8aXAJ2kqB/tXPvRvyruGi3KvAM0URNObnrkiZYH310+fI
H80hGnLo6xHbmn/wTZn7KkyTIVJP6KOPT7mtWTKpE2bqXzFfX9kut5aWJBwO3ijaoRSmRPsVOQm6
kSfDyv+Z5UdOS9DA0/vyvIADaXBxfVf+M7mPA0GB0WZtse7kBkTKUCHMFeTPLA81ZEPcI7HzAbGe
lc/IgARb9ChOGTIHjxokZL+EYXojQ7xfRGYawvK8ZqZZ30aA3/iiE90c2Wle5GsUzhfVrWOeiZX3
eGd0jUxow6O2JlAhvuq4k75fexGpIqo7enoDhiak8JTDukD381yyUN3K8VT+EbLmd18pKP8pokWm
F3cYTSoODrBJP55bwyvR54yERlCUEAdwa8VN2IdFY7/TBz14xUEDUjJaJTkzKnIsWXY35Ywjdo4p
Buq7FFa6CgQpWJ9848Qzpu9lRmvUB6wRysLHZQFrpStLJYMTCcGhh9kGduDjbzngocdiLu5rtvCi
MLbxd63g7PJvXhUfCddo6y1gk0L1aZl7UoZnlz9FQYDxqkTsX+5CIB2oYWEubROUUjNun8lkcgwm
J2HEuaTpmeQcRAsEP7RaPpzGhCXniY+VUCw01KRe02TjhC0pBVJC6kcPi0W8MygxQDoWw5UvVNLZ
WdZNtrFuB4CekovRr+2vD0g4Nv6wesXgiK38XdBEY6FH6F4uShgWqiQUcw3yiCBpoJ8594sxOU7C
FNQ6DBgob6dGm+aqrEKo7z5QFa3EVUkCH1VvYueyVZ0HZ5famgP01c0U4BpctgyzjFsWWVmJ/RL3
smltotFxjqAfqiS0nnC7mRzFJVHke+1Ahv5UrXNlW7/8TLxYkgwVkit1iUWLOCNnEolyPMcHdPfJ
gBsv2xDUU9p10rXjmmsj0TqHQ+xlk5lrwIyczmeKDg8JJNE1u5OmDROzevvODybf0lnItNBjyv0C
3NpR0+WSQQM8Tpw5lb0iRBSUs92Zoe2j7EURW1CMRt7LMlUVY7hq3o8Bg729PwGGPgqdACohfX2P
XxUOQBB/j7kNg0NNnBnOGHXLhWoRq9Q9X7vj5jZ0IT4fsBK3rkkC1IdBIhZTAwnR4jodxzQVqjUk
v4yJ+HsnmyMKLV01Ane5k/+XtRgPhMQjrd5ojYaknJlIHcsr2yTRpJQPb4ZmjALGeVQvBluaidWQ
c9W0j9xUjacawlGmMgPE87eSgTtc1cZ3LqfvIpStC9qTgffUDX+lk8uU/B2FIDA8hZT/0C3Jgicn
ZdjaZlbwSgKSuX656a9YcMBnWJAcd1Aso/qtf5hCxq9czmS5rx/8S9KDBwzd2w2Wsvi6lrw1P8Ll
Xz4V7jGVqG9Iqbt9LLtKyOOeRHguwoKjECFB761CL4Flvos7HMcU4wqb69dZq1Djm52XpmT0RAss
OKSlLO73HIrANv2W7nv5W5SHLzWsukXuHEEU5OO0BC4EOgAWkWIYF9LszaqwXr6TEjclHsX0nXaN
kpJKJ7tqxWOCAQZFyrUdryQtDCEU1u6PH2iDjKYGdYVf2l7y7YPXGSyR9cD1X9PKloOuPUVbkf1G
UuhDPvAgBULJW9M4lD7Om9mat9tKhFc03MBNBk4QWE8z0ZvmgddIll+eJ2HSSSkokVE0V2KrOYQD
CfN8fYdExzmrAYtmCiG/3GXyYu+lxPONpVzvEzsRxKdqvGpnWRzAEW20LUrW9fWelrRaVKQfddFk
hHawpZaPb65nvTrwqqY+7vk4X3vp4B5I3XG+QQ8rAtaqKJ5SH9DBZpzllIkNoEOdv02tStz1gqwu
2eqhnKtI05PtPX3b8SzTvIB2haU+7NE4pNBfACiyAMmBjleqvHN9o3MHrZGCuOfMceBsdYvZMrAO
BD9IQkGyEtHfy+lHC/lRQQBv7+Js1K/B03CzWOuobFMBBnOtXy2GIpVMDFW1bxs+V8amqdP9Uqlp
zPqgA43ZGwlyBkZQ2ah0Ooxt17F0SvQeqwu1a/MuAe+P62RCEoijMBYAsxnhRIwjtxu2kGY4fOcm
q0fooX/wnkDJ2Ga/apjBR093f2u5En/vn01VdLHOwkLMiq9dhFkktHMkZlErdHpS0ML9UmPOqAUi
WJ1LU8QAaloDA94yX3jmInFRFlWNGWEugNVFPgzVf/OcK+TGK4l+jZTve7u3i07j1biEmvKwIR2Z
nL00a39XoK2wyhI8OgKH9cKBmNgZE3/v4f5WSF71yDuA0+on0rTMqvkXdK3V6czQ57uOQh21vicq
30936ho+rJZi3pr1nhkNsBWpCNmYupR40yQqYczo3Dl/RHrBrLuD0vNQGEW0Ap3NUF6ZyjOg4jAu
HfMZuzFxq3/rW/yWbOd9iVmufZzEsZJYprATLSJaWeulOeztylVgAUo1x8Izc74y/Y9xGQBEV7/+
eZ9MC/vwzlzn4PgjMXY1Yk/mjtI2UQCdwFZqlvaP9qIMBEVcAYU+iMoZh41LOKJgBbIBaCbBIPei
vOKteH7D6dhiJrDfBYYqLjwhFtMqEv407ktNOpgcwDsVQWjlj1LpW8GcNtD/SMXRYqsSdAeaddbE
s3AobW7Ggt+lWDrrHU7TnVNNUiWPWYGbGkzdbOmGmVfjJ8onbni54KEFsx+61eRS6HcSFvl3bRPH
kUcCn0l8YDC8KvlrgSUheFp/ChSGnTkafNwxvwfnk21jOpGyFvviaKzc+MV7hBvILNN/mOnhAr+T
PtzfD+BeCZvomVLww668EfiX0cPYVEuHbNAiHgOrB2iMtEUzyAKxXXABm3gxBk6qklXSG44Dsfyj
95u4eTndLEwSGdxthMCiFYgdOLr/pBUoNT5E3U4LAQCCycm5zXPSHIuZtZgfX0OncKJ5HCb3BEto
B0PFnwGiBzEu0cW+zzyV+1vn0tkVP++6ViHQUfm9DPfSTQcvdoW7csXYCtCvMrIZVt5qW2VlWYg8
qxsEJxz4S+WZZtK6jbhja7ETbDX6va1S34ZdJSRlzMjb0HQwiW1Pvk1kuO/3sXS4yt3Y1zmeUDKY
cnlEOF0OAioOqe+J9g4++vPzYfnmBnlyCDQAmWSgUpMtSi7eqs/VM4TAus4QxNaOilRZBhIMhte/
W47uxok5uK5dPMDTxP0oDvwP7d0d4kXfAa2A4wM5onSEqIrLmAUlIx/3XFrpTVCgGwwH3igXxgeF
8yPeuE2FFZz8d2LJv6ExtkoxiH/OJ0tdGXQc8QDtJQuqpKACwByM7EcE8vXl4XcJGIJDog8vVhrj
kOywwge08j2X3UEFA1dvmsbDxXaCdDfBsfVSnvYrDtCcJG3VutDykZgoGdDKRZtB9yAVOyPIO47F
wI7CmFuzdN9d6kICGPmtxQE6p3cp26JA8zkEsnZ5W54F8ilCXi7pTP52ZAqpL8lW6UCmFaU3w6Zz
6oNvXmsOAH7DOtvJeMirEhnwq3t1l5zOdLA8Do9Mc6uplD21BhFj7CkEhJjbH0SaEDTCI85fEuuj
AkBsn/5AvH9TK7gsHTmVlJwTMTGHpkiTUG/9PHTeO/xaHFn01zh1DwANd7ZgjCyPzVwLdT76c2F/
POjUUOk4unzB/aWa30swgCXY9OI3NOY4irMBWfkVMwep3Hoyf3Y+22CIilxS6WSrb/52/j40QIIX
rrZNNjFXj84hqZxpEv64e6b7qshElB3x80hGVjMyd7On+4iJarhuOOAtcdPnWnGV2rTqmdmDjxzI
ENkXE0RGPui7+DqDQiwVAvkd8K8bp9OVBALBPSOPMXf87TDfbbdFUzs9vNbW0LE77oBc5LZHMou2
M77xvVfdKiZu2OTPkbVOpILLM+j+0MDUxZWft97oIChfStPaErpaPfmBR8kwX3sInEzE+xyNTRrF
nQ+u0RoOQeb6Nqq0ivodjYd6Enl1rh5UpHyiVZMvBIrZsQVmu09cuTFio8BgQwTvp8UWMAoZTJo8
m+sl/ZMD+ImWJzjEPubgBx1cBo+BZhpIqp/rJczbKA9jPgIqWflcbrf7qvbtVnWMkNnCakI75kYD
rPuQUCv48DqW1TbjM4dq+wDB5A9F7xVGlbGeOJWZkKoI+prX9Vz+ABcnGZDU9e9zB9f74cAYwn46
KlQnggA+1KV4T/r7j52aZtcPGIAc/1gRnkIb7fQ/h+eBMIcut2jQhkFa5IU/Qeis4kOD4dakV8jH
clfRBG7SQ3Sg69y1O+sErYpbG9Qb0m54r6nk1X3LZ/MV6hItvRujXrmVRGZgnqjKCP4kk5xJk1zf
urqDRcg321eXLZrBJ8IXsibSa73pKnTj7hMOB0fNqR7sTJzDKHr0Q4DCsFIxOwbc6TFiYsTcdC6p
FTH9Ncbo2JermyaA88Xe5Mz4aDbQ6+IyTLbLQSByPVgiZ2p+V/cgJk46TRcjFm458Vq3Ifhj6fvO
Y7yVXqAd9K81uTH3Qn+b7Rrk5PLrZdqSdjm+XqoZv/V5L0OScE14J3LkVgLxrTnXivNoyxtJaSRY
9AKiueeIbbyw/EpNx8c52RZSKXhS5+4FsMomd35UjTCKbN0fH/qXNkyh5At26c9Piy8Xle6ELAtt
MaH1/RXIe3CqulE7MoOjBJxUOqJs5gMXHzKs+tnMGJ/0GzJzDwqp1fuCK1KbFZfyv1QiuQ1L5nla
9Ny7g2VxJOzu4mnQFiMJFOJEY+NrcjJW0Hp+4HOdr7iKKdyjqSmV/waE+xYqkHmtpd9si05oxPGn
u48DGz5JQFRZ5MVhjKeiRWRKs1wJPmkSqeNo8iHdSkflkgJ5dc9TZtBTQfMLgFQzGx+su3gXOh8S
PaAehogKozH2o1y508nCMh32PQnPtdRnYBpBvyV9bwzzfINZwnKt7TmfFlVl5YXreftSjazEdJ6N
b9B+0S5dS6Rd7IcIMlsLjiCWXC/44rV7AgvfT0BLLLsQ/Gx4LNjiU8ddW3P0rgDLji4OQWe6Uvr9
h1WjxoJMsQQqb4jwjWsXHKT3JrVoBTM6OgUSyPdBZ92gucemq8vsqfUMQXl/PF5b0F5S98GNoNZ4
oBHC+V4ARYvxxAU6auGgr0DqIQx4sbEn1wR8YaZT8S/T0612K5kamR12kzO1PEKXwPUzTMPpECqW
H9FXj7uFo1XRMnfd633Xj9WzYOiLZBOrPFQKxGTUWV+zpPACRUOP6TfFYkDnbX7eFxK82bYmF6qO
gskYygfFzcH7yCpy08tg25A1N4Ajh0VNKm6Ux3ywFWYuIZAfSiZOTew83b5XgHJ9dJTFMtzf1GyE
Se+jradlP7KM4hw/Vd/4X2vSoeCOzNKFSlPQ2uLipOu6myryahTJ5XtcXtYSr2JoguZ0lO2ebcAS
7rrDheNHvlwn4joC7qQLDewT4qdKn1noPIwNtfeMiEE/QsuqGabk9w2Obr4jOTmETb+dyoxbZq8W
GrpxZkVoUwWjTnEVCXh4Yp4CaQtYv5ed5w6irNA1evKpqYm3I7JRGOLFqnNPpqTaGSMMcxzyo0YV
RtZG8cNatX3dAqeewqn7v55FWGaJw4oL9TJPZyZV4jYlHpxR6UEIdYrerZ4SnKUN/84POrAsKE+n
m+uL/c2ZgA2H4ubhxhn5vTchqkdg3550tODJ8XcZ3Q0JzuovqIvtjq7MltW/nF+rXh9zqGKF/+vg
jxfM43Tj4mLhSuceYML0MbbknoP4uaG+bx4jTTpolgZtU6W1m+GiElZJT9qkJyHQClp546/YgOEo
gArEEbhK4rFiQwrqQ+KYOLCHxaGUrFZsZzqjNgwxBYckLX9qoP1Z7N7WN587w9lfhZFTHC3oY2xF
6uxKFFOpjgA5YZNyftF+r6PtXVw283KrRAL14FVxDghElWMx/ju50JCg03VrDJSBmTjbP7pMk0YA
c63lbPaaZDWQMQT/X92tmojkH/dyW6ZjmNG4+zEq8Qzv5ppb2ns5UuPp2bzViNGnmQli0fnWBUDS
g5NN+xui7FzeP8NaDic3lOw2FDmgfHHXtnBZLpKZysQzXrsIkeOXtdLKZ+r2bst2WBpPhzINXZAE
TzM/wVTAFQ9Z4m9QZ6/ElqjKcmX4u2emSuwFS3L0NCzp/HTcn+euiXXr3CWmmTWMeT9S6Jp48LNZ
1E3F1qUChOXd5oJO71ENZ6RpghhhmALECXyO98uFi7qSHxI2aDM/nizpgsR0mwayLipAxudlz0K7
7oqz8Vu0rhx7/Ht5vcklvzkWInGKug+xvuQD8ArdQ+z8hRn1UuDUoaGVDT7TMI8j6JUlml95ZyvI
Ad2ROlhqFoRnbXHhfvAlm/1uTxfvCVx0Lmrk1KrzmweuSLygk8zG8IqOd/qrAmqFDu6HOH0yssfc
HMC34TzTnIzHn2FdBT51FkyicnfSGfZGZJBZCQVVZw53mnYtlOwM0I41OnL2tx1eVHdMvb0XdMva
djgKrMiSrLZJR7Pb/iKe/pNn918w4nUsFxISygHAOUW/Eh4MWyuaTgxBPel++VlqTHPgb/D9KBjM
FtRFzJ5Lhhz+Xdywut0l434e7MvF/uxGFaBX+VaqSpXems9eQaVUo8SPhl3m9Wy06ArU+Fb9jfiu
wQU7PVI37J3GVgPFRVaVvdfUzRmN/nBJz/6VPEnxQfIrs60+ho15BvSSKW8B2WBTDr2QKkQyS4E8
BYH81cbaprwa/+hVRyKOq3/F0+TV0hD+s7oK18r5xVfj4u7gRG5iGCfYlnUZTZ7YajRRxOeiboS/
vAGXQB4dlrmNur9GOAo8t+L3BzjgEOYVaLeIn5/0fdiaXblI7gWDLexFvO+mUy8PbKEJnFK8mlP8
7FWFA2KpQoXu4PVk6u21ovVKQUiPTmYLYprIxGtbTWsEul2L46WYrhucG8UBihgGW661UhUgqZPu
/FEAKdmQRuLrz82mrGCzPPbBeQBmRI6nwscY4SEmXs/pLvDPAcc+189RPSw9STEQEFBK6pfkBmh+
HyFpX8VQzNzwW3Dn/SntgPLSEcEWY3elBxaVX6Bn3zsxgorHLu4aEzU2+Ay6hA5cKoeQtiIYuwof
avYBN/nqeY3r858uZYlt9OZYHCxaSZw47NATRxvZzqwk9zmpQy+FKScQtUR9lbGmFRT81fJXq6Cm
no2UtI1CMmqZu9jqtyn1ErVm+TM+XpO7v1ZlEmGaeV84JBDXPyCnq2a9bZ0ocVMX057co0OUERPJ
+Q7IU/wJk4ZSb/cerOOx1CkRSEDxzw+HAM0kX2LjBmi9d9B3GhUK+shb07XXtQfdgSvykK3kuDZ/
5KYjyJxthL3N22m0faoUXDSAL+TX/2Rv/kuujqg7Nr0+QEu3Udf6tDNibrxPgPTlsi6iku6desKM
iVmcFXDRerMekwplA2rVobztWblj77MwfxIYRcJ9DAPWSacVAKj8sPUeH+mv8HKJBT9AQQRfBIbs
7jXer1TssLh7pAa8F8h/uLSp0g7prFwMwW8oO1NePqWcLNRaPEYa8vCQdPVz+xHWfHdhrX5yayWb
815Vy78pifwTM8S4Z4yzeZ+rjypupqf4YflV+Y3B4AVOOynsV/3yMmS7OdEVaodqPTWRjoNa31KE
uFOF5Tit8BiQlSjwDUXVsMq6Fow7bQo0s4C5fcC5rJOx63dFmA1hjyaDHEspvR77b39smiFQQpyu
sTn0r1qHDbDh2yyVL8fsuqyJveeU4uw8E+DGPJLCMgw2YBzt4fVAkzxzYo3g2pW4wY8Dn+dAPI8/
a1a593TNRx5mSk6UPjea1iX4nrQeX++OZqrDYWcRDzb4zSPXFc3EHbEWYRQXwQWRzWYidWjzsOR0
1rWNZl0WKIa1NId8Dg60WYPHCPKJ7pTWZjS2zur02sxs91xgfN0v0o8fHolu52g2QjGmRIfT2ieN
OX2tl1var6V9H44suL8A7Xd5JYp5PW+5iUttaLiPe+95a8gBCODybLDC0RNv2KCIwmM417sXl0Cj
uptNM96MXH7SjS5Zzuz2xdhkkwYMghc+R12w+hFP12tqsIJBcl6MzqRHX8aGRMoZtrwDiu/4ZlgN
JWJvDNHCni4JIiHl2XsVf23edtjuEm/5NUBufPyuVb5SfDZ4/y1y5cpoIsL0PSVWhukBBb6Ap6c2
nWW2uqpoIRA5yN0JxRIc8tzz3hLQz5HhdgPZzJs/EJd6hhH8n5/RA6MFulA0g7qn7UpbxQGlGK5S
SyoDjVs/8qS1+0UXUf3u4jDWqUy0CusDFbB/sCx1e2ZXY/BcWIn3msBZzB2v6vlSVP5m6VZAbf2L
b82cExc3XGdzJ7o0XNZruIScFAiLmNgC7PrtzF0CHkN5eK3NFg8Ck6QhfbKijlipce9tBo8HNLgW
N4Ph7txTeKaWmoZGOnBpD1fF1623tfIvjk1BB8cBNXkAYLPhdqjjEizoqpyltaM8qaJxJYAow35W
VSxLLsq77en3DHkgeNqJHqKWgVkyQ5Vwt6pt2uxgdqROICioGVkbTM4H8+wLuWEwHWDhYC0GESXE
wd4yG1nU4hpJ2PpxG6+OuhEHcULwK8GZ+wLhlaMeVyy9OQw87GbOCLbGDx6rp/NWt5KZXW9+0bLB
H8gUwi5s7g+m/nmteDXH4pn+nP1bhlvtGzwkhVYz0vFhRwyifSvCmg2cA5bsT4WBd3O2jl82LXmf
yl6fGOslSoQ3Z0IqjbyYIupcx+rXp0HUMwOILcerihw3Fn6t2MUjqK1BDrxiLzB/X9ayFw3nvqhf
xDRYXWZy+KX0tk5h3Cltz5wa69VvrYkX86s8QUMRJ8P2WlJLz69MDMa2RO9cSnyqqX6FjYtdSfmu
lRyl3cRJ7yGjwCQw9j0CvEVHcZAyAOufycapUFNtQi7ICiWZmEb8vXoqgKt+yr+Tn5rDXnbSp17s
6/siUFJUsc9VJyy6QmJKRek/WhEp+265DIpIzXRseeDYXZ40hLYku5S82bQRAXksaoz8JzmkuwC1
kuzENxLFCF9t0XrafIcFZHw95oZqAX/8bHSSxDF3L6uti7YWg2eWUhusMTU0Kl3Sd/Ymj4WhM03I
m6A29yAZUHuqEtwCI7QkCl8F5Qk+Vn7jM6uErD9W7eRXdKLFenIEWbbfa+ya5jntFCOgzvSPUES3
OQrly28+O/nLvInoX4VVwVFqLvOK4TbETOXgYX4mDDf+EB2xJv7B4mSD9lyX2FOYA0rMK+FZvSmt
O9QuHIAq4xTFGVMV84NahqB0S0w4s3oIh7SsQW//lkPPunQWWey6h0cnSn+K0cI4otDqElPgJVWx
hm8IOKlsfFuyRHGi+p7b0VighRr0eDBvNwc/QIxmbtwTooq+j8qxHfhR53MMJadFK6UKZWQP0bkp
XTH4KDMxhVVs7GZ2blfdkcJKy6szkZiwmPT5/Gt/Gt+//YX2XjGnTvjHY90e1OUewlaPW1MfecGr
W6EfY2y7s9sSZGB8su3efUL5/evPjBwUHjgGqhXDdTHKYK3j6R4I4rvdMDz1BGnJGRi19pZ3sMRc
k5o/6tcFEuzmJNzvmgO4ZqlgZmqyQZ5f/uHNY7FSpA8G3WhSQ/pk5j/vVs7JHvpXwh0FbFYCtq80
my0XKyBpwPneOb4HyfSLmzibp3OncHeZxWATk47iSFmy/UEt9jp6g3ZqcaoPRyy9H2f2dwMXnAvi
6cMHPXq9upc/EI88/+NlQhJhDOoUzEsG/MB0a0Piihj+g/X/fHkqIwjdZBOaOZvtKQGd/fKAB8ch
wS9B7UxMJYGDKuoPxFkO883fycyREZsFjHf98YyGcc/rrr9aYckfU8w3ptvfIg+Xmm4vHvXx/Kaq
Mg55L4K4cOS5na5007mFzj4yYau/Y+3GII1AvrBkDk8QqBJpCquL2GlFkJGMnjguklqw5WLWO/1n
zCmdYIAJELfKXu9AUnDnGfzwAQm1uRpP5dDuEYXb7C7j6BobkLWIGltfH0INK+NZqEdMLfEdzslP
fBD5s6bRM0QKtSLGqnv28LT6KT533qQ8PL8GUZgkDL1oWLJh1T5dgWqu7Er/sl8J70payYr5B8bO
642QbLzb3Z82dIFHlQk8vKTFRuxJhODEK7jyl+ftcBvZoMMkUsG7a1MsDVJgBy+gMDkrkBlh0XKA
GnWzsOSXoQYXLDgAM6hBXTj7xtxaqEi8erJW4C5c7XHHoKeC+QkinLAlJ3XlzfCN+SuaCLrHa/6L
vVB9yb5kxHZzEsG5CtacrfFUbiz+RMKvu0EVIDcjg+oYoqph5b4t2WtP0Cax9d/0Q/VRFv/+ZXFf
RvTrKMJ2uQp9cGj8wECec+IG1ejIYowpxYHOcJ90AgwQ/iv6LuVIXpJH1H0Ie4y+qXK0z9EaAsgS
TX8anWW6A6c2+tcAxoazDXMmeWzDta6mxaSZral63Qbqc37v9znPyi3iV/vTYBtmUcy6cNq7tfhN
bd4Qa3ys1QqGHTe1XXoB2X7aL3m2vj9Y9BK1xicZF6PB/oCOKLOLbv0xiy7BfzMmk2K5kTvJ1xJR
l228cdfo1T+5/BtNbBMxWiR1HzKMN1wxWm8+yFhltb/xPpRN07GtxqvM6MBNnyrgrMJ4eRdR5xr9
DXCAozrjQmDr3vtdMVhtmSqZGGhuHzFWpeqBXQrK/ev63w78Fc+Rm3lWneymOCZgdPiOxBuIaLIP
AeCQG+TiYWUQxEy+/iRCk9giFdIOECD7ptOaERakVTdsgcn3NXkE2Fzwb78TGQcwQX5WDuzfxHRi
q6Lu9f/Yk5wkCSwMPQfbKw5fzQQ3uKMhOKoA9iPE0SHDVGMkwSwoluEA1hKvSem7TeNIL+Mi39MN
ixnFQIBEz0KyWOC9MMDG/yHCjrv/6Q6f2KCw2WYLPsN6BNqkE1XA7WAOaWDNDwl2yr3dx5Fz0kXV
3cDgX9C8307iita7N65kKD203XKxhg7pQ+7z77eD1iYSRv6cGKvfF5g7XpwolZWlRHZX5NkxySvy
6ccxS5wwAnM6jUHnumiilH/NmMAtSADdkciWFP4NZWIHxNwMH6F9AWLu8SYVFqKMJApAZlJsTZKT
qwGksTu5M7eUt7528TkOCD7w2uTiHkVbyqePXZ1PCHifJIeDEhc/o9gCjS5hQCE6DdtBtUQ1rWC6
qPZG3kJtMdBwo6HYUHeP6EwHPm9msnlNmHuV2nU9mbOmXk+RWaClQxdWyUni0ooELPunuOdhapPM
3iNHlSGkmNNSXibTTKst8lYUHk4Pzkf54KGjYrPSxTTbnmH3Gmm5MNIhpS+jSVjHSmIkHPLKhubY
C1TaD7zPz4wUfMv4GpD7W4OhX40RLrYF77aMXakZvgtoejnOt6bEtpuTttWXW5/WY6OWOxPXARoS
+vbM7NSeKVL9RBMRbpqMqE+HU3tl/8sZ27K4fXaP7Rkf9Nycv3Or1vhMtL03ouEGYCxFQtwCR0d/
5HPGb0QVXSJKNzuBt/UEl8U5DXl9p/E/dmPEWlBR/YDSVWM54mPqYLIbLQeRKhnPwLCiWOJOOWW4
3nh0e6Xz+nQkVODJ7v8IsHAGGlDu5FAIZPYSWsonbV8SAAq5uH1yDuGpskA8SdMJhu8f6+GXmZ8E
tcWLhYYnLuAVtGUHKWEwq4SwzmhXgn6qrOVUCPC69OUsw7pF12nKE7KW0CBcnTNKaRq8ls75b7Gc
M3QPS/sRIe0NYVmm2D9Wv54qRZ1IIYytsZfJIXoT15uI4XXhSEgf3LWc6Zuh65XNc1PDb8Xtah2R
C3by5FtK0eyerzqXMJPWuAFVq8FIfg/Xsw8nO2HJu+FmF62T8yNaxaRJujFOrTYdvsLOpe7M/SXs
5Qc/dkvc8uGsddbE2xP43adOkWjn3H2QZC08Xa8ZrbzRDrI4laL9RePtwf4SjKbdjUQKP9rR5NHw
4LGhgarSWUoTX81gmanjfeUtPUlxH8HO1FkVgn3w4a2Dweo2B/qn7iPAvfP1lHQgaklOSuNrLdNg
dhDlnkdRvF36EkPf4d8d79fHqO3YCQ2d+4N+UyBjE7+kReFxtVlfRgxYSayiwoYiVzW3RZmcSwCg
wcIZE7+LMqkUvY4MDjHaq/T7WRUxmRcCX/8xSn/6n09xkVNODUprNRsB/2x4wiGxd1e/0LWsYwKk
w3DrVVtferWQkZaJNwlTRfbr9SPA4CUxw/xBaLNofBbk0/rtNmIQB3m7pBI69O6S0HZgqZwJuNQB
IbHbX3OmrKK5E2SW2OCAwRb28ZEW13reJZHxRNvamhwPAqbWMAYFy78k7VsqfwzVsZlMXsblEbgr
Dx5mF6pfMgaCbnht+gZigpDReMFkduI+/1RzvfUsjBHq58cpWJ+cWiFt6t2SsSERvpJJkUZiUlny
UxgjEC95fKpD/qKEiMk0GyQ2a0UNX6t/+FtFTklvcB6WZEWaXn0AVl3Ki/PH1t5wdePe4ngpf/ct
r9MIf0kSJ5qB4ZsPbahorOmlKPfBA7hpT2UmzTpieWrjUMphdsSMQGeazSVVvunlou/KZA+n3wwp
ATQrZvMtnj89VUNupxbpijqKDqKuZkVBRGwD+p+7cDafL6y+mMLxRGst/s63wFyt2ODfOPStPchO
tFvgwVNymhvBf4BuqIiiM81yM5m5+Js/16wKL5qvB2y2DGE+WLK9B9je7K2SRVutKMQVJEJGHe2D
Do9rg63hy/H/eEeKLOZmytpIsFEU556r+ENqGV7+QgIYHmatZGFhaTJMf2gHDu4p+mxsHg5POTEH
qR5WBSzStHaMRducTG/j8+lPw9ZH4hsZwplahUWDlSgngFBSHkHkbojNZC6iQX+81Ww6T+zBP/1M
/56bo4CumQ1yITIYhyM4pC9QCck26N6jgWvqMxlTnXUvnh9IKcEZaSFu126aQnaNZMwGWbhEegXZ
qaCzCZeAK8yYFREfsTyWVYW1LY6+bgdYvWFgPUkipyei2TpP8y0dXyOG5cKbWx/l0MDhv0GNc1vb
oGve0P0ODAsTMviY4JAAZxvlFeXKu+4JKEb4gALnt6A+td3P/V5UjegZy7xZCesktnibsbDPezqX
jWtrouzbzGzSD7gC1QgDnRte36/1FU9u43rdFMmOr6YPVhIvM0LETULqwXEUYJr4A1Z736FBt1KH
S/o8IwXYtsukHeUwSFSJYSTMk1OfuK2ZpiQHDMN++Rt9rKtWH63rNKihIE5KtNxqLWsP9BsYbeop
1IOuVcR/+p6KF2XmKUYLz99sPStRAhXC+5M4WQ/vEfZBoFzI7Y4lLkqNZYm6kjaeWjoozqPQ2fn7
vVdgXe7WpOaunn1+xAcSjsD4gYq9E+0HkJfMqoCXULwPtEL/00NDdK0EUedSrMhkTShj/C87m5e0
Me0bB3hUys/oqtZvhD14n5b9TCVaZlPJFzEGgHvWJMHHd1L6Ki5HY3oxVplQJomuGPnSSTxw2boW
fMRGUvoe3paCx4m8ZUldetEFPnmB1WpzwnIW7rqdoBcPrsb2KJnnUcR9oDf9w7v5xewgFMCXge9x
eIpjA0DlvlfYvkcdFMIfxvm0bzca/fk0TLaOJuIasuHWQ4GdDjMiCZXaQ72nby9i4QXjRl02Yy5E
odZZc2IvToOuoh328zf1VD97MkPgHj9JnUQRzHS/DiFT1T71RfuFW/dj8WIZX7wcQxXdBnZ00bC7
2vStvQXplZl0/k6Fsdylou/KWC1O69JTGYsl2x0CyTiDpztCZhT27LHesTZmmZWcf8gSkBB1Pech
433thieXKNbMtzpH46egvMJThKt+iHGTv5B2F5x3RHvFDKWbbnzyi8CUQWLxs0foaLZzMkZ+u5sf
PEDsp+Coetv3wpl2FXLj30FfvWwWX4AjssI0tqRi9r7I20CQA3dUQCYNHIm1d1WGjxy7i3R96Shf
ODbzTur/KwiltTUUpRF8ITd5A5psoq7sgio15WkSTtsS+VODTJ1pNPDO4G7TBDFiD/HzbSbHDgc4
S3Y3kzRUREG7gT/jE0KKW0nrwp1geqUQVpoOd5X/jyflEp536b2BAH6quijiQhBlpI6OjxnBD5+8
RmafHj5iImBHxYsCQnEluNV6cjhViBPjNtRfGxS2XTXT6zuJT0pY+v+59RqUqAQJCt7lz7ZYJMMT
relaby+NAZmA7iJC4gAlfgEhgAOQNsbQsDmXW08B/vGSQV2cdkJlZuwEJViJSuckpiZXtUnJn3cA
oBcd1pBn8UlPCk/GGp5oqVDmi+wFAP2jCsFVtKXFvRQtIWRH4KXWxL6LwUsJSDBAmlEbUCT7oAY7
GmS/XoWXh2gOEttgk+WD11tttMwY8kj6WFXzSOlP7q4bP4ogkwX9gkgDf7UVsLaYUGn+S0wWPT+E
zvhgJI6RInu5T1H+Tw23KS3grtMIHyUQiO2MCxbe60f//HMX+9zURRoCN+0hNzvNnTMzj8bamTy9
eGy1ew0zlctRDhk3aDy5S+fBbkpxVC/ShdVl4Jpugo26wOBfAseHL+ix/9sUGLzn6xZxPOjZ9EKq
FUDRTSmC7nzovWZItaY9U7KtZHLjNLYnfcBKDn8IEqlVxzvJ33BYzlu8+minrvZ/tFLMvP10hYCH
rDfYF3EFtBhCalXT1k3WxHcbaZR+RAtz4mrP1PX+jiQa2Z2BjKQfvu408bDU429lr7/CMLg+d614
NRpwV2l3CkA7w9Scnrxis7AQfV8mVAt7sRq2cwnmRV9d1t3/D5rzw+M1LnungocM+v7rWblciQUe
54AO4FVnIlCOTwqePWIUX9B33wz/PT5LGtfxFsCGYt779SxPHE7JTV109hWYpsJhtI6kQB1NMtXl
zF2lx3qOJMUNEEXw6/PARjDZlWNjyCe9TjD11a+WkrAci//RoTJjwv2bn2YXlmBbgefCuGrKjhgV
f4UM70/dGZkuQ0IVY5I8Tz+XVdtb4T5k8VvtiKVMHDhOImofmkTGz+tSMcwKoL2CM3LI5WgQT59+
kV3oAjl/6LQV34bxYjVvsqXoh7CaRLSkg/bImxFliIZ0Ud1CZVT7PvtGBxE2HTxqy5cEa3hyMkLi
CgezHdj5LYjKmp5jClP76fHkDhrkiIvAkvncnzicyK7Pgl8Odc5+YWjx1NRkooaJMzUbLyTntz9Y
1k3+NW8upsRtENae7XMafHYtt8OvKUdDuQ8mejuuyfg8cPSAqH3kXkL5IOtOx+V3YpM6VRea+A9m
UXeqXeYCFOw/IWx8WhippydCoe7w7EILR6Jd1fmmVyddSNAphVwolsW0Z0LT3c6z7t3deSahmDOq
CWCgvSKONAqH9hPDxLgZVeWWWyYjARSgXQxiIxPXh/FR66QePhy7VopxdqjJqRWVv2IHyGl7Rl/U
ZHbaZE/ng9hvcciymuRQNhv7p0l5qQ2AzyRs/BwCciv7BWskGHrTpuEg0/On8i68P8iwzd8Jr3+q
bs/i0xJ8tZA0vYsRtdBsxKKYccMwp/Cq+vYLK3l12m8QnNJa6LsxjpkqYM+oIaLMB/A3Gg4dzVXn
UgsrXJOUqDLG0NB/uREZTQ2ri00F/q0cjomT2fSDK+9AmtZG1kfcjFfY72yVvij98RgNUNS8uyt4
ydcTp5bzOtumJ4fVV11scx5U8nZQVGTFi6b6Z5bk8fXzRYNCHUJkrO2MNhl0HXU9QrXLtgnLYF+T
+kyE/TBonSlorJ+Tj5zSPP6sOG3W1LGhY3OczRcHyqrZJe2qmD/Y3WZRAhYhp/XEiQxQq9s/o2fA
0NmxbuPRhCU++gQWRm+MqoMXPjiyGqHMIFYLMk+1sQEQASysXcKn52/8gRN3KTFBQDjU1b7FvtCY
90M71wuVuDe/KbTx807Dpb3MUglPMeKMuQOtatkwGv0RoTBOegy/+1xwMbOiflQKPDrOUrx0xX+3
s5rQL7/9fZAQSOjjffvzP9l6wxtiwRjyNIseKtIyLWW9Bx+m3pBWJ79OfFer3RxkI0mNRTM3j+Pb
jm02W5VBV6Lj2fYf4ydybkov/P+V+qqso+UzOI48fzBGBucV5jF3wJ7A9MoLCy0UYAOaFKkRC05H
eP6NxFdWrrCz3FFBi23Jm2Jr7lrGOoHrCXBOtLw5UbgLm44cBRXTAGuvo8VQoi19PmN6U0fOqR3K
/PZGhZJy6ZkdmxWi5tmtUVUmJVlVSSdqcE9P3vRHMqQcMerqNL4T2Gj8iLwZ2iSrcusYTQon6ynF
gYtn1vatmeJ4xJmtysJ23BeYFnKBZZUKvaoGuXCgKR0hbrXANmBZxnZxJ3mRX7ZUvM9mJyuK9rRY
J2JmnmzUOe+OpTNIbQpQfMgutI4zZrrwAL3UKv+cZPAdky7y4dVVJbWRxrLPPZKjrKhdT9dHwFJg
0i1qtUcjhlvvTb7lwyFp2jYIodYpN947zrBlWYO8KbiW7F3/GQW2aT3Con5ZkF0+ageUDriHxZzY
eEtCd+uj6I7T8irrEs48+KB/6cSwIQ0WNL2PvrPOVGzqkh+1Km7xXKJchC3NoZ1ce9/V1+EFYjgZ
AQpT3Ob+gkeGFRoS2jgNoXAH+LizW/h7gOxnU+18WJiIx+N/zcetEoDb3MUaFnYi60UGAsO9Yv7b
vzOse4raIJIiBO7St2ouRfSBy8Ldv9ydu5Tj9blwqCs9tjZkLrqH58EXpTc/Kb4dUuQAfdHB0tfJ
LXS1Is1delquEkvPFs6X0ooQtZ8TvUYc1VdghnGpQF2QEywQmIaw4rSgN2XDVWPtM8ANuLUfme5Y
GjwhqSUQJIh9aiHyB83oN79PrunpAC/qqQ/I8uDZUuXQsWaQGrsG4DmLtcVkAdvQ5ud1cQs0o6x+
PJVthPyH8+zs1VNjNUT6c59RcG6gnsSU12O1BqglnbynwCmeNZ/U9OzActVkeM6tT0FroPmg3V9F
BQGNGDdXgXU05eVUAJokxyVuoUxOdawyQgEviCXnaA5PLDaw9BLt83Vo3S0L/L2BS24moLwup6z1
PIaip1T227QcQSyc55tpD1TSpSj/SR6nmEu80S2JD/jORRCBpS85VdaVk3hepxny8wAFrT5W59Y7
xEdfuDJCsbbWJ/ycrNbLeswWO5JnNY+hgsVu0VtBvng6TU2AuAbCYk6z+9R2y+nvWu0EdtPNjkEN
Pr6gWH0gkxwxLcYvDZUXPT0FSALCRq1l9pmtkuWbQ/8GY3SbNEtXwIj19ojpQSA7Lo+7pGmaOVMd
7RxYBZ9anFXKdSXm5rvUVhooPyFFCAIsCz9ZSJ2KmwWkSeaO/S/GkT4rFxe3HdlJpolO2rhiGKf9
Ds0WAzVUUqSk+D+yGBykPk5Wn4tVL84qVnWpckP3RLY+ZstEw5i3Ku39g4XVu/bS33t01wzu64Oq
WIwtOHxTVIG6+Oek1pta7AH5BzWI8d5R0TVjlyM0v1URDfl0d980oo5SkPUmIAvOq98UxPbfItb4
TVGSmmvV+ia/RSlVdAjJItBNFh6HXM6k06tiUFdxemxeqKOb5ic8/hORaUXWoINiQfA2u1x7wfNm
uSCChZMHd7d3fWg32P81s7zkvH34RUUEC3odT5vqps9T/FE8IqKtHdJK5B9yO2a+BM3DilQ7ctMG
RS6CLx6/0L50tNKkbsl/dxFQj4K4Nw970vffU0SVr983+nClHliY6DzUvWIfn4nDci0faHiYe20J
xYwG2j9/l3lm84KmJ525jk/beAnjGrhUQdeNsjHqGvo53ANdK9mLAzzAs5zSrDlx9vKnAQ00LcDq
u1kbRDYLFKnU+Pzwbk36l5ieTFh+h9qitt0vV8T5M3801sUoxjWMc9F5aTvi6YyRRSMv7DlQbl06
aO9uNvqDsDPJ4sSSYYn+0wViagq7RoqPMeKYU+++SiIUjMPsJtAQXlVLnZguGB8Bj/6Wgvj/dF3V
ICy2emvq9mxh5C14dIMY7+hSZPo29hr3pMPjAzf4QCqlfWOanwjFlaHm6t1t8tIseM2zNxjAV7nG
YYELKzsbak+kPzLoKvSTGJoUMaJ1UrVI0TTmaPGse7j6QU5C048WkULBl/0PtuMEFXu2wp2iMtei
Leq1m477jYOa9SG92tg1LNKfBf7QBOIc31Ax5YxB8KSPpY1islFcKo9XR6z7tfaqTcnWI82X8a2B
EF7QDAswWelheVBvYEOqsrLVVbsEEbGpxal9y8mct+a1Chdw+B0Li+SmIck5+pXKmRC7GQPY/EVc
yAAzAGcRiC79mUk9Iij6+KNj8lKDwi4pnJTGhGfgzyiQyxJBrVW/Xk7eVh3iH93CFdTDVI8wQh79
zxkYrlVpzK+VRTbaD6WTC40NbUxa0q4Ckt+qubfJ3OIrRaOAU7kasLx0nES2H+PKzuNjRKxzvWJT
2fKwjHDwAGw0K50b16Lcw+QoXnpK65vwhiahhMGlTiWnJLtSfyIFyIrYvVc7qXJVo0NTOqRDMqRr
M+gAq34EEitMw9i/eFiEizq1vDQTNEw0P+q+jyJCwGZgU48IB0tEhzGVjPCy4RysI2PWvSFrNVyR
KqyZCnHzv/siBE+CPwJVnRkgB6x+dLi55gNBeRFv7q8OAQXUaINsoXrc8RQJHCVKfwnjYbI8IUNu
XLFIddqbP3rg/79YjwSrhCk5qwhCDc5O8sjtFaBQhzfovmQcLas4+fFdEeQEdMXGyy0vT16vjpx6
M5ooXayu/lbpEu+5jf+KMfn6yKzjqAicVmCTEqtHGG64j+awnUpk8M/Zc7+VK065ny5t39Ons2k2
bPWLgYsoyR6Hg7DC8kcqmvS2lPMGd6n8R9MGpoio1V6FTmwtGCYPbcHH+q0p3fT2cVoBrWqHlYPi
4a8Aje4J8xVE5/ZWMmnFAh7RGvIUqUvXdPjb7F3rp7NwTwUFrEzzC9rNb9JDQKmddEfOTEUzwmMD
wLFGsPQp8KVNnmr7pg4tT3BFVlYSFCUDgUiFHX/r1kbT7Jw7s0lRUj6p8sOT0dYLbs65w8bSuv7c
nLtPNOg6ioVsGPc87qFELAdocl0j+Z2wGRYJPc5HBU4z6vTxaKHb//9SFL7fqtu7+kvbym/+ugQs
YwLLTlO4Qv9vERlYA6ZTU+LDnzNzWB5TxHkOWycHS/duxMlN0spUISad/MzvFuyRwFIWtzVtfwrP
HOusmynCvC9LGWXanXKWU/kqZb8Vuu2ppZ48GNVVCCNRDvNmDgTqYTHYfbggTGjN+AjG6zn3VHBv
MhQlG7bi7nX1UXxDsUo7pJ9wP5Yz89ntP+uUcyxO0IvL95ooN45Op99xwEzcSk1REiY8nQktgS7q
6S3YK1MHgknRdZ75z5DjfmozTIaAhXlHx8bzMiFeftFzXQk405lZ5aFwVxtvOKph47amhB4vOeiC
yrTC8w1wrAPrphbJAqa2DAk64gzI3LqvRFPYGyBmt6d4jtjxTd0V6SMNXPyoxiio0cofNldkLiJY
E0fi533HcX/4Ub1g4L8JoEPQd44GOgksZqUuH5RVl1S1ndbDlTC75DKllKcZsK3Z53qG/GJfHSlB
3sLYvZ7N86tEXQR+V7yiVVCJ0brlTwP/+HHWWcf5mL2p7usDMkdzzDOP662AGMn3xCxpSezTfQHF
n2qRsc0l7ri937Rf0lpaI7201L2qz5zywR+tW4mU1KgvBJhrUtLCkRApGiY1K2Ws1X6j0bzsxDMk
87W3LZ3l91F2OVmHZXSf2odBufHIcLv8vIENExFVVb559A6/LhTBdcLe6mduzsfzLoFwuXezlAti
Wpr27Zz5Ce/Z2ClMY7YI0nWFV/iM4li06OuKb92BSnsmsbKQzuQqAV5n4TJnUBqCCuG6nvSPRntP
9RXx7gt8iyWGwLXkAQ3IYG6bynpVdjGLCq327TJfwsAIFQ8mNI/Zn8oj+0N8op3AOOeSQHDvr8Im
ETs65LnoGAxYAJExM6C05sRJ0yO0uRAs3MQRqGYDHMwYgux1wWcUwTsud8ILe53Qx2N0CTo3UVnc
gIRSeoQ831+mfd0sao9BxrcMkYTtQ4115rdT7VcqpYMIRBQTyBIvaMA+opH6Tb4qW4jA+Fmtdaln
3t2GtoLGGVkAKBaPyKBbJ0ylv6rmhkavJeZ7rFV6JdTE43GJi+anRXtKiSCCtnQ+JLF5ZBp5bPln
zP7k/KsG/kfXhuaT79zymPEAuvghLAle1md6LGUiuLoUqtjgQSf/M9CxUlhVoBoVehVd+YszSb+b
7dqDH4O/S1pJeA/xr+sAvPVQw8WY0Ar2kqZ7XG/pRLjtqwKA2Aii8EDPuSnEnWShSWCO7u7Vlz6a
FzghzaaL2j74hXbJEPH7gyJfJBEL8i4pZ5tBVqTOo7CGMbSa94OWivS9fqSamuEwR2A9FS+hCd4I
m6B5vygrB3aTmLX32gyPHowM7xzjzpTax/5CLstaaVEjZbg91dRhoEoZCZqBuNNR/nRWI+WINdrm
SMR+c0ISqhWSRiCXXtAm61HNnkuyx42SXB4HC6/OrXGweVYPrPFwNy5RMvvbohsDCZfIcQSraUC+
waN8SEfyAnOk+EF6/VdXgAIH2bw3CqIk20F6DAs5pzLxn1IlEqo8d9v6/oE4YdVDW31gqIJEVcDk
BNxFWAkln7nWO2hT335SAvUSRGaXyjkU62RV1+lzPf1n/XQSDeTswEcDuTowmV2nJHtneOZLPiuV
A93oLQZE1Vnz/e9VI4eRyqwep0CpFCtcNx/rAjhHoWrZ+SDBvf0fWedR7WdkMoAvtBWpOPWYSCO2
BheB2HK2f7cwTCRxXC9zpAfYtaqMcEgGiZgKdrhQilrFE0YkyXPX7QEmv1pRXrO9Vgb7HRtNjp7d
3koAjkE2Yaj1v5YFdvvm5gZCKHNxytLGMQbv86qofkbjw9zO49PvG5kkQI3r2iMOjfBXvIaRqDkX
bYOdj7Lb0kZ66gFPdusjpYQa1o8fsuma3p+GR0YyZrMS1fXz6odnGQMsmt7f9K5iiZLur2IezynM
20FE2/ThshNv/q5EF4IjQDKulgsv/HjfsCqDmhH9M41fKtWwI54XUkesSf6ivUhQI3pWl7by3mh+
3MfjBdnFDStoupeOkyXQ6VUn7Siph6FQyHEoWikqDYAXcCzwjQjtIUdNeThngpvyt0S164JXx0m1
MMkcZFWZ3krWIyosBOFYlRQvrAI4bZXIhynP7CCotttf9istE2SipA1Ous15bMStCFFb4ibFnmxE
DiV/XAIbyxQEpbcgXqPiJy5jw5oSTx3vKEHAKKYaOy7Tu1cbFoaKdvz0Qf7xdagF8siAENnb3Jec
HJBFPMdsKq+dn+V7720x/KOgvk4kIAMlDxs+WztArEOeHTZLoohcvcolgu7LrzKchoRzCWZZYdtL
lYCfTmuUNJ2/Vk0Cet91Bi4BJ7v/CJ3NaVP0B/WYLA3SoOMce/bouMyo21stoFJXGXn2UKjEqmTt
Fr3EUbstv0rtnWUmPmqBc3grYAJQeAWoqa/sR8Se/Jmr/g/aIjYGMgdo83UdEBAfQ6ALQHoLJtWM
frMRUjP6EZzfLd7x+qZvZHjFNlmuU4+xYW7bZHPOcX9sGtjPdW4ETq51Mb03ApHjnsnETTYIBQQP
0TEiIiFKRaceDJbGGRBYiD9MWq717SQ5xMPJMm06VX7WhmUqNTPFfsMRgKeOkIwdT7SZgHfPUFAL
s8emFn7rjBWIzQjoQsVBlYFmgu0CSwYakm8rHFJkh7/Tw1Aw3Qur9pz4a/ODEhqwzQ1WPow8O4AQ
90m1jYAdFODKdbJIu0EEmiQTChZdrobUb2cecEXPuJ2wic/WE0ylv5by7YmhN5vStmQTssRCDqAI
xZWZHX3g+gECcUIObI44OxWIjPzsIt0NNLFQhkaXdOGVRmmpMWxyhbR2SCC5V8WyqOdvyiYgvHJ2
+0eTR84O9apV6FrDhTFrDsGw8jSHmVzeumZalGEgSU0bxqHo4aj5Q5rmZ9bQYY6q+r9jpGvZNKpg
9kXhl40rGrP+oUCGy49jftKnImLn51AhjNbuybSd2rUDLFR8evcV/OhXl9wnP8fFihdQUyGGPJ9z
O3dhyF870X2fcbVT1s6XOVjPqp/T/kWGxgWak5v/Iflu08//QIa604m3I/Jo3Fc3vIKtwIX7+NPk
ji0N4QYK3h0s7S2pSqS7m98r8OKIuIBgupk4jK1zs7Yk6ba2Z6j0qiwwjSPoV/qySzcYugqNHBUv
jB/ThmueYIkU2QRt9qTgfz9SSknUTfLzrnewkynlobG8Zf3hRCFiJ5i7RPbs1UOAS+9pYb8/cg5B
TrJmk4nc4j72d499h1IkMgBpSaTZ0C5wzsn8G7YjLUb4vJNbMgCTxH2gSEcIM5a4e2Cpz3yeTrSy
e9kIlt3wmYmCL+kPELGdRU0Wv1HHTGZ8b7Zxp6b8Dw1snCQ3pbIBK1tuldvwPBuU8n3XN4y6kQHN
SRYDGvvm9yYcKHr+UGywAAu8IKxLrGEBnXxhkKUUGJTQAavVTRidNklUvswkEVoBL0r5LhA/7aWg
R6QLYZBQachXrS00ig+D8V0D0xrq5Ex2wKqF+GemRKzvTA/fnhvPT9PIR9Zi/VkjC2iOAzfOFgEJ
JrX1bjeCWl9ALrWoHpo88NAg8TEscKSpp+g2f+WKXaRHavwHQNyO5TrQg7KRfCkPJ922ECQDb2re
wI1agPK7jDbLpPUSDfewiSAgO23GasVOIQfzLShcKheWXafdWQ0+iXas0OYxU0MKbOUEUYDGYDL6
NwagVjxbECFd4N7rfBYPvYEA23S4QbSgJ8ymYYdnGZBWoamfVL02FzJqbS/Vzuln/z0vG0BmvOb9
3wPnIhahE4eKWtLFkPpBR9+pLvnT+0cOMZ1QJ0v0KWBRR02XzdOHeGYLYBQnswSTkvS2H+pKy0V+
pQHub9PgPFKbUN+553vq8ZIvvxO6p3HiK3YdShDe4jCwrDw17lE2w9g3QWHHjjSoNPep3DA/luTK
ubUlfee/HYcR4nloGiUQT1ulyjpNcTw2m+292pvjXDml9nnLocjDAI+qb2LSpgB8pGFmmDmkPHpv
wG/H68KH32eyWNtm5GIf3Uu8S0fFupu9YO14SB3il0iSnxNYAhwi7985dkqXBDgbgDasgzPptgMj
sBCH/VzYWMs9O6XPs1m78obzqGpgVZn9b+NjOWd1FhAIdf2UpJooaqOLrwLGHQWwfxiFYL/pz+ot
OLtqycjTFuHDTfulus4ay8I9EqA5S6s/au6ppD6NVYmTjcWLWpoyGy4aMQ9TTu7nPR2wqsUF2J+B
rzNP76om7Jo1okNFbJWoWlBH/EXFIxTIUicD0RsU5sZAD0Co/ctqLemm1ZN78GCeuPNe9mYZyVUC
PTZr6RuuCyqxW7C5M8gLpR9eW5LU2ObNpFB53cDzgaZ5E93eUzW3Q1v/m/HR5KFGbVq2WJD9V0Sa
2IzHr9RLImh8gg2v2Zgp+DYacZlz5Ongf36XxZm3o0qnpMPy1ulKN4f0yxSE7GBEZ8juN1XoKAgp
U4qKWGzvMie6xNZQDsFQCB0qFcJUWoSYQBHSmglCRbdV4vsMB0QukTJ0KKtasqySEARlfUfcowhp
TEFxbu48UK1AChdOvzMDmoaV5ziPqpDpa8EZqvuRqWEZUcHk4jxwtsU023G7rqg5LVldv0R7pIZD
7FrA5zvHbJgQ0JtXa09dscoAHCssNYeDljvcm8vjioSugolzOugQXkWPTGADb02SX71hzdBqdpoI
3axZKWtIPqK9Vd0xhJ05f//mKsr+LVMhcmmivwzSIej7u6XA3EwvqPz4ef6V9Kuqd65xyYva5LAV
zqHRL9pPL3WERFhsa9uPTEMwNBOnz8oy2VbiqfsqQ/2Oi34r+BcWrtkQPdlYcjjMRFsgUYwbN2BR
tUBHfBpOEUz1zvbzZecLbDcg2HvuF8NnDaIZ+4hpUuRMFkpvyWnLWV8TjhSkS+LxXVSm3X1dIIl7
/PrdUzI/bju+Qs+YMr/ULngiQ6a7ri6kbHSZ79FY1xV3k7THapMOHClgjAOjIipkjS/Lj/pGDA/x
uBRO6Lsj1+P8BkddolNK0Y3HbthhBFis9TyHmmeI175bPAvq5iXjhH2Unh/3OQuAwQdDiCa89EWu
NQwsZYljQuAFKkGAk1vxj1msIVthkbzuOO7aV+hR3ujbAi8MYbODlP8/5RY0bYH7vq7/b1ooh43D
S5ToEyNmYXgcTAe8bEcCFWnlEPtz2n2Bk6t+1PusHXFtu1LRCBx6QjiTEZxyYMiemMUP+/UZ5c4V
UJ616EgJmarFFhjyiP788hFxJGKB3wfQuiVIdSNar0MW9OEViqgf4EqY/VaIJqAiWKVpO4a2Jckr
gWg7KrZHIfvGAtp0+jWaO6qh6mLDWuBN3XYuATv6/An5b0z4ITDRFfCeSoq9rrtY87/lX22Xhxop
Ie2oxfb+W09gOLLR2JNAQFk/wXnkMTVQe90PpbhMBZ3zfEsiXJwuwmLk/DevXWgnL19yiyZMA05u
QRoLFtAyEv1OsvH8UEmEwDA629hXJXQQaPPo45e+MhWU0XiRKpRUR6EeQ7uAE1gcaqe6LayLTNly
uWlaNxezJqGe/yjRgIl6icCiK/jMrJ9EcytE88ik/i36rRJNCjN63V2egQEMK5EhIE2ImFe+F1y3
0OLWv0mgA+uJNnB9DQd2V9yORkJmKvE0A3UZLpP6mbcD+ngiGY5j+mlcNMCkSsdcLkNJCgUa+8ZW
bmJEqzKx9qAkWJ+y67eVMtLXKWLT1J/P3qx2FM5lnENSyRPnAZpwBPdQSLtUzGkpo2BNzB/oZLzL
DX88g2SbjMaNuFas42/I+DWjX6aJ/mhAV8ayS741nLSbZeYA5Fpi2EYL5DF5s0LnPWi7HGU8WHXU
byh0wyJUxKqMCt5aiwTx7eYlr1nuKtKG8JA2Zqugmylen5FJoN8N9VfJPKHNJadPKCa1OEW4wYEE
fEm1k7kB2I4HyhMZSweF96ls0GH+aKtJujcDMOLPAFoFdYh90VvwvO4fZQTtBbUgmCsSKFC67bSr
lLTJxVoK4l41Zds2o/i9K8AiU0Tm9l5wFg2SIK+wg//FIDJyG8Ly4ltHhwq0/LjIX0ZhlcIx0xni
owYzFCDMhfyLy/T5Kd58Bv7l16SpATLx+bknefItrHHpo9TfQfUVGwJ0I2OgiOmYOrmbs8+cintA
BLiX692BpmHxkx/JvMsqBQiapmrPb3ZZuS4jLAte7T5ADpmBrMDlzmazZ3H2qdi4izWDYak4din3
QY6dWiXfMs7tNwgFRAV8ZYTHUU/DbASbqi+JrgaVnnGEJrO+yzvrvuCb6wqrbfpNDcTEgeihyh/X
zsenItGkf7ITICslMPbFVKaexe7ASoE5IeobRiSzxj0DY1/Lohfhr1k9XNTr7BZP5keS75vTAQAF
oyXc3YUB4dtt6DnqGcI/g04jMaaOTdYkNeS8g9Z3iLkA0DicPGPKbSPxTsATxOYMQujdzEqwwnlI
kO31Ibk6Qi3chtUXhGgoSn/fqmUm3w42Nzd+44DXkSvQ2sIUzDC8L3hLEMQYNF3DnIQDonzI53tq
RyrvZLxMrh2In+hKdcgGWJKePw/mjyBgbiOMvV/F4E2Ix7mK0m3YaBExiCOoTsmE3QAgh6X3gwVh
QO1HrFR+7hjfSUfWvLb6SPzRucnabCD5PTiZ5gOmQqKDt7Qv6gI7vxQYEapwMMbIYrcAIJamBKZ/
vmDZ061Is6r0T/rq3/y8Sb4NhTbIxD/6qudA8P7gN/Aeaf2gnuRpJJJ8gCFLUHzhxfe7qYVvprDo
Yf7BX3HXbJ0e2YioYd+8a7PfruNsuRI3uFDYZbb1ZNzhl5X7bxH4vwcqANobxOFOwJR2dCLnyAg+
9DeRO7DjYJmzAAjWevYKo0fyGKve/PWFBYXqvZkrMmVBrZTHtbsbPQV04FnThc/FRRlWFSxTWhmv
lz/QHmV0+ntzgFHTdB6f73e8e75AIUN0IAimq6ng8JU4zEv0nxWaUP0gKLOu9gR9SGBj6SMgSo7k
yddTd9Zf9Kzx9aDxHj4yu4ZeuNg+IkPWVV6pe+nUpex1Bk030IsUa2Qne72xRPXD3mxhk1hU8ye5
VJBlJqJzlX2EBAjvc5KcVHChbq8cDzoovoXKb6+/tVZn1/b/aJ9vUAJgO8AQzv/D/yGdSZFJC75X
xMQkwArJkeC3stAw6N/BXuc/MaHdFAVfYyEOW2BXICooJFubKYWwrQoxWp5UE2wVKPF9rlxfO/2w
hY8rMJ8vsVOU+Z+/HsuKsYopgJ2F05Hf7jg9SAjOcRtMuGJ5svg94vD+u0HGhG7ZVCvJdPSlTkGu
xF5UnMCmK8shJ8QUQcMQvZAvaYHKGRvH/S8iJoikNTPB3Wi0rAggDGTq4mhJGR9uZ4Tk7otTHQaN
9zx9gCISBVToHH2i/t1YFlNcPaj4zrMFN3rFwWsDjgV2CG+QkbUqLzndRQsOKOaZSqvMgAtLZdqG
GpV0TWu8ChlH89dGEJCBIbpVGlVkQDGckgEQ/UDb2knlwDTSJ8cl2EkOlAR9kBLOZT/4n/TCmT3k
JQUia5cQpAIvZfNDTFy/h2Hb+sZ1JnYeP1naUY4166UIrNKNukYpM7+cul0dFBcgIBRCUeyE4z3c
4YBJVAgO13R90fATIhKlvqisBbFkx8X0mzxc/bkC5AVR0DzcIuKEc0R3LfxIy41LpgE5j8lE/XhM
04X494AsCrIKPUsTUAnHBg/ArLFDxXV2sWjWD0dpgpn0Zw82B8AQMWJ7hsn4R9Ax/BbxdUcsli+r
o69/Ds3m2pID6G4TIozFZcKEbNGwl4UYRUWrefyoKYw/wP6ZwnimcUCj/JUwImAU37sd+6NLoCK4
QGPUnoe0bxPda/OzK0r1LGtLrKOmkzWlEo0BtP9gE5T1SLS2ucH0Fd7JordYu7v+Wr4GPITxb49v
WQdnVfvm6ViNBDGchDJlWQdqEq0iYFKMkBwiZ/JOLx7NBq07nm879jgrvPoeuCjiX+syMi7C22YT
/ZZ01oIA9Jxb4+stYL8594dVWCURHjMzv74NPoFjci0+vh6K9YqAUSTn0u8/yNSWx0/bzuHmKmX8
7kY+FxVvqz0/+ymavUELlZ2RWGM1wrBg3b4vkxMTODk3wZifwN2OOtgcEtgHpn2tkIkO+t2/CDcX
JQEaJezKWUap5sXxTUJaBEGpAgMVvVT9oRhfUzVDj6x1t1MMQuSljhc8BiuMJcRq58p45xi3G//I
oVstsY+b31fJI/ShZclPHQl0XwCFP4tFcw4ZMPlAwMVx8jhZ2al/L9ptthyul6c55ifsmsI1VWOm
pZDP3dppSwa9252AMMddxSiYA8Bv4Pgs5kLjbpb/uvmO9ZgzZj7XBDh59r1ytHqqkHERpNXtN5Cf
CcMdjZF72Ecxt5lBomDC9v4ivCNx2WAjMVhrqK0/Zvyc7JXXzDOChKuzFU2IhKreU9ffXXpqVLJi
Dr1Z1NpqlfWYVkNyJT0vhtu+2xV9hUGofh7odCnMAHOkOEIajd7hFZ0xuxQ20XW8IlUklKnsCJn1
LUAqdxxUt7ZinGuDNDlnlvNpHEdP2vc9Pux2h/Yks85kAeRSsA0OXi+OFCwDAvL1YU+FSn9vdPo1
eMUyIxGafUAeGm8/xF24+rmzu/RHOnPPgKdZTDvcvWIThSBy7xYAgb4uPK6fDYqJHS7FofbhKk7Z
Zvv41wMObP9+W4Qx2AMrf+J8ReuD+US0VCXDts73fIyNJRUT9a1Kl8yK/BArD1+HY+qtDVI6vcyo
XRrO19UlZKzBqe3F0zHm5HPu7KtM8ToBmNxPE6dQdNj+tdbBLUPYIUN1Qzc/b2h2p2F2rNgUyM/y
LRTZ2aT46g+WosP7bCswBbhnZngkpvqDM615k84X7Y7qxUKFjnEObUUTzomSKkOuaC1rHvY4aGkk
Fnm556Nql3Ze1DEN2P5YHOKSD3OmYydwIDn3ma7d3NHZUbMsDAIBmH2tT0b3Z9AZePSoqGxA426X
aqLILqS2U/CnWoOkryJjWnk/zdXtzrNgdw/NDYtRP6gdELgoVr/i0ridF1FdJ8GZNXTYueqazXjG
uOetDTDtas82wM8FBSDFCmGwZ4BdNQCGjObxkDhH819wIqDjWaE5QPP0YpBA507svJd10gk8pNiX
fSDNtfEqbmDs7qJ1lp0uEqdbZdjH6u/qtbSEdEvW7E6onXEozXfJBKfXICt0FMufzognZb9MvTHZ
PjtlihG5xQix9/OusfnF75Vnt5vN0jxoFjQASdPpmrDNyU88YvQYRuLeqaQu9fu6uozgInhQo6t+
KJ2pN0xDf+3oj7t3NF2kV2txFqndDXN9ReVROJeemWcHrf/wShizS7xy96Jrzs5SJmuSTECzLoYC
+EMJYyHls1PikdnEpPXf3wwWfno+2lE5YYWY5i6SbktiDED3//G7zz1DCu553BVo8I40IpIYCrs8
HLghr43P/G9ofQyUEmOFTCQsJjqwejPD70wN146y31QRsA/KQa9dWjFX/rX2hHejApH+Yy1t6R6C
zSV4rAryJlKkgk+kT8jGLV444E7O/vn1aoBXyDBwfYahLuGn7VMFNe9PRtbbKSypynXQQdAKYivV
NLjjGY9Hir4OiukMsGzMhh2CO7DPTAEkJ6Iy+O18XpKY3QDQJIbUIKdhea1kSmQdkdqrXI9eNP61
ck/9z80QNxjAy2rIVH+GZkw/36c1eg38hMShK55sXY+f+nWpSdKtALbh+QqUgcYmLLx3SWRmRfmV
+pSlvngm6rtvVw89/eKcTr+NXsEROYGuJLUVhCFr9w+Ei5VttSZaIaTihTjUU12TOFwdAKhEIAGL
/8KfPpRxtirxtZqKSG7QkjQxvtN20azxc30hDZIbCZRBGuPAvzdZ66S9iE++o6A6LlriDYCcD5MY
hmExqlmPXMQQtG9Ex7l7hgufbxZneR9dcRo6vrt4nB06Gg1hhbVsF6hy7BxXUZTaBJKGCnWK03/j
JYcgbSfa6SuNzo0k9ZH2E9Bhs36jknrSrjLBymy+AV7RgIwrz2LPOC9AM/h2VywAG9/hZC/GLkWY
MPuB5lThwYt3J6wjtpplXPUsumC6yimTGvBF0ST345KjHRiwYfNmdpiWAPPxWAaMnv6VOtYKsJe/
Q+7wWre7ULq9kPyZyy6DvJx1DwnOi93cULd79AkvVuaEfIC7rKOGbYjN22Mk6V3X+yHbOMIytBxT
NgCPo17Ls9/68+8pjYdTXOhm2DtreYslQfZlzbKLYPLFF66bPlAa1UEmBu4ytEjbf7TBQjTt6smV
nbBfR/IiHXHtx6W2DSWObpT4mHTkShM98NL22PF/ykMG8K6d31FdoyH80POAVgJh3t2oUlHS/v/9
vp5lelC398M7x6NnwwCBxjwKKV5y70538AeNOXuAEFQJ4ewc9ZU4dfCYXmtvS29ndsbjfX6XFJl6
zWDPYdv9ewug2hCW2h5yxSKjFuSxOz5NOEilzX09toev/NWoeQfSR7tP8HpBG4dVZU5bLgT9wApg
txXlyWaMiQ2hSzFpKYWZoI0dT90AW2GWokzH0yFTIIbaHfjXlR0IuIwPQTjb76mPlsAM7HnSHdSG
ZHsJQr1BHIDMYRw7vEkomo+ZC+VGAdH2xhNFWfW11ZpLNXf67mwDgek+85pAptoQuJ1NiPXqrTsW
Oo0ufsJm4mWH1RLE0S2JgRzAljRhPVJtLNymcnxBgjAsDZCjVsKcmd2UfpBsT04MTBoiQIq/3cDq
5fyWhNyGSnH6eX+Y7HjLLqn5UCM307atHy5cP86ZffmUV/Jo4BqSKvb5vBfBZ4ZUduVfSZNtq12F
BDxa4q4hyrQYp4WlSyxA7kAVz6Hw8VZRulQfzh01jpbldz4VX58DWEpJKE9ntC9x3Xg+9loiOv0/
UwK1REnYYmN+eini0QKUSv0g7XodFE4CmNBvNvvgFKd7wRm4klYqsBJXP7/f/rkj3bhTMgnTzUHc
gy/yjHt4mCK5troBGeISLRJdtVF7QM9IGqSxNDXLinUKrSvlm5L3Cx82FEJM0DRwNjHbY5YLcGRY
LxcNFfO1g4MA2lbXb5ghVmxKAQZs91yzjTCr8ZMA2++dEUkbvKFa+YBr8kiCplMbyAkn5kxQyw7p
ebBKw7Z2tmNaixDSiwYzmpfZo1dZddShIERcj/4yBonAwfRGRIvOpTK78juzMcCuvB+8F6/q+Aic
dpPqDq3ZJi4V5yDS1zwPFEmIPHZXqsReCouvJDQHCMBgYMYK3ZbfN7iNMhUV3FFYkgKzQhNnTkiD
YE1UrIBgECz29x9xUmx0JcKHcXd3jACwme7qJNsLey9cXY+swKR19S+QrIhK76AZ7YlWj82Hq+ZZ
OsMcx8hcdcuNRTl18AWDvceVwcP1MxygG+vR+rWw9uI7GfMEUpl1YIdJSf/HqWbaPPKXeoTCj+3W
AztTOEgPH7h0zvcvipp/tl+N3M2ieBUDH4r8BTCMh1j0ozaeAjKdfeFHB+I43sA99QnMr1pcl4U+
CrAxKpAONQiZ52xCRFKt1HD17lsoNOH3u8UkVpiYdRRYJptkiQh3HvIbcU9qzUtujkiIWsTd+z25
FnkoWde/8vrUpi5uiKJiecejFdl6yhJmDYp7uetudBgXE4Ssi4QxLzexjtnVIrUyUGayxGJyFKoY
UfbzK3aA80h8ccOr4tz2OaK9MXmEaCC6mifmqCKPC72IfXnEOhkfoe6coLhe6WqKe77QQu5REZyp
wgE3epEGSYqis4kY0BVDg3gLt6e7peIMlw82LQQWEdgr8E11hfqMg5rI2rxGjhg84DNIo54pbgUQ
cx8bcIcdVUrmT0VOuOJ3noY13WWm785CjTmZEtrxU/cBt+l8YA20676p6gz7emeWs6f71YaZwzvT
pnLns+puvtEBp6ItT8RW7cLmdAe0uK9LfACrRcqrQEPFpe1kldMZk5yEkWqmwL3w24W0dfuyxeLM
RYNMs1t/uku9rGBuXYyEL9n/Q9vd+ZoBFDU7tqrPqaXB+9Y6Dz/EU3vFeYg9TnsQwvoKezBh5s6b
qXHtiquMltIZtTFdEHtd2Y4ROpxz53QC7aLxHfa5XBdO4cp/+Guje/PpAPbgQX+pbSFPGazsPAV5
VDGTZRkO9xUt91pX+98I6BVT01AOUWdv3rcofC0nKgUMQfboFqVOpi1W1py6C17jsWTkqAPLDYPd
S5M9qDtBoBvxYlyXGup4fwt43iGSaCMQMh80bkc7vt0DDzn3PhliACmMfAzBhpK/4FdQKImUhZbB
gj1czZQ45dGbyYnXsyIAW+h4E31bHAtMQ1XbX64dmmEHe7LxB0A3QS5x8xfxFSfH0v/RnucriCA+
9BvxK+VMn5OsbfaaUo8zfOnQ9FDdT0zrgGOCKu26jTLrwb2G8bfMb/DgZEhqC9bZ+h4M+b8OtkQY
gWE07lhpgi8FnV6FIZV020Ar7tfUWuJlw+sCSBkZISGSffe6/at0ZjVwYD0/LF7OfOBsuBZ2BGcj
bvJwwX35EYBnTmWBUXETARrQlmxWF1ZjqsJgs9OinWEq2/Y2VWLHRUrp1DSnExfP/4vwgPPARjXF
AZpTLuhmGq3vEfqaA9yXGVyoJBA9eOY2D7xOx7y296LclZWTguIeN5GN5lX+PLdmvJWTkx58ThyK
cY/kIvyYy0T85jyRL4XIE1wrcVcMp0kubld4G93ygP7BF+iJcknfwukQCk0MA9W6hoyqt99E7Ksd
PEwLN15neuyLhqJ5EQTxWPQj6MK5Vx/cyNx/V/JCDOGs5OmeAjJCPOv/64noICbbZ0fFMEZq8U3T
u8a9k1WT0C/9Rnm6vIfbSOeeEGBNI9YRs9EA5Vwb6ZfmWo7K8X/Kk6bG81eFmAzr+3bBVOZm5NrV
MeTEwhEm/WMtFNOLwh5rAnO7gOcd5u3TWqGAcXUugFId4Of4pGB9EI06hk9K0nCI9IrHuLdG8Qwt
ZX9mK4prgpHM+gXxpLvkeCN4tRxQuiJaperpusw7ajoZ7hVIZDwVfCyJ/q4rK1GlkDsTqHHAWnzd
6K0AnQubqEQvC3hilCGPACFySwCh/iiroClDj7SqKdzBplx6qktPrGtW0mlyuIB7ghM7KUWDTNqO
CTUMhxaDuedgNPQ5Sdeq985sLIde0qKeHxfi5MtDW0MWxMqdxxCRs/Xqz2s0IZSHeuVVMDL2cCAb
HzQRUhdzMz/ZPkpx/pREe9qA66kcsVcrk3xS6MiCOruDoWhO5OPIsL+L0S7OpM+Mv5BtGBIuq7tX
aK0LfZVA1T4mlBOBobPsTOTLkUbHyfL7oJFaEHDuUt9Q9V1XmmKCcHnoB0S56jL3MqXEVhFUnPxc
2ZkMrOMIH47K1PKdeHFdgDZ55Rpd/4bE1o8be1e5/Z28D/2jVc+FTyXqWhA5AnqzI7B/vQgwJjpz
PIEEUNwJYogLfFTDos6oFSHwDbYhz+6gy9s2k1/BVt1paqRM7M1NQAG1gkzzpier1N60RqgkuIeJ
sDt3j2fbtABOsF87bXCrBAuBZfRuCOHupKBPnUiwGcrNZd/LV9euMLStM8byqi1EdN3wjoeFIXkQ
ANpxt8MhNwsLU0pAQB+yX+ZfizRaTvJc5VOLyk3iZSyWPEzNa4yZa5qp0Qpo998ZraK0qERjsB89
adehWTs4xIlwIwNzAeSDLs0Whaj2jeUfIxtgtG8ZnD3t/SJYfp9WwUOPepodOhdMVP+doAcWlsxk
JrY52Q09jwHfdIJtB0pmw+cxDZrPqcIZPHeA3TZYvhGXILUR8yfx0a2yls3IyrK8PxArgtfOSgW/
5ItQ3QV0rj0Jbc7zgEuVkrk9hTkIJfWeQgfQgcj8pkIqZ0EFVH6zppwRKcpPcFtBhHvrZLVnY3pL
42clnmwXzgWXvN/KCtMbtoWJTIbJY1K9lAzLmee60Dq7Dk+cET4tP3KEglLGlqkFdB0BYV35N1jj
2dX2uwdzDU5PEBg5RgUH6JKjTTnkcLE8oISHBlZHaj2hckhOqnxleK/5lNUkzwFJ3Xxwlb0dFWwG
VvgC8SxLJ4mChb3+6QHchIfEeX1FgzURAaGm6hQ8uEH5eDKzTh5TnImeTMoLKS9e+iBVPUYF+7jO
DC5CZJ5cODAyVYesua0TBgcg1Hva+fMAjhtZ4YeGyzHvjTQt5U1J4QtN5NlRyDTyReO7/G6OnCiH
VZlSnK/ckuVGJzm2wIzs9X49z4TSpA9cZC8TAqui1+LWrjeSQgaqAoVlYhmKOjf/zaQYBV+02YYN
bdUFoUNtWUsMKdgFnK70zUZ5qKeb1UK0ftBX5bscHQN4l7Qz6CPECf7KibxnQ41jjIy/IzRIZ+dz
Q4bVyymWMEEOrdqoMyqQ8HTlUNmLgJ24EfMt2PyfQ3Hz0hCtsGqx20JFTqtwHdHWqsyZPMETdcaZ
SM+sSwZhUE0gBRQyH1jq2hPDaWUuwhe9HeI7YVh3hP9sB//+/m17/PK02VNNxhDwSKbVkh2cRtNo
vnmI5JV4K7NMtbV53Zc9yS5IJw/WMEaRf53U66VMlAL6uS/YXl5QYATsu6Lw+X3mYdbbXbskErTS
VpooVyclgDXqObegqnOP9BtaEpCJss2Ks2g190ZwdCrDApPjU5XaQMYfi3eQIttuo5+UsQ64RWQJ
+4s83itRYlMeJ7Px9nkZF8uknTb3tvNsU1/V8Dtm1jXaUIuSxEdKVuB5rQ6BGBlRVznidPOmCEYk
+mEKnXuM/hG8590CwAB+WBCkXA66MsqC5pnf9mIHttsYmZHA32UXmu00AxpnCSZEFCzQuJZqvalY
yO/FYHTmlYahKoF7n1l5atr6BeLbvuopxJaXRLTiK16uSgzsPZFOKSvQaLN6B34fXbrRXUr3jX8X
R8xDzpYirwqOzK4HpTlthPby2fwsl6Bh3zhrxdDOLwZMvaIotiMmvXPpt4Hormqdm05STJbYdGQs
gXxIhS8adTLL/NkSHi0Yr8MaOpyBgmkXMC/8E5ecvAnMWVoOSWjtsqMMlroxntV66DB+nlIPhUzb
htnt7cBHoB1NpPQskiJtSgCV8SEP/v4hvQq4k+0oEITa10Q1C6+ozBUP4aS7AGU2Fz0AgZ2++EQH
2dhBtGSVWmO8MRlEKRLYUhE+ciHwHcqx8TF1jZ59GPmOeRg9z1L5d+7Rtrpp1DBm+W2yb8IJ9elf
5U2z5PBojtJ0avIApB94kZ6PGX7Zg2bZ4nwG8IE3Km9pMKhriFg3Q9mcmpCT1BaRKUOBm+s1FLWJ
GeRxTbapEsVKV1oQihlaqNN6rc4I1JQuWjGkkrXCZu3Voyh069drsTHOT52La0s6UMNk049GRNPm
nDfHekM5+FhF/h2iiv9HUgtCW64jBzV10718UeWRAdREqs1Xx6Zh+hvsiJxcMgtQoB6hHc50AZGq
/zHqCBostfKEuuA/f3KfchPEvALpW51nHcuuBUIXOdg2ZyW1+ON7i5WsRMdBNcS2tVHMfskcLhwJ
OWHN4vuP6KxFwlFeqYdNQiY3jExrHS0CwdiQrUjGss/sGiemttr/39/8VIWLRlQm7/IDGPOI2VIj
TDISeNDWCuN1xo5bIP+ImROfMq2c5c3Z1JCe07Dir8+ZlEhtpyn1qydESlF/VxfUa+SNvkLCmHCV
QZx7SSGHYURTrxWq2pXhALJS4+HgBMQelrB6HSx1acAqia/ai2yLfi7RhX6jkzIOynjUABx0nIaq
o7L+9qBQOOErIgtxrd6aZjzQ+h4v/1pBDNu0m8N/K7o/xZY59SRpX9WZNUNjsj3ZNu0k3tZ4jkA+
FOigtaNFcj5whRklzKXOiurZypH68kM2FOcFHspmsQjPn04np5MaINUFdL0k34NajFbOaixFZin8
dihzSgtQrrQ5D23Elm2iPaVqQF4JtMLOFNNQhTH+QXe1le6cKKYnVfxJceP8G6MBlRg4a6EEDS/L
nkVGDDtYNuLfsrZFjfAKcTFIcd826Duvmfdl+BS4n4Q8S/jHIxDr7OlIBti+62791t4Xuc4mn1wI
5TFO/pVbV3twL5Mjq2IKrunPfFnIo4YfFgaxKd0BzkM82anFbLgpplMC9ZfbV2DL+t6S6NuSU/5t
GiGa2AhypTKFpo9dXGUbgnPDwGmrYaB9JbwwXHXMWhPYkFM92ISXdCqJavBRXMiX/wWxAmiyoQDS
NPR68WXtWTvvKfv1PBzjYVQUV+tirfvAs6TwPwPPYrPj7ZvFGhxLBYPDFFxyNrEf46EIPVJZvuh3
gSaGunPhS4wkAY9aSzbraLjeByxmSpNo/l683QRawqR3LW4f3LJkxKPNGzEgMOKZssx/c9zVdT+J
QE3+FE2VspHz6tN14f3/5hYDSiuP47Fc8MXQeo6yGfg2MHGD/qtlM/7YRMZdotK96gebhCpyucWB
P+KObq48AxFlSdUb0oYvStQCCqN6q8pTgWsndhMM7HxlfjQz9c0w0CYorcqe/Xu+OUg0qTMRu7lm
JHi/O/k11wjTXWCva4ptK5HxBMwdh2rrLaISrnlAzhGbwHeYfHoITBtrttHAkz7bFSv/07TCRVJM
WLGuZU+3sspWAD/Y4AHKy0wy7FRUWxin1TIdRLG2p0OFIMfSx2vt1ie6z2tgIiqaToOjGg87EVHg
A/Ev3mEMeGTMO3FhNE0YRpQU0C+cPtpfJ7Nq48Xunfa5m6SoG/zbFC8qxAa1u2n9SQeXE9ZYa1/Y
2pEmoDanXMcrZS/WeqDN+khyrWNmEIiMwjgwte8L5udHQUDolaXMbC6cWbu2Uo+Ya+WbJYXjdQq3
GL2TyUdTzOJrF6qEnI0H9Y7UMCTOr0lMG5B2kXzA1I7ceLEsSbUJ0Xto3XaI74/zY92zeEc4Rsi6
CgtQiw5KBZyxjAJwHmQLcFK55nVgIwyAYoxnX5kQywcUkZmsIab8YAGcEkj+ZfwJ7Ar2MqTNK0KV
tf6EXIyNuDevF0TJmJzY0GBp9OCE4YRpQd07oVM0rvOzhQ4j818Bj0tCMHQFMf2a5ywXP2NUBK63
SAoEGlY2o9ALcU+W7qQ+TLi5Y045j88INvsQRDkq4/aEnVQkYPEj+7Ou7rr+uI1mzE1wAL2HSnap
cN9UmWzW1Ay/LoKwxTs62eGkjpRQDlrQTLDqykMRWpZaiMBwLdiiUVWWU9/W5PZnfBGD1wBSee5c
PMpZ+D9BLXBJKUWHcdWH9BRWOkixB05oFWftRCHtlvaiNpJ8JH/zTY4gCg4bEb74jSqhqHfO7GLu
8OrRxXBTLwKJ0K5yHHhakzGiPW0EX7bYLCev3G9yulcP4T7VAjoPByrHJ6V2uKMhcdfSirk1CMTK
sdK5hucn77vP7mGlvPJe1vys1wOQ1WWXK4sqCFO+iZh03MjI+mhS2dgPP5tduZAJY2cAP1779LMv
9h7Ok0ZqNDCd9B53u9nv/5kv2XRPEQQTSmOt4gdfALhzzLOuXJnEEfj/vJ2UH5BjGP5inB23F80E
VSYuiDDO1EVyKUMy5/o18RSnBu0dphYWOYGyHmbbv5Oce3rCCS0b4qzudKK6FEqS31ABcUoV2zs/
venDWU4/fN5nKnyWJBFuAgBADY7WtYSTi06YFvPg3nKU+OzUmpqvpIzTZ8qWjslym7IB6MD4gv6S
MJT1yWyGf65JPGmKlHB076rkbOT/bYYM8086AqRXRFdF8xWGYUNWJ9S7wyQ9TF1fOf08nInJi6Mm
ooC6Q7c4gAHsiTSARP1OCXvR6lcbYxRDsGWkE1pFHXvdjQZSKXqy93474VBDHmKygahEIvtmTQLm
tV16bMK66IaDYR0INX1V/UKy9JTc3xt1OglZvJGFDiShNOtr+DfLZLYVhhu3Y8XBfKJht0JMueeK
7iyuvGabpiy4dzD6njJXdEf2xFicacrNq8dZ65m3QNla4VOxZnrss/K93TX1OES+26WtfJANegUZ
s7vvE7cvE3lnrrqFxFh+R/R/t4PjzPUsLYJ6xF2SnzcMKjlZlyVoAdPCq2cNTMErnJCzunaexSe8
7fQhV9yTf7YYenR4wnZW0/OxAiHhxkr2m6B7rXzwJEaEl7oN2T7FTEd+8o5gIohPoOhO6iGIVpN/
zWOvpEb6Wak4yk6eHwWbAJfk1zr66YL7l4LanttjfXQfg9Wsg9AlciN+VSDCMr9VodB4BXTtctrT
AlRTeLfFmjPZeZrzElDxssU0WBzhxq05L0DIoA+P2d5BlfJNqEiqx1ionb4M9g8i/0uyFdXOVhUw
IJx1CuIGz3ChbsLPuOCO4LVb4zu6Arhn94rERfRdG9fVP4oob7d8A7mJC34IfNCmBx94gO7mG7Ne
Oan3yiF5onolEcMZX7rLhgCbKCpaW7Sa2DnoTx7QoPp2HjycoZz141pCqudAomTTywSLs1knGnF1
2DgkE67Xxn26ibHvPa+Lfz/EGRB7hCtdhjSzKAGcf/mnFSbVIPJh80BthODU3rD5XaBIvSbrxht4
eJkAN/fXV9RprCCRMo0pZ2jM9bs1waDyorWjcOe7r8pW+ax+BL6LDyT1vfZgeJExgaptDImVcsI4
ENJgl2e+wm5iMBMFTDsnxltpmvDri2YFd2Pk7QNV52OWKsn/fHu8NcJ8hqE5ggVVQDcKu1fafQXW
AVx2cpz6H2JxBMSclRefyq/WbRAcv2Rgz/sCqpGC3qbwQv/JspNUhiZbINbxQtL566eZg1RVPbaY
GPJ6ke/rX3Z+W2AKAN5xnA4BORWk5yn48Dlh/hbQwVEBNMSNk+OHQY5Rp4rbWs0jRKlzRw+zlC0W
U7HduHVZ77hZI+hWU49PfWZ376gbCpd4NQlnZkBwYnq7Z/4MLifBccezjklE+8Kk3Oz8xbWTz+QC
I3aBUKkk4yCzA/AULmzvE2W02I6XV/ajfgqFqHFDJ0WwQLiGoyX5m0yZuJllDv1dxDR9hHn0O4kO
d1y9AUkBt1BEATUfQR+i+nqDo6uYvGZuF+D9y2QNnabB6RfsmeuuI1v6NdCCEfWoD/EG2LDyd85l
7Vjq4mwsrqsSK3Oixvu2INtC/urOABIOAlHw8Qb5dl/I3dj/mCE8/WfcYUtr/GLUNFrl6uWf1v86
1UNTDA+PZ3ApZLlNiNO84dDx0PwuzqYDBhnYHxpdnFjUP2NzpoWPBfIuFZW4d2OSXbWjE+FmoKOK
8N3jTgwBjYBRXG0XWBtSngUEz/l9gThT6y+65a8pIVt5+w7G5AKAnIDOdkn66oSwSBy0KCiuJnsk
K+Ler1x7z26H192EpyMYndqYXJnWZgqsekqsvmFC96l9YBSdI9EVpPgvOe+8DFvBLReMmQzZq3Bb
TC0N7tcIufzSHtTRMRkZEuqBbl+HlZASp4Nj8kC2ZEbXSa7fapIuM4p97QOyyWuIu69Q4dhLhqIG
BYUK5JBVGMUmjG4PtDhTkuEhFLsy52BGMYyu1vZ0nSmOVhE2k83aNNeA9NcZ78mJSR72vM0hPZxK
JRfvzPWCiVI5E1dVLz7fjxJs99t6AosEBAML6I4uDeRrRnDq6nZg+IEwnggkmgxDHekFz7gwfnjN
mOzA2ncoRP8W5IndtUQYK1olj01uuAuTZPB0TVVtIGZngMCpU9V5wo++0hxFo2rUvIPANxT/p4Rl
VTjkLrH+wHEJvjP/kEBL21QYZcMT+FMJcAMQc/X9Yu6Yl/iXVwBb1tUnkRCRPz9nj9VRZnYSwceX
d6XR+UK7+gYH9oUmhTvCX3z9g1rqiCpkcpwpVa8oOJbfymRxMHfpE656fu2XN0jv18RIxLyGLWvV
J1rww7372umDqX0idmS7K8tyF7Sjoi4BdMDNfO8TCnYzE3BF1IjlPsTWJItRDqYL1jaVL6RRfrkT
QKjvf8h1p+R2j9p4O06EPe8+h4RZGB2nPq+wDs0rqj6C9/OOLvoDOFrF9vNWU+lRSItn1x8ltjkH
Ci5zqjWhGIThy1hkh1XMXVWPDOCuGxA0IP1dUmOSfbpt7aAcO/xfp7YLYaOsLNiQN2EJwbrPpUS/
k+L6VNxOM/kypIBTzZnnC8fDYpMW8OaJKhujqHMf1WMkeEmbUGyXAO7zb5Z4SN+K3fx9cHFX4vrZ
pJ4Z7mTb0Kz2/ki0D9pvV2RZfG/YB4iAZ1TzeYPgxpc5o0Ib9LgMspTfbbVfVZlSPioJORY03JhT
hI93McdEAcWd6oMaePwgOmXurM3vMCqv2vl2rmDzqsmwsDqqWS5dnIo/mAYK3HQUdHjbGf2jbXE7
1FmFab3SJQfjnSS1hq6t2hTp0hXQ3BGoy90ahuDU89u4KwYvx6BBtb/viMJkmMDOvQN62ebopmhS
q25xey8jjESRxzX8F8gPOhazgM6Qyvkgc9QGvN+zzSyzbVPEucy2lTu4uD8uNuIRIOllV3bSUi+H
Eak5DWBTU+lBUZdNciubzUmH+N5DC5Neq7iWRdwhCV1DII2uK7ghEOrAWyzYmgSQD83Nozr1r89S
QLN5Jh/iY1oZaonJbmJgpkxIMS6UqFe4nI+1e9J82o2ZeG80Tgac0cSSb5U+uZcp5pb674CjzsmJ
xHdOgVmhUfWDnPUSCFWFJ7BCirjttiQq8tyHb7pUKwCwvQU0KjnDJLG4roGGxkrwl231dr4vb2RN
CcWtMC3srFFTOxsCmltgR5D0stIXq5FXmTWMLQeS04wC5Qden6XfXXlazI009fwIa0TpAg9y6y/G
XRizhZlonRPox5IbtUvb+JrsZm3GM7/mhoyDmX/CJWsPHEKL3eY4zIZcL/EVne3xoITCj4+wRAzm
5Man6df1sGttuzNoD1R1/A/nTNyxtiPnIhUXwVnJI0tkrzRm6xNI13l6GP/WeT2j8gz9Nv/57JHK
B7A1PWafp+HXERnrUVwDBIfDMIgtcNISLK6YcOnpC2om92DsQsRHs64U3JZMbnJ7by9NvuAA1So0
2wMsScG/mn2YhdhyeH4e7xYTSkT1ZoomUcYgbt+776jRkHhk4I9rgINSZFnOymfVZfS3IQyJvGa6
SBCNyKGQ8LUJ/8K3wm0XM6yZdaW4MTckWwvGebZd4LS2A/7U37kMywGfkTfazYjSDhRczhKMUx+3
PWhaRB/i/44csY04f6l2qOlFJnritpDb9oxvXbJkH2lgTfijQ3mfS7OL7YNiShC0vGKSZqy0J4Ut
mQRHhqWfPHMQzeTI7Gcacno3KtJQdUbdVO1PZxWWAUttT+7RDoykkCiQdJpXdkyQqlAnYdwH9j1O
eBa9vBDvPHrwM9cLv9jtxkvWnSjIzeczC8xNrcvBF4rMl/jF4U1s7GAwjTAHy8yn1ET6KSKwObTk
sDaRde6k5KI0H4eYhzXZXSPiKO8OD0rWdjs8bf09Gx37EEykXexIUXU965WY5kbBbE8vwCm8xIvD
jGZ2DMvERejCq+Z1uzVcaeQUggxaoB0lSi8GoeVxzHjdRbtllJ6A1thgaQLmLizHcXxaVJk3ui6J
N7/fPrMjebpLHF+YK9s/UULSwAMvWtfpj+P41cTHGVrLKo8fvpVofH7Enlci1KHeGtj2sEjyDNAs
WRXDZ+zJHCDFa6reECBRWM8xrh4XrmmTM3UhA3gMK7hjvHiqfehNVa/F+SvWU8hTdcpbkS4FtkHy
md7aERaHUzgctxgHpLV9XWt4ra02kX/DyfGasGDOjufwzwR9QHq8dokqUQ17L56IzZP8qndHjx/6
W1O9plQR/Gb0zfvSoJ8y1XADmb+Tuq7ELTHMJPy8SrNkjt+OlZOLBSwnDP1EoV6sM8asMGxLYGSd
wEw98l+dQL6w/1/gq1bdwExwqcxw1g8PC5erJWcuY/hy2fmj5RqkOIwsA6DEJ3zMKYlD2FTfsqyi
jpYjP7DxkUu8BnpydRh3H4G5GNF1eUKEPayjJodUnk83mLRWACGNPH7z2y4NFZXUCDY9Th5Ml+6/
BtWYBtiuhXT4njKbmD4z9KfJHhdRWCNdhAeoocSy76biWG3ubvoLoK3Qvkx9WnKJRzqE9xWhGhEf
cRJ1REL9yYZE4Boa9Cux0jUzfZC6ODK/EeAUd4bbgGy5hkEjVU1i/wW10gC87jrFKea98A0ZPUh3
qHg5D8T+vH38sE0BNFeFkSrXfIb6Eiy4hVe7umIy8WXuc0GFJC9VO6gK8FnOH9dnSCj0aYnsNAZI
JcMxfB0tdZwgxJ7laXL4WGXBy2+7bGjvuiNU8p3QHeDNXscB0BdcglU+e0Wp2LX1NAw4PGc11On+
FZp3ZVXp0XX+vSSae3sIje9Dn1RYCqaIHGi/ReXqYoqOOCyJecl3ea6FD9UFi+isDXd0b1ZWDzSq
82WgymIFgliIQ4omvwwDfWeqvcJKsgv2CHu1FvwQaH0HXD4IR9oX8TLJHqbQY9fzpiOxeB8E5y5v
uNmndh4Py91i6GStWP9A4G58WwRuVN7IJPtvpmvtaAOlZW7S5Hc8G6yoOOlS8jAfin4W+tiBwAdB
zDj1OXJOvxvLxdKkMmyY19lPJ7414FVvwGmHjx5Ia8IMY9f1KDnX+KYURFgl8necKxwHrzexjUYu
oHlGKvUExTu8nLdMJnnmKkLfkCWqJRR65sHbzGt8IJgDm2r7carpIrKBWT0yJpcM4HT3RCDXV1rz
D+s0EP3HVz0oG6mX/fK4zJ0vQgnyr4Nm5HtSZ0upyHEfhsKt+aIDaulla2AyBKcDnO02xDKfDeUp
TiuKpaJ9iVzHkPi1EApornqUZvw9p6pUHeebLUEZ53aHMlEwr0iG79ilvtcZmUSKqTutmbyqIYBk
FrhXyfbIU25H5qBMIVwLm7Q1JOE0EuePGoXTH+puM/hUNh/EDkmKygcB/Fv/cU1nKGwit9ZWGHrx
lqMr3VgSsQ1QwrNGK+YMDKAFolrgHKidUso4djUdHXy9lIlceR8Jz4AAYO4gqL4ukd2cZ4l8BzCN
qBKGH8xWDm6dIIoF+iOUd+6b3OzljDV/PBNgRYXRXMK3vCR6PI8Y7Tev6mM4u8S51S8x8VDV3lH7
oJsiksF3qRbW3Tl+q+UN48SBmermKkT+tFMQC3OZCusZrP1mvhhDDuOEMsf23P6j4rcUd5dKHODN
D+cIcykL9IlRKLFOIN+pSgb3UFotewAL2qULs9CK4kt7BQkSrsUfyxReuNFUlWVFyPTtxQAWUJib
+E1webFNaGtneKv63aSaqi6eSYXGEW2xkbO5/0stTDP1vdtHQGojM1/rtx9jkrxZglS+7KPfJ3YY
eZDzpvZ0jEqERJ4R6kKc3kTihagLr0A/uSdL74geWzQEGmcVGT7r0iJz41vT9Euk5X4ImFc3k0q8
/6zmlVjDAQItECX6BOzEdNHhSABHdUEL9UKJgGKrsyizKXnZueTTCHSSEX1REKfKlyEM/WMOY6/G
jFajRY7QGUmGD7kfrJkP5m61dZWpw67drYmY1AzQn+uobfFhPHb+Rcdvx7+vb/zC2vj8J1TyfmeF
7g9WQc6mqnyF+ZmMMAtMiToXQ3oCk6W8rdx6CYBH2fja5xhkPtx02XtZOXDGS8KkmQ3cZFoTfWW4
arhVPP5nJWqCj6luLBt6nREoyrpgeoC6Y6rQ7lmIK3F019F5QM9GX571ySGpG5S+1k7YJ1mgK9J3
2a8zl/UufUQdMKjrT7JqIKF5E3uHG5EjC/jyiOVF7lrPsHoqTZG5MeJHtVSpCskEg/fHykr4ANUF
y0Q0NPY0y+eeIPDD2Gx/b3O+vPvsaOGKfJEhsVfO0TPbZmP4KTQvJXpZBOuKCOA3+J8Hfzu8zipA
P8gkzdRF0DdhovWr95eQKxi+//aEPwNMc67kQeplm7KrrrDegYEZHfVrY/qQStmaw+FWS6z5FgZc
l6k6LBO8cU9Bj7SWN6etmltWR9DKNlPyZU2wjAKjMP49FrTm+z4QmU0APnPvMjXk4vRmBOxforh4
dUlju8KfD9ZWxsl7sL89XDFi+K3ki7H6fDfjMpvScJQtB+iSbGeynKs5op6iubupdo8g0ZPf7HEI
CwgcK39jpaY8rRxDBZ/7+P6K3IBPSTpjpTcT8XtRDqlKJy7SIJ+5MRzsuX/BR3kxLrUhCkzqBZeo
38w664wBy00ivVnHQ69oriBP9qE1t+cOi6MYNB9Uzvit4kHXGyuG4g//GDvhLWwzjmw7ebWMw93U
sVDQBHED+1Q7Bp38oZ9rg1UuEYTQqjy+iqnhna/Gl1G7WQfXcDI3oHwpRAsvabWC0Ve7TCLw8wuL
YdutF3zyH5mrCVMlpGvinHWcvPqLKWwFE/1/wPz9X02TkGo0RZzKn1/wHMoAjqR7OX8sTO97TcIz
IbvGQ/gEbFA3IOsFhfHoWsv3H26sJK7mKbTThyZ4NacqgoSn7SgaeIR+95yMccQUTIKtnfaEK0EV
fTEy6lC7fUWlBF0kihneXWOcgRmuGfP4iqk5tl115L/BqoveWCW8LNz5RdbcbVibAXqv/jkdNM6w
wTyGI7sfPeglq88h4kmnkcTX+ynQ4XUUHcTxIBIALdZzueAGw2TRDFnvCoFPLfCVzhJCA7P6RBae
05TzpgLx9i6643MOKWgmpYQW4VXBJRYWN0KxAXtTVamDQd3tS9Fx5AqZo7AfrtDpqKzwLmubbzwo
cRcM6zy5Y3d0DYGRMKg62d894wlcNqzn2an8ZcrhdUHV7PIk9yFDHalBx5fkccv86UTMCAdKQsIo
qGTSHIqBieQk4ovDIWjrJmaYZTEIWT3/IAK4hID1f3iCJQvbHwLwSq0I0o2N7ZqZAvQ6rw3OLp+S
PBIW0RtA9QB/MNYmvVB/HwMcSJ4rvT77gmxr9uqc/Gtg9AnWOytb54TLJ0ZATzvSRgwR+hvcigvi
H68cK2W+Obj8WgvLnAWRLh4FtrW+SMNpN92YvtnjPIkgyuSL7k13il1zECxE+HstaIwwgUa9Sczl
N3GK/hXaW4EEFSGQTjLROpxOw+0sog5IdSE3c/YmYBbgt4ytI1kmxvnC2HH/L12EglXCo4+GDJE8
Ve37iGd64iw1xI6KfU8kdRggVJrFAS5O6GJvTZsaYns9b06MR7VdUZjz8sjxSXOwP+go//zSt/G2
+tSaaKXVS9ognoZZ4//nRLRk6C8i4trYWfOJd5Wl7S2Z56ZSHX408qROzms7y4ZI1tNSJNfWeJ29
oUtz9nQMl5lFquGgSnI/u5RdUHW9BzpXJ+webxqNWgj7P2AaN/KtayNsu/GJtAxKQXVjzB3v0P0L
jJkMI2mUSHqHDF5XpJQiuN1iDcLDxtzj347Ezf44EPgXGEzMFcVZ+Te42jpnaGNzqA/YgzZn6V6q
F0j4aEEcjR+AePkNfvsdCVYFSs6h9OuZhhovqe5dql1IGBliNrRPb/c0c7HXHsKog/vtLeFvWFxk
Cx66OL9u76bdSjct7L4LW+v+zieerknvmE22ttXS2IZWNqQDn55SyySjwQxjClxnHosXdm5BQT1a
m0JTS6wT2+CyOowCzQEE3UxjAUxowhaEIR06Ydshm6hR8k6/lOp5OlycxgQguj8E5QJnO6Qp4YhQ
TO4FMAj3QK9urvGIedFRtD5DeKOogGkkxAQ5hrSZyqEAr7cijXqpSqXyqXUsOrorpSIwzpuwawiK
R93GW6uX3u7TLnWoB9jR2CKMQ+DoC+shyX3QuWtonr77s4DSkKynyrfLmDiUDrJTJ/SVbkQ6BnqF
T+EzYjK/vTxgOUITlufYXRTdWiVdM/jCAGx4dZ099Acjhwjz2VjGqqFsaxVufyZqjCziGY1FTUou
KtHFBju2bO0cSYEzSsc3Jwm6fwwNiMNHyW5BhkTPG5EyOokmxGZQMVvy/Csc81FxKQJZKFLdwoJr
QqwwSEGTJCVBnuNjhwmPxtRjMzibY4dl3zw+DARffl4DQSR8nTjEZUuVDfKAqu5UYqErKKl4V1qI
1oUTsZ5rS4/p6qW8DWuyrU7f8K8dohjmn2Gy60vajLcjkymcS5JouqzlxWlDSd/ToTgxQBstaFD5
YIbuoVv8aXt386GoY1dKEnas8CCylcJZqFsT1r0nTo5ASR+LUoJutYrIZb9luzu/PRJyjvQFfpca
DsLZcgOQm6Et9AjF2+h9EaBTFCyJDlHoRG37tu5612oHB6R2hdMay8xFcKCrINslUjnbpQdP/tgA
BjUXgsyGs4YPo7Dhdp5mAysd3hbvuiofnnEYweT3Ntk2vMITbMdyKWHqV5HDyxwyStiCQNcF6qTH
dqSSFiIVOsgjI2hfYgMGh46fjmmjbbtS0qFv8gRdiChmZ29bqZnJ6VrJWIiwWIQenHuhmh10T+Mt
OBkJ9R6HjQ6IfBjJSRX5yi5SQws6fEWmDXX/l8exQF+XVaJ7GJwAfHBT2cwq7bCiNQ1qVSs2Wmf0
D+y8AzL27JmYrdNqVN0YFoNlee+28PgpclDV+WArZJ9LsZHzROVGNVAqC8HJ1mfyUylbe7/FyPfs
JTKFUYwUFkdLONoD/enzYslwWDNRM+qHaXWz6Mfd/D2G0cYZp6TPmVPgyMMAM4lx0gFd+goDee06
h5qM8Ug8m3cUyCHDWJYTxlzkFk+uASsNRUxfunWHx+EB1Vk0t3kROChOpd06YmoiXdzEp75KNauU
PFgahr+65BEdKSN1nFgOA6iJM//Dn5e6pyqpDPBSaSoXz9pvObIp8275MwPSNmWB+3cVkU19DNgB
9nzQZVDKjiPP2yBbvKwvoaxRrnPKmnx3nlNdnFPthOoCvgKIRUtamq4IjNyYlkXahBioYoQ9ngAZ
J/vYJiM/MUgkyTdwfEX3xSUFg8rezJwvJvA7sngZE2NIKMTa8DBPJ/V8IaS4GOVfR/S8PbkLphLV
0bRKYMOZY+lbIlr6I/zyNcvwxT20aceU1Od6BzaSqFXWsKM2nhVkBihHryNeL0X0moKQGMl1GUk9
IpKPKTHlhTu+ejPOGlw/I4XXhU3hjzF3YOS0tFViKUG12XK1yZtMl4J+djAmf1E6RZDyN0N857V5
Ihpem0pmQKkd9oKuf8lAeBq3m2KSKxNqcRJGNh9wFJ5wseV6zGdqY3AC+XsIvQk7HyRRTI/WKiuD
4JNMk76KHDcgj6pAriGowcyyc6XGsIUjUd3Pd3JSXInB7omkbUu+U5PEsyqslSHA9K2HkMNPp0//
V4Ti7oZqb2jXe8bCWiKSyqyRhSI66jSCRXZJ8jwomZOW8UbR2AQUQI2z4vLHWCnRCpzYz/CtcVlp
wma2ZdhBt2KpqkC6SAdTMLdtsUdHCemf+L8dNGq8f3x9aM7jS9eLf0b/LstBIQIIAnQL6LzITMiy
D+ekDBg38dmIpTW9uRnZMKYVO4Rqv8JuUKuxZkFR4Vd1sWkt8rBCd3tJpgx/JQKKm8Hjl7K6KQT6
njR1dacJQCJ6/UCkirhoNp6CGDZ7JSTViikJWyvtTuNbv1Y1JKmg/qRGSJ++/w41dcAKdPlLU1bC
0Zhz2ZLpc0AWs6QptB3yQCWZSUsvinxpBUC+FGSXlg0M4HJLedmlK1nl1EECOcKxnG02UJ5QFcz5
6h8ulX7AAn63clYfxH7FFGLIypUdZkRm/lqiIE3YINul4ggLqbkuH8BP06OvKS600T0lRwlFCL0N
QV3OP/pqPbKXvKJZm37ViCs2zXIWXNteSZT7E3QCbeSU+rMCcdeqwtAyGiEbRXxuXIbeKDZRvHIY
IWgDftggFfpMMpM4E4gMrbkTLopYafxWDtMlnX/RcIr67J6PdxcTZjyZMJ3FhsU0rVzmEqP2HSIJ
be8nWnJih0it+3hZB4kWKMyoou3c6eFYGZiBzwlclV7W1zQNDfUKNZQ5u/f3ionvenXzZ0BD/zU2
lfTL1JHhN3ZVjP6LpzOh6TlN2psmIQpeZn2pIy89yYSUH7CckxD9VB/lQhHlCuIZpZc+ie7nUjZ7
OD2JCpRuibeCiwQ//pe/UgQIY4slx2z/Suz3Aihz6D7hiQOQ/CtDmqVNpmJCKsSpHLyv++4kWqLM
qii99OYaHb1XZtTNCw/KS8JvWrbSyNbAXb8mDbZ2eNiRrQw18Sodk9M0u8V0RNFpm4qSj2yeBk+v
1zG+ekWrG1rfWGZ5o46X3rg13m+OpvHRK6QXfYWi/Sd1q6T3Jm9A42RovXHYKbEAz9BbwC9KoDQJ
NLgTCK8uCPRE2ASvp1Ci5K/vZUrCzlJVcESbnxOPvZ2TAVe29/czyrILNDwVYp6v6z1ENxQwI0n/
moLajWODvwlBbFgNxw0WZcgmVbDjiuK2CmFm/NZ6TxT7kF/XqYu1wi84Bd583wZPYnEIeYbgmCse
BrUq+oGTIywMa8KWoYftyHYiswWm/ccZglBpJjzYY82ai2HlH1n+jRie1vSgQ7pKpSkK/iznX5ST
fUm0VCHuFT5JgqOYoiPn1WeX4oHPWqS+WsmzFcusw1/SJZzuxjnlUCyzUMjYvaPGsYTC16x67cgc
Hn99Dd7h60V1f0G4+RMK+Wvb/ev2LaACuAhJYfeQq9zJrRHuooRQ8Vx19nn4QHWTolxC702rASXp
sDaaH17KQiCFcoVytgfy6VDNI/Sls3Lzc24d4d7ir0gR5MP20CT3dLq+pKjA0mfhCx1C46P2592j
R+c3K0hRtbXZ3rN3q/W6+ozOFphcKQVcHbFhHLVUBUFbq0MK9q1BW8kQ0SDJYlHEMn8uHpv/L2jJ
fOhRj5GBqs4H8sNClbTz+OuDqm5vCTRTJ4KNqp9JioxuL61ZBnOmZzAfqM1GMei454CmdxDy5V/b
vVpwXpLiCEydOcFQNFsadvMSMDzM9MulvzxtsrX5DkNvdrGCpnuZhj2bUDwr5q7q80h5RNcaz0Wq
qIR8HN/NJm0FbB8PeczmjAVrvEkSR3rXhLlA7s3oEcifuPGM9o6WjUIEBrBy1Krgwcy+ndCVDs0C
tnJPIfgah+UM2LY2UkXuIWgYngfsgV6i+6Qf4bqJ59SB4jrBJ3KsxPcsOLBHQQwqPDSedUgeaWiD
2TlqiJK5GYyDDm0xefhHUq0ApdpWFtmwEv/U3cms2BxA09LfblSHi2iKBnGyGhY4M0OAwC12OC7A
8RenI9cnItFWelCXUHGSSWO1SVYZzB+5phztAuGEo+i+Be0Gle9Pnrn/t4MlJOkTLbxDFGZtdyFz
EkmRxXjhjXa/xgsGM72vOuGsDLM2re5V5L+IQFN8PZKXUk8DjmL+u64WLOFfenE0hSA7EPxYc/6o
8DhA2HW0CjZapPE60T7O3Iev+OYIbiwIuCTfi/MntMgSuEVaPqktPiZ92yLCHLwS2W72cxStcD1l
QMTOOMWlQ0esVnGOo9Ai0Wu5pl+LyguUnS2docXIlJzY13zvoFPXNKTIVAZWUmJS225SCXTzv4Ch
wrQr4JZsMVE17nplNCwpn5zoN4rNpjqLh6QW9X+xBciUtx9Fc/jZfZ4tGm6oRpKzHimANbU1h9kL
bCa64Hdl/x+cLklO5Gwu9EpPMNj+8cEQNVBSydlarL9THfE5vMLazuJsXNBHUjycry7Wq+iasMcf
Ye4dmogtMgEe8fixnC0hLC/0BAZ5tu6lmttEiYSiHpFHm4PVDE20Xo5ABBTSi+KO5LXGxdSY9kIF
d7WoU9SaNqo0KcmAyLjaSbNdOC4KUeXgjgrwjoS7SsUzCAwqRT1kwjnZZNTewCYltYejJ2zEnqtc
CPURFVGuEOczAyNl9SWWWdB9mVoW++pba+46vgf849voGQH234xc6R/K/jknciG4KTtDjjfaehoe
E8E6vetJIRXlFq/T53K309z18gxgDkh5UFzH05cr9Mwfn7ecUYaoW0fyNtdi4VxdlszymYyoGdtY
ogZ9lYKVx+hDaRtT/ZZEgD8EdlR9HlXbXdKmSOn9CSuEPy0qeY7QNFTJ9wvulzLblrRcDyNsMall
dJCmKeLglS/SawbANuIaOEw8/YnoA//0xHzOsakCOoBJ0GXjn18MDPDtUvJ8Jww302GP9kx8gq8b
udcGAps4ru6fkvNJrsD3ITBvjBrDAHvsQgkjwtgMI+DCBbv31wJ23pdR7EFfKK7MYyI5Y2AZgGPD
KQVEt+DSZyyLFvFDtGk2poNRPqGGYt1cWpJZ5kp0J1qVRByC8hnzpv+hKxQZT0wZWnV2ztDjtJ9W
FHKgEWsQYp5uS/yo1VqefbU63JxlZpha4JHXy5mGWMvM3pUA/9GHQ0iF2Y+1mf6tYfGUQVjHZEbN
uuwiFAp9V4ZvRkjUSPEFv2YyECfsGHLHPjhURbigesdza2XjYXU8kNggkW+x62Lr0GOJzP/f9M1e
CSY1OUg8R/NGJlyvhfH8Y2oyFsNS2AF0S0mpbMRRx8w/NswwrWoCd6UY39h/CoVhIK+gHV6Sp8wA
cjUNnKw8ePPEFeawJ0w1Al99H1dq6Um+5FzyyR5J/P1+0KCng3F9rJvU9Zqj8alOcRLrI3LOeWIY
PHvuDLyqnHMHOk9SFbYoVVuHtE69Qtb92vsh8Et6F/++lq6x94K9GRKTogXxDsZC8ycSdHeixZA3
+FIO8SpQqabA/rsyP8J/afQocPD5dLadjcAMWK1igBxnDLXtNlpXy/M0wtA+z6EB0jrzipO9ToG7
09VsCfO9gpf7NX/QCHnayK/N8Ip8C+nA/ddGXVHnQLqLmDyxV49NY6Ye2fng8aahNXB1VC/6152t
jqCFlRn/COgTH4d+QyYuM0J0Fz+8Wa463S5XqGHsbzqIo6/heLPERuEBc2JBBWe7hw0puvAxPFr8
t6fHkWxONkYADtUOZWe+3zQFBOhUDdYETCDJv6mml+qG7LbRZMIzFFgFxMoQWdT8qMrFg/J+Vt38
2qyeypuuJBxOGoUixYArbx7PWp+hDIjXiQUPrQZhBXVjKvvbj6yrF29qzX4gHSngbOXf29UkXbqv
EpCc0REkJCYe5Wd7lxJyZC+SItXkz+v4iJgNTUvNku863YKsOM0GpRE6KUCWG8xMLu9yLoo1mklD
PhHhd9m6sUaRG7r6ZaMDkeERWSwSOKZ5suBgUs0pXzavtEbqg9c6zIfBGmAM2yPOwEKaGLr8gC6e
9ZwD4nEzyWxLPY2rhOlNb4ZWS+jq1CP38AbfhMVU6FAKtoGie9JgLsCdXEDM1iaKuFCXm89LXfuY
adNAE0NsgtspgAIAKgS5PeMV9CnnjKzmrJAzYUa6k099Jzs7EAX8pKoF7L2s0eR2o2Jq61sQlVq7
wU0g9v8Aq/45PsLrWRl2pH/H6eXV2KqyckwmdNJu8+5ptDAt+3N1Oe6bt3KexlrSpeLQSHmbjkt5
TWBhkRJZuSGLgfCmFrlXrlPejQt3GbhbG09FE/MTpvdzFZY8G6p7irEze/59igZhreVA3kBc3GMw
M94V/NZG2erl6kOp8IOA12BqjZyEDyKM8n/BeSDBTKvKv5U+6DuKRC3IUbZ525LUrXWc5po30s25
Pq+aQ4l+Pg9XawaTgxx4/hlM0uWzvT7VpIMdHeuJ9qldbyaMeHjlG92LcpwPkUPpTJQnQnxCQxJ+
JnUOKysVbfNZeRGk7yLqYQJjh5zib/W2/zK7EsBo9gSGi0zJlWWNTnkODQJhL+RbCgfsrXv26Lea
fPGBU08Z0fTD8suZ8X4Qu1kKZ9W8BZOdmJOZQZMb9v645FH5cmi3Xk/pf5RCj4FJClIm1olAyPCh
+LB+PqTPZavgg+uhpdDh6NTeREk6edCU2FuCM5V3SjQPwU+jMcsvcKI3Dd0vMLLFDXI4IzTTkmlf
iUJCGuuuXaeBCxKM/EQUsCRmuIN5n46bV4l4JZUcBMhjtEI9TcjGX/nROO9K+y9CulQr6OUv9YIR
/3fpmbvbWTl0PkGcLefwCJuA6IQaVpYOr5yK1dOFiuXzeIJA9ZIvObDtiSDVYOERoI8QzvqMaEiQ
PWx+xKWnTryKnMBA0bkjRlGSNQ0V08TFE8iudlbxRyrPjkRDI+aAeWs8iQVZMY1tm0qUpm4VIttd
qAwpmqd8lSB8hglJLaS4/d4LrMnTMEQVWWlEHA3aMCunXrgrIWg5945xKqCFQYfWJd22OZlBPZmj
63kOWfvFnSV5w7g2x0R9JJdNSgCnLFBbDR6KWIbZiWDf0M6lAQnbFnXx/LYwI3VmCo0HIXz1BPUc
xK119aLtA0DqC03aohSmwNFaOF1BWqks08+wIcKxwkCPcGYQddZ6M41uOgaZnB8N6nDu2Zg5NBWK
3TYlYHAobK8WBE2lPlki6JHYTLKD9CZXiBXoUfqljCGOa0v4Xmu2TmeRgwQce0DirSHFZ2K8AF3d
L8+IxfQTvZmm3lWsl3ACzCJXy8nS5m0UCaaixpgOuRSQ0szFNv32+aetn1vOeB3gmVHngj55wbw3
QZua8XAIsRYFTKk2tm3mXj/K38LvgY7fVVZdNAA9Uiw0RLQpmE74wCfskNxNeqaZZcvnSi9CPaYx
yim7+3FgPCUwEQBXTP8Hl7ZWPIdYfVkdieDu/NNtme/SzYSpuP25882JFa7j+HNiNnyIijmqyOtW
m4o/RXFUsBPzCTj6pn4lua+7sff1Xg8kOmVvX88SwgtOURg8H0LP4h87YLxS7ytieHrjLNcrnQtd
cpdXT2ikxM4aNwsE4KFgCR0FizfA4bK+8rqMh3HFnLPgENvvzeAYolHGdJpjxK3DeziNAKoovOlG
Q2VGls2gvq1v2ZQqi5COJb3J4pzNFO5M3lAKE5rKIctRsSkkQkU2BtZIJVq5C29GidCB2KD+FyVI
O6C5MeSIhwSEZaLVwmotN383Y2ASOgzWq1YfHSQtF4FDedSPuN232gGYmpcSR0yaC38uP5laF2bt
gJNeSbGgYnNNmhw2uMcf997e75sKrGVCreMghJDKWIWlAsP8nNVW7CQ5ucDyyUGqXcMeOk+TvgUp
BP+7CrIr3GyCqOtFQvc7YP6WLk7KjOVGjoAyOsUUoLYFTn6L45HmYigy1BgdI0ZYS4DZue1F132y
/lkQI4qkYdR72j+eDCRgJ90BA2Py5SuY50XW4ceCvSgUNFNPzEeWpQPZsakS+YRL+gqQSEan52kq
49OMyZN9dsaRa8/kh9OSdeOUwKneQsE7L9nJQZnVphPlEmAiwQ884Hfk2yNbcykMNY2tv+SAHYQH
RIM/DsYVt6HBfcU1i778HgLyKDSQLYnGQCGKFzcQ9rP8kbGqi5rzKxP+0ZTCP9WrGrjb08txqPwW
JyFbuWYjxfBpyzgjiQS64GeHA1jhu/7VAEePFoADlM/F/p9rwN3cZ6j5EXZPyN4HmxQqv8ucGh61
HqWgju3f3nRaLorPilnzoFkkz8oTg3Jg+1CbWHRaeyRK2THJ4g1aZ7SsvARjbN6FSFykU4kGLAMM
TpaL+GxJIPKZAEjcDI3vAOAFDl7IzSqZShQTeRdCd1/hYJx0Nvy3Bi4KG1sUqc2Mq8NFQW6jPGMK
S8rYaHJIYSlJu8MxStlAokVyj3KP9wbTcJPtFFm282aPPM3jIA7y1YPbE0VQAa85gSHbxbN0C8Zh
FmFnXQWXdkWfwwrD9rdKPrwBaNIk7Bq4Mqy9O6Nj3gwMZ+s2CImKkw56mK3Rtx2BxM3LqGT8NGEt
gWHV3iBMlytGp8NOnw2omrntMTQT+S5qkUI8i3KHk5gAmV73/GFBWoJRk1ZI/pgvjZg4kRy9aXen
bM/Fi7Qt27B91rwsZCrNf51cGkdP4ugCp1hdZT+eosWxjl59jeSzclZ4dKQraA7CSurlfz3Vmh+0
swmnyfk+V8l0cdPItm1rMX+dQZLNE0EjF0th0iv/wQr3KyhamlEmII/57XKGjYJiGaWVdy3caU5S
XpmnKa7F1pFDFcjVwUP+A6YZqAs/r1ixTNgi+B77/Tp4PuyhDHYG9qynO7HZMKGxMEScrh35GhIt
bEIwR5qvTrZ428ZwdrlAJA8VUzoh4iQ0fUgvXA3v49pPJcNUjODokvp3BxVX89RAabW8QJbZPSq2
3eqaRBvGP5R+VqUTJFiRrql5l4s2f5240s1UxWiIRfv9cG+bNVVIKrJ8csbhRrdCLqKSL6wxUyIz
mNdarjkjOlZHPUI1TbqEKhA8l2l/U78iXE0Npsbb5bon+QsjSZN4BHQ+ge0aqKefYtnIQa8nge9+
ifGRgvM679El4LrQaRYGZjwo50Cya9GyjuOTki/anzPT6dDo6Ydn+OTHIt4sXJy2Ojpo26nldKrA
pnnbtN/YswGQ/V31lUZpciHu/A8EMpiQFYNnX26umdL1HyD3H2fN1yoWFgNel8sY7vMY3DF3ZR3W
FCYl37YAzgvp+zntGj7ls4q6GNaBM9UaUrfklqf7gMmGUBcMmMAoMJullzYWEWGf1A6xwOO3FhAN
Nlmxeeyjj4yC6mvxuunO00N8qrRt60s+To5yVenoz4umQZhTmwXvj+8fBrPdM4xp8c9kt07G+wVH
Roklztwd1v/YF+Bd+uvArUaeNc7PJKgT62Gi/kvCAmiPLudv78neoRZpOXLSPZl6mBrBekk0Q31F
/1gjzjSi0a09BcF9l1Shzzmf9RbavoEGHUzwCz4NlfHRQxDdAyRYig6+Wg0ITtx20NaXMJNXWlNm
FTIuvLdeSQxsRi0IbztyLPjGZ+wmlajCWnJ+VL8VTSwdXinnZMlLsoSLrScJK4fL11UkRsfnKRTB
fwKMJ+SERp8EJw992fj0dGDvApzM1AcWOC8dMSYtc4MQFu/YX5zUOTXVJPvjzVAuR1wdrhVlMTrx
LeO3TTR9vmG9oXTUwqJt+dcbERqvesl+7/MXuT19hQc53jKcc435ZPJLOoSKC67WtdGODDtxwhtv
gIvqePoDv8GhF1RhtSbqg4l6wFvAn5eGZj5cZf3i2H9JRWSmzWtq/GiwLM8DQEQvwXpawNxlVGR4
nTSs20X5NBqZLrm1MEydzsdYFT+ZIvrjTtx+VqvExvpJiXsTfqBIL4YrRYqIkZdFXqy1qCiAUpQ3
F1RF7qkZV1AzGZ5nCGqbVeltvwCsNAWWt7nWucLB99yFDFkG1GqWA0Vm5zrN+Mp5mmX3nNIebVNm
8a4ElVbwCvdH4qj9iE/U1s9Go6w05pZajykT+Z45BDeV5Vt5RyWRvyZEhbubIEvTpdG/6M8drSoR
nBWtb8iUx6CAfJMtPEAu/6L4pkIp4BEaxKnzOwGy2P18V9tDnjiG12TySfc4lxl0mBhR+pjVFpKK
u/PF2H7csFNhExq0x5r6TjKgdLrKVo52XQESRPoOh78DDoHWJUgfn5e+oW7vVAoit9tKmye+JbLQ
NcWOHRkZinjqH7e8dPv6U8n3L/YojUfN23GHXalhZzWEzHnUXdicZoQojdSy5skJBPugQ2QBp3W4
XfibT6NgvksF/msMZ6otMXSHL6+yj0AdpBtO1AsAfxhpU4G/oaEHuYXh3QiKKD28b3qjvNkth21N
CGwQYpHpClivVbfemEOWxpuZz99NLDdqr+0tIBhxB7+X3gTHWFzttdhbySOglgeH7wl8O3GWQliC
4YGQ2RrnwJ+T+15u1UducIwx5U8fH9AfNRKatOT+mxS9tRRH6PF+RbueY9iBdxXD4LM2P3PoEQvD
wzt+veRcCUK3QibH444rKnuqj4vxu27kdI6rrTVFDb2WqpbrWrZnu28wzKoy8nkklcXbLyESxS//
Z2Jf9UiPhN50m3LNgYCdu528HtK3smdiMRmr9MHx+6lw90TpiJp4uECZ4FL20gSrsxt3bvuohjPR
FyE3ITeYUu5VquX+Mmd4P20Itx/9kLP5kNyXmic9sZ9gwjub6TeOIt1OemApLql+Hjh461NCFSLZ
CQ9W/wH+2RQzf6olEk32oWrSM0gDTti8aV/mJCXurcbfSQV5Dmq864i7edLW+FPuYkBYgGSOZBiI
Vm53M3Pm8wOoXtE7AZCSA89DlCd+e8rQH000N2OQlCmLTSgg3rx/hxGUAqKZsf4sP+hShL2JfnNm
N7FPRaofV6rtkGquLx5qTGAo1LKsRNIwwiWLyEjdoqRHeG5QLqArywk6ltfhizhJt874tWRv4Bri
qK0JaTKfHMVAqEXbl5KVDCaRW1q7fnkjJ8zEqes0F29CKfQct1sTSDbx7eYdXja6r9oz+6lkOgcO
MZcxAu5IhlxCt01KYIsagN7oVcJlXOqXtvX3T+S94qXKCZhXgRL6Os7musUNcJXJwjiGSVNbXbiN
FCp3ZJrglaCckGbL3v2kYACxS4lJdgTJ1hcsYY5PVg6aXvOh4ijoWHtjV/SGkB/KqqYOETzkqZqt
NKehtmrj8j3GAduOstHlOc1ERv9IwydDgwoDC9FV+7sNoMoBP6B6DbowWvuI7Rnr2W4Bxkdsf3z/
7ZrgWe9ch6Bzz5gjWSWM6VfK2m2RHsfJxICVrz+13C2mARwMKilN9hCA60VSn49cUSxdaEgejx5s
O2kuyTzhaWqsCXW25EEa3/jrY5++AkjQaQkVm71tNkfIthp9cxOf69BKSpA/Qn1svw26l3AG6G9+
8YJBxFWXakk+YHTNftoA2Nt5Q6X6GrtsH60PQL37ITyGL3ncI/asTBeS9QMBJj72NteRUOWX5j//
SVTMMvwUH3y8t/NAFXsiprO1JrzEyAc4HBVOMZ3Jn0vuYUDxKwrUpIpSdiIqzSbri9yYzL6HGQjq
2E7NOLTPRopeYKt+ytWPtl90YcFKZ5zZoJ6MxT/sc9Y3xNY+BnZIWkRBkxIx17f4iXKtxQ8Zs1X3
PRTQn5HoGQi03l9qDHjr6qQkcKKDClYod3oPgiJemBbsw7dRDmVfxmU96Fc5Ibk+v8LtSb7wWoNm
LJ5m04Pf9a17I44FYRYhuBFBL7xdvlGm76sSNDCRMd3R/FD78JNWMpNFyWvO1WWUeI+7sFj0+89K
VKQDYiRCgV1+a2Q05PeVGnJQIb/hCp7gNKTB0jKWJmjQLa3Q8E9NrUl5AJUM3TlpbEv4zJuCelNC
sn6ff1JXL2eDxB2aEWi4TSFZ6UnXLDGZVknx0bJFrnpnlpOk/CmrmB7/1/ZIveKYmU35d2epcdsH
XsDukvSAOjnTFDb0oJ77whfTM23QviPPgsXVCKd3qtzy7j7U3+pUm6qmUL4lX47nDULXLJfFb+xF
zP8nM+TMjIUjh9sO7qbC/VwLyn0VBRd68s+woswM4QYwONOHldaQz5iCaKHiHx40QxE4vvSVd7qJ
CCi0TcFxY/1MSi9eotO2jWOz2z7BFIP4eLUuSJh2ynKmK8UnKh+P3e9y/jZap7m0Q2CMxQ11XEtA
NXh4pmdq4j0rvBlWmeQ3q3JB44PZziLWfcdfWXm3uXb+5VVcxHYQkuF15bti80YOuDnCLhA7GEJb
+g613r7DOZ/o9HUYmBP4utFv28aof249y6V1m7+zskvf3HuR8mQDmLxNWzNWm1Ca0lsnXkqSbgqD
M54xAQh2IFv0upf5NdVuZ7iUsXm2qoLtA+SBfCIM3vhvsGpq4qo+dKrbxhy3NjQkh85OtyBqPubv
3YVBKLLkM/bvpUFL4QcYwi5pzGIQehXoyqT209N6ppIFhqAKnCei1xqx1fqaJvLJN3Fgyxwjyk07
ZXv9RKGbeF1T1HZfVqkO6YvbF4Q+Svl3bN7wrSQxhF5nFzpwZ4gMLCL9szxgvgqUxHsNAQT65qPP
PGp4vAjXuCGCTUIOO85n2xE7mrjtIhzq2MBnPm+N41Nj5LkMWpYRsMx5v+QVm1KUjIKsaLQXbPsT
cVCWl6onuhGN+u/VJbqa4ArNQQwwwcvxtJhpA5UumMFkHBeVxXeJoXKVsxq9WDlTZi7ysg5rBKvQ
m9qmkFk26woJp3dBpIo81R6oD0zzDZjyed6BSKxWrK+KT+AxCwPcOgFj+MqIFR5Y7PgYD2hr+IL/
UBsne0pm3QqpCgNzSJGEQbXL41Q2tx27Jgf2mQKfQKFDd0+6hU1ljp8vztdMAnSbYmwEW3TQ23jK
tM6ly2t0IHBZpgX2xYQzyyZ8AKz6C3D1q0P/6tPJ/rs0valKShfMHSYsG5b1rs49k3pyEwP3PPNQ
mxxvU3cVIkZcAm6LHoMI8V8TXxoopHEgg+6XI4MoqZdQ7IlE+0NgVJxN5UI7vch/ItJwiG0Kv7Yb
iW1TLsFDnbiwLv1S0EqHT/c8BNHhh/u0U3zftchDI4lmr4pR0OqdgZr9L5fSEFQnNu3lyg0NTMSy
3kwLU+r+rtPPn/Kr01r1nUzjk8mC0RmDhJc8vc+mQmrnTKEoJqEWQ9Tv2IfMY7B8yABHN21+8Pjc
1swaO5FJzc3ml5mDmlQnKP0ereYxUK0M2mHwsGxGY6Ovidphnzs4hJToZdg1ch2gVBvkM0V/pK8n
p9s5E0Qa9apojWxSuh3MJ+aZsB1Hlv+WZOn0SlYtsUYPQJd4fcmbw1wE1MnoXHQhfH06NZY+SGwm
pFTE5OnXQGS2KTdgx8TzGpoXsQhEBmYJQUmFqHiFME1NPa7skI3AiTapWoRb35CrH6RI9ZT1R+CY
eDJA8ICy5E27iPFo86pVaQAk6Kouhb0VPx8v6GdPUXZEHHlSnjMFe9gtmdjW0pefwo/Q3HX3KVq7
JKI5zwSl7eWvyiGHiIwA/VlhU+uyU11jxwfNDGpJqAQz8jZdSr2u3yWyu0flA9U03fCuu//2WHxx
yihza15EUpenbgtaIeyZgtgG+TLTLwYAuFTUN0EZtKhvfEWHxUi1qpGZ+ktYpb3fNTGIOYOXgO/K
HgJX0Jd5/5L9ZPC0f4x+swFu6TU5ZJGguhrj8K5lNMBVkqMLXzur7fTeLwpTFHGmOR8wob9e9zn7
LiP4miRhy7EZIMFHwXCSCaDuwZWzVLZeX9PfarYxa/XICJaS4e7jAtg9V1s7WIa6+Cj5JzgLBIPO
ab8oORNM1tBBNw+Izzr/dR/r+Yf2Sx6VtquXU+TifHdui0+Rdxm7RyyDi0x8AYJR5ymLSUeeDz14
aynbGj3VbJKkFCRRf2eH6Stb2vPsFaMlzTi/Az09ge68gyhbPNHPEf8eo3AkacxxxysJAWH+EosL
cqs6UEyxNWhGPSOmn4AnbqhISuwzC43EIVfHQvx7HHtOoaww6h96aPg/ppwFoV1YWBQ/CI7B+tIb
Fa6T04SfTq2n99G08WeskOYK/B58cdFD/WpHW5JJp2NQnaTRRXF2ta0pyIoicPBuHng/zv9tQ2CW
A4T/KFZmwRHPRfwy8p7Bg2VFvoeHQsSKFcEQUHqVm6qdXIWjVgxF3MrO0TisuKUFXb8iFzIbb9p/
DA6wJ8O+LIaNglFaiuI8EP7dg8oMqsUTWmDu1Mz4V4flCmxHGCCazWxG9vPQ1Gu5DCccOEfaoe25
v0ri+GSwZcwWtBDSzz3Uq5ego1cN2B9+xff21/xWCeyvC5JHvUtrgQmphGSXDbfPAeswP/QBV4yw
zV9LJqJ9FZynA1KaD7ZrBLEnis4CpK0/8/SpMU9E+rUcuGpts6lh7bcLv6fIYEAAoRJlVDzP+uXR
NBverHOyvo8aXLqJCkrwA/VUYbJ/02tiW85SO2elYnM+F4Wd69t2M+ekZAV0yMO/OqkW0zkBhBQC
1/Q7j1jF+AOMRt638Fowl4Ylj/IXgyfP9UqLGSH9qNa1VRU9Z2heNVZ22AGw9EyaEgJmwcWzCGnq
ju2CKpH5p5J8eB0aJY4QqlCd4EtQ1E+nC2SJha1bTdPppvSGoJOF3TPMZNNsfI77QGMONeg8b49O
DhxLm5ol8LG/Jb0zVbmSU3fyMRvmj2e3pl5grfYFN708g1LwONY/RctqF1JsB7LH9TjtDU2fjpG3
VsIExmahY2inljcMumsLHzLtHFq/dxE1h4sHHSSAjAUTBl3yaWXXOJovHP4kLyH4IBF0zrIsoEnn
ecQD3DHTJiHtXGNkHB5zl7KX0KV+oVS6cXTS7r2lclOld1kJnJgJBERN+6kwZ8C0CSfo4OrYR1pq
NbJUdDGECmm5Sbso4OXq4VV5xaZ5DtZKxYQpK1WjVleGgLSJK6D53sEUhJuBUvNoLJJvywPgcM7E
p8AyO11hmAtOQkjP7GJffTtGVgJk/f2mjZGhxtzWA2GdYWPktk38SJ+bEGrMMgu9SB3+00LxWEQJ
FCWOFS60OCYl1q47qTKeWyLt4OFGuPv58zf6crsltO7pefjbdyvQDvJoYl1XPybZAmcXtdb0L5MT
7dzcDlCyRII2u9oR9HOOXe0Tl4jLkyfxF32ZLNGC+bfA5WO+JptmSugFxvw6ENSqZfR4q8AZaXpc
E+xGkMxenTlI3pnT1cChLQY99/cKzBZY0zhMtAZEneZU4KkY0flpl3UDs3Gc1vtLJLwC8GLlBF3m
pq8EnP3HlF6E4oHsAJPSa8IvJrV1FfxRLPLcI01jEV/O3SugcCfEJp96HcY4gMGsomNWbH96/U/P
aagOMEwDUlS9kakFiW/86sALttos+1MvsVZ+Ua9Zg95yj+6N+oeGt7dyLW8+NOZKWrJSdGolcVOD
Wx9Swz7vtzKzObE+m5dt6rh1NFhgbWW/72SvcsqC2PjAGNgGQ2jtiF521l4WFSrD/lMwh9ccMw5D
3t+53O0I0bn54DLbtNNfQDtqUtnqUnBoEixxnWPbmtXJ2C22Uu13WVQmLsxPIfB7bpnXUFT3n6Xq
Sb7WCukhw/KioD/EflQvob1LOkXNPhDJ9VLgsFpD/bOYQpr+ncWME8Krar4PzF7dkp679Edl3KD2
FgxFkA72ruTkCFAgsU676hRCYx6PGgaRPYsjcZwA6iBgFlin19bwgS5n36l+Tep+9JYXdG5Go2tc
Lp1+PWcVCPopskHti1a5ewxJ3wd8psDg0wNHf1c9NDKKuuxYpj2FNI8ZOtOdDgHhlvp3i+CcxPZi
85tyQ9G2mrYB8bQ8r5OKHZVForioKhjL6PPntrXHRSQ6cgi95OwfNNkJKf13Dnf4lMmEGhFG2dXe
XJQdaaGJ4NbMyD6JyEwoVgRnlkwlqg7m9vA0VD8lyjJlYuS2TNkdHBee/XpsYFO+6rbyDk7RpWkd
U/HKlg9yQSmE0xFR9CRwNrUrdg5xqvCZftwTB5XkhfYoZPbU2uRnl2NDOHjWIlsEw+MQZCsi2TaV
uplM71XW6bQ/a1nlw8kR+ac36+9Zw3CFjxVPNgeXYEONilbIETPvGYAZHQKvrhiFr5hRu/LnVnva
WGEqeApec5jD8oTZuVnoOlfvnOHLNXwDZktE7w5cv1XVOlWWchadxWzQORD4o9CReDs3Qwgg0XxR
cQyq2/LIfm3RyH9Wa4S/cu99aLM9sQf4i64OTR+RKJgZW8e6DSMbeav1lcgVdOC/aFSmb1iF+sZ+
6FygSEqTMHTTAHRilm9bNaz6E/12KJB1cf/02Y0F8YF5Hk/LdHdfAFqAa5BT66vaw8nwRieLwvHR
hNa4b7gX38l/vYFsgGyNby+qHRFuYI0NSRPEH3nVhWhIAYiAuKsd1Oqw9St+0KXtFw7ST0MYHd9P
ua6XDAGrIe84FixdlOlDpg+qxacF9O3iezH0yHLPfm4TKZY11ag4rBC+UFZolOtOkU2F/7mdASyd
kv8n/+XuOg/eLlGIQuG2d+FcqBQNndPy71CT22D1peP5PJzCL8czIxJOm7tYJ52p5yvi/4mRJEzc
iQZ99BWoWmQ5piODSC9tr/sNoeIUzst79DKucNF58JPslR7SmIY6KkwFvbHfJ39viMhtlp5MKjMv
GAy55Q1xbsR0qFQModE390iXNwaefs9mjPp06BArNLDsYkq5NCWK/F9rKDviq8eU0zWwOCWrYSoT
nVU6PmknMhS9lLO0G/1N0othYZ5TrBp4MjN577X2re40taUehQeKbHlcfkOxC8AArDi+fOnvz/5q
WdNKkgQAR9GTmLF0ldZGj1SS3vFWmKtLpWLXfM3eiz25xLtbS/uzuwMbqzM03kPuxE3ITYWLpmhG
JmqAI+9byseVR81PRMRgJX599U72IoiEPRjdjzJc/W4KPPqrM3uFLBOsc3K0l8uVSAKrl6rgDKJ3
/2bPUY/X4S5kO8KK+8mu1OGYDO6l2O//hllt98qotmFVEW/t8bl0oYf6cOhYRM5cwuhRUtWfawYG
WxxmqhHQZJvkAx1uiBT5POZlJsRDxnwyyT4wuo+AbTSBfw/wfVc6Si614WKr5bKW+xm51XD0thP4
IsmRe2MqLstSOX5dezmvCAbp/8q/YAv7yKz5Ods+d4RmDVG10D/71k2IcmTurXYJh1K5rVb4YSHX
WhiCyb+PNyBuEqykrR0kQ5ckEdRjuQ97EUnu/JLzn/YDgxkglNRhrMkzpwM1nBpGTz3H/6RtVi93
5fiLsHB7qTOyDujvZmWfgr2NGYko6bxB0ioPvBkgQCCgLOhoumb4hPnqF4nqHhJV5CiKxg90m8re
ZZcemE1gsMUo2kES9NdL7KHZjfzVu77E0bsNfiZzPaPH0jcuI6Bmx27PoxZQZLCtw0CyiGkQc9C9
CVMxJdQEW68dpLDAagm3ZnUfsjxEZw3NmqqQz6hlCh9CvG1JDuCeNZ/onXZdcWCWsd1wlnFu/1HA
mOZFjbxOBjfLuDr1cUZhitZZHF9PBaCFVNL9f9rMETZBnvtgnnbuG0GTKnqhvUXc2Ji+8L+YC4qg
CrT5kltCE6FiVdMWEJJghdbAm7EjUXKpFkOBpSTx3BbttV1kcMfgfCnm8kLvmj/Nx0+5UmM9zynv
FwTvsi90zjFZBKgaLcyJ34QI/+qahnV1CFXj9yiV45lSl30D/RNZT52UsVG0vBsHwu5ULoqraxqn
s3VQ/BpKR+QUQ1FdvmhTOyYq72QqdaAkaWLSP3QVSgoNufT0u+e3nptvj8A7B0lfAniHFWBw4tal
CYrcRd3rnnqDoC2aoNbjvplQe8NBwLfyjLp3pmNJERXsEuO2mc7Vfi4KRi3RuB2Z72y4hNDYNbUu
Wio7/ABIpdvjuV6svsxTugVZi1XAW/BwZfn7VGD7tOhQYGQ9d7+SAAuPLeJw+Xc+B34ADI2kEN4f
f/jaT6d5NwkIZk2smxYKliJ5eRDhwB9hdQL9k40aAhY9chaBtxEnRXt5FWRN4oIf2TcMN2o5xoNz
f1etgbVxiv9FjpS1+Dymz/5oPWPc0peqwnissnVg2Kl52pUhgPzA5W/65mrmPSf1eCtTWe0kGVff
Fdr5W278jiEY/ytXF/KY5P8wpZaGGTts9SjYRTqNh0eD006Gu9LXGHcy+J0w0npj0k/3ZopDNBfM
mAzj0pU4LfVbjnsY2flx6JBVtQlDNQqlbWd5TL2RZ3pj+It9YXz8YOICxRPiH2L648abQLH+WxSI
dry5IhLKxAy5LWfwBkW2PtMKZPT0mTqkjXctVk6Cbmf/fQxaovCj3DbU8nZxhv+HDl+bTX1tRyaX
pfoexm0U+JakXJgR73Rx25UxOUfEwBEtfRO+pd4uaEAXGFCaftgUXSnFXXx/A5zkOVCU+pBcLZ4U
loT1OH4k9agZmsQgfsUeG+uZdf3MW7Xw99ZuYialnCQeQJYPCpSO3akZHdhQ2mQ+Ddd+9euQDInX
YZRm8I00D3uJAzpdnY5T1XcrDD4OVxYdEJobLxTa1xFCbu5QGRlAwXtsviJuT8Lz9KL73VD77yco
9QT2A1isozz1Y0Ad97qGUZTvirAJL1oib1N9ySU7l5W8nzs5OWaIKDurnfWfLJDw4imdn+/Kv7eU
237WJtgMAzeq5pOVz26P02DmUlGSAHPGgbIlH5Q4s40qpbPqyjoVpoIziAiuinhBACqn6ejNRFLc
wNo0O2DkXw3ecwhnB+Dw6fvJ26VPI0tXrty26vvtL6EERpGjRhBLYF7wY+A1dHLXRysU/3YyNqRw
hgiWf5QTGBddPfmKqIXg/2ZVIozt+6aLnyGme0Hb+nyp2RXoy1Wp5mWBgWK1nxsi/lmLzQEKizxe
IASnSSOA6MT0MLcwkyjyr+/gz3MionIQj/dfZicL3hR5NiQKgEc+nbEMeVUJ0vtSqFUGxUL6AE2D
M159FswRbd7Uyv/avXrk3iRZMkYKzC7TBnY8c3MIQ2Eq2jQlb+ybvxLiHan10GppkTTWrJ2R73Jl
wJtATVoUqx7RQrYAiLXQmfFZqATFhX6/KjqdLaOR8NevfvMBMD5/B1XmjcG3nStXLseEsKNF3KWZ
rqw9k2u/ZumFre/yf0VnJCySIiS7pUK6U5XZzeIF4Hu8vxlkoN/rCqCFdMgIMrsWCozlzYsg/8Zu
TtpZOEhd2Wr2zJw7bPNSR68qTUZECdouwUQrl9LL1rlYeO9LrJh6wvM1M97K3bgZ3Qx69Pf9I4Iq
w4mnMS1/O/6fx8rY4VR98MyD9hITq63Xybn0btDhojBBA0uQryuvOc/urjBII9HKYhk+MMmZZavC
16p4rpQ0ey4EdgH6gtDWE/sjtUGUW679N4JQQe/vMosYvwOfOpwFPRjFyD/rjBpVOpdIjItL8wtj
fVmdcdigw6QnyOl2dD1VhoCo2wGe8Nmj/2Xg2phNuX8wDYpoTkJ22qeMGFVWyNTZT9pNIj3KuIXq
jutTfbH2qrYxM9aKcotTz1dWR5HIwMdZTTbR6vriukd6hHCW89R1HbmB96kaqRNZhiSo+FwRnVCv
hocLNndKpzEnwWCviVXAYiIfEglVUyYRB7gLvAf/OFlsDmHqHQfoMtPPMlZVjnPGwGoHZum1PIwv
zwE1q+9QcmG9JEpH/cfJ9yNGNKiuuPtD85veEFmTzrzkdegssyHDRorAJ1zMR88DKg6AUJkaj4ha
j2INd5KMWn3/PWNHrB2ZLrKBxeGZrPG/H9Vddt70XHeQ2iwT3ci+7GzuZlF2V+h80i6GPEacmrGw
Nkf3HQ+9NIXYeHMp5StgldbYNGNjvpGRsceTN6jEt35x/5DnPDWbhdFAv/CZN2KwXnpWiRPYg7/G
CDJY9MkaQ7G/gAi7pGGRRvrGeMBHlCeZPxCifPL0J8iv17tRUY2IeA4ZRKHSLSKNd04ztX/pTjiM
aQjabYRHMbt4JD+zAgzmgjUbNVeqMjt4lDFiaX+qCAd01dMAYK+/0tDcYVHK9k9TEoeu4uMBR2/t
GfwAU+nqZmu7npGlYbPgdoHqpqf9vCZ6ThYuvKUtxUugMx8wwxG1xEJ3yI7ASIPffrF008PUPGIJ
OoYA1PTe/s5acXxYqASKMF3iTQmihKFE7huOwpUJ+Q/L5A2495zAxaJyq1473KRnHNEdo4g4+PUY
KdsrM4EQ4OaRR9/UgPrLtzuU/rr9JpJNnxSw1RyVUSnDXMvsvimBkAOA55gl0bLbjFUBCL8remHi
gWd/GNyR4+WK0dZITRMu8quamQMFSJa2agM0R/x9Um4JVgO7vpgDFpQilgg92bSvVYIBKesa+GHX
r/VETQ8q0tG8btCge0GV1pUAdejlg/tfiQID9kw1jsaXimNOuRD7ujtFsthOwxJr3S6a+plB1O83
iP+rW7HyEmU2VD14Tzmr5o9zSGc8FHQtWvzpUlZ5vLm2rcoJDsodWhMoY5V/cWjA+hGfm9tTvLii
7J3Ew/5p0TBnhSidjJTVDAQt/VSSCyZopFImCS6PI9dPQGwnguHQdGiVGIx5ilm4d/hCUf8MIE1y
VXVmqPqDm50XJ/AFPfZMrm/WYQvV7Z5M04mG1UW2VU+2pH05R2Y/3aIDHavDctmRsJt0IybwtEnk
VMXQxaFLEz83Qu4Tx7XL3BKu48+bKQaL+T0SLBqOIgST5o2epy1ryOdqCGagkI4b6AUcY6yMOjHv
41lqucOeZGcF9oVJsfYLxVptl9XIwoFursAVvgsT2gI7r7OTIWOSOcn1Gr8QeguCyQqCJ8eAfEx1
5RXPMrB9qmLBdv184fKFFVWADsybsghso9RJ7J8XQsizGSWL/3G2B5xS8zdaMwW+TUZpYup280K+
OwMW08C70A+XkiVKu9T2pHeq4leiX1CkK9zuR485ivztn99idxaDeahWBYyrnN9SOqV7jXQce+s+
Sul4psyOH/ZMmAMjNqGpzhiIhgIVW2Eoi6ZRj54KperXhqqwF7tUw0KYVwknOsEokC/wCt/wIT8p
bQsRGSjwxI4rdSaHj7/5Q5hj+JmgLcOdfYBuExojFIi5958nZDB95C3+CKWeOry8xlhpcrYKpA4g
5O6jxk2JkHu25h8QClhbIBiav8wkKMXpgU3VONuLr6FDyXI5z3C5IQHilHHQBU4tPRzr05IYKMhk
0aQfu368Ebl+JZ69YlJk0OutLnXyV9UuN9GPIYdRwp2zpiU5/h3McKuy/LDXo+OGytQGxonD5u7T
cWdiEcJZxnsxkn5F91uX7MukBVxZVMTaDO/vzjCmC2GPaEjvz/pdkHDn6qCSHcpGM8p7KEKUvH1A
BjF8nsJkWtfpUM8JYYHQD4haeOpHzZs1vV8tOW4ib1EvEFF7gJpsFQSZ4e8rlt1/wquoNWGfxhNY
Mc+MPUeyzH2J7a+qvIyQ6aFoqLodZX1cVvwpclXxHlENQ1QA5FLqAMbmr2yc6F6zeYAedhnr1r4n
5kX2N60mGQ0pdO8BkfIgft6TqzJFSnW7L4MiHB859jgXJ0uLYHHhstlGSS95j1PUJDNb2hD7sL5B
FuFZeJdmtUFC0DDySaQVAJbAxXabwc+lqJ1EdQDiDrnWWljr7sSdz2PeVbMKA4w0uA/SCVMmXd3w
M6HV4dhecYmoFxarriTEcptP4FX6ryn8S+EfVEcxCeouO8n3YA6czEfdPo3N2irv/YfpAw+eCdi0
mFdSKVL16wTAF/Lth55yFyuJlTEe3Sr0WYngx+qnsPE/wcwMyyluv9GYOGGW6Mqg9JBlJ+WECCDn
NOFFaAugGJJ3BsBbILCqgatkyYXsq8FBhgue16LnHzIhwL7VIGp0eshPgYNIwuKNYvfVWNQVapT9
fpzDKm3WOt/m1OOmoSvDERNal5DXzi9dgDQPlQ+36l28ulPhxJo5ij0TRXLO/KQeLzKiRp5RRi8n
tv+ZJvDCXQBHW4MdM2jYiDHe9GVh3eYD4VFjnPf/23sEOs0dq2NausmwmbDuEyPCKpoxuE5YHOky
buaso0GoRXJgKeuukguqFh4zkJzWb3h6X2OZuOXlkM9SkPImX0V3v3qxTUozLN6fSolDNFiN2ln4
OOBwFBrEe8zHqVciTG+0bdsmw26eow9AsQ9LMF8uLbd8KonL7vekqylsYtDrayqhfX4xp+YSpDgt
4rE5elBhk//PJBEG+AsujvIEFQDL2L8345ZqUOlRC4+ja9Q9Mt08d1OFIBYiku5b7h9J1YwWaAfZ
QS54xXkj+VOzc0MnzjZN950iiB8UcV33QsvkPp5SL4dXwaWs1iCJAHR/hyeNZwTOGwG2sWPx/Z0X
NtnhgVEiXLV7r88+rWE3zOu02L13QnrK4/Ph7X6mG684/LtzSXT8fUKBn0bsNGRgPoxWUS7844Vn
q3o3LeX9gdRn6CL+dCdmY6Cs5nIXsDcn2ui1iSakzQl0T33B/XktpKVGxGRnuzbGGqhWsxjDuuEm
Scxn69AXNOgUQiT0s8uXp9k1YCb63VMNFnJy0Fk7Gb43KMohqF36VGCYT/RFnXUhSRzzlELE7cPC
RP/dkZfJSHwOF5Dd2/K5l9EZx5v/YZf3cYSkmk6IGGLpzM2B5m+cjeZ5tjK4BKPLdbH9CMQ0SKdg
hKSC0McYq1Z7lgncE1kXHbscHWYv7mhIGexMTnoNX0vdg1fJ1KfdQOB8Ks7vjpd5sgO5fveqIF6L
32ReNuiIvYRrYNs7sCKIflbUi579PCcFYTHT6XlOin4cW63yneffXAA/w3gDmxhnjuN1gA9dxYXx
BrRDkuG9/BxgJW8DmLi98kA2gm+mqe7mN1I8HpLdO747QPLiIlPIfU/o/VBk8exf5Kfcg95UG0SJ
dJcCFeYhTjIh7gFVDQlACOUrEl5EqvQCJIyMxzaHSCVdGvoNtCrVIyWxCrc0I94pA8AFDANNQTKM
n9/yCJfu4u2QALuYNARsd5Hm3aCqDUREhdHz/csDIZr/WhyXRx2YHt+b8bO27WF2Mp/xe5b1xxAo
jPRF5HZ9BwqIO+nI+ypmU+l8xiwgLhSTBEMgVyZbR7BmdtxhcccBNL/bRj5nvngMdjGPHCJoHNuQ
2bvvicLOCAPzQSJ/HllqQMrcvxDq8Pq7Ortvk/CMPcumolyM9tkDnMaCWL4hvLwPkABfBTwuxAIi
ZiABpncI1FyZhprEDTJ6LEE/7MLjgbZOP6iyExPvfbcRYrQf4Rfd/dwWW99qE02wXBHn9v4kFhuz
xK2OGVJniw6Umq3D37vRtDVWPw5mY0tp+dZd2D7m9PKfKYyu+5p8cGWhRv6jTcgV4bWdt3y0urq4
PvepdzMNz+n6mMJ7EyxjZC6/CGibtMP9y9z2845sbehNrudivXvV6Mv3FomcvVWUMZW9sDGa7aQC
79R03faafBappd09Y4u3SEjUqqpTth413GxWC9gGVU6bPwH0NSh6Qq036OFSvx80dya/jNMfRxWd
qUYEkSvgg/ATLSyLrXlyUaX7f+qKX90S7ltG64sV4OTdsD6sUMT2Bmg1IHCsPKc2HjyqtGJmx0JF
tVNMOyfnFSgOXDgv2+Ret/1IYnzdID8vuVQmNWHwxBZQ/83YVwYIq+2fDo1gqogddMlP5T3m6aaQ
ygBIE7PNzfwmqYqbnOoWbxldve+lL7zL9cTLXGOfHImCOub45NTjxqw9AKkOYtqF+ZWO9Qeh4Vh0
sJj7cw4sZEtK5QNh5eKaRLWrfTC+DhQgf8gfzdzI827UAzkTZ6cFcTn2y38aQQZS9EvqDl1osGJv
JXAGa+VZWy/9ueFILNUEhpKF2f4eEC5jm+SbtzWcZ4ZtJCO4MckLfQWs7wGJ/BTG2d4+cAcMEaKo
Mgv647NmuQ38s/sVY8fqQD3PMA+BPXe86pWYhVhZx+zjjCRpaRDMDeLEzLIM/OaT+CLkwom9Oa48
UG1UOBAqnjZij8ppef31gqd3IxvLQe/VPOt6+Aoop1JHCBqPyo55kQixWYjOfeoFUfNBeWMBxcf2
fkb/Ob0WbiveOU90t1kPlpNGwyMoRrTVjDSdlbE72PLNoRldqAAu912/5CLi7Yzz6yBMSumFIOKy
hL0XXeWB7M3D9W1Mz3qPj22tLxQZ6B2I6BcS+xGhJGkwoFq/yP0AtxW65DyekkKQ5hi2h16HvFLp
36xTqVjDa+YnWIMFZdP6XUT7kL6pauwzglH8W7wH5Jm1OKpFaF4ycZNJM+mpPwbOJ+X0KTj0LHw+
n2x8CeiiDhm4ynNFuSWQ08jvdMOWOzQYbndcmZJ9stUm4DaMqJ6R1Zl1P6jvC8Nq/wSbEQpHt5cb
p1c5xVaV0owr3Ln+ti9wtgRCj6IqLBrRBehtHcMjk6RtBy2Abq5SJVCO1QXGt9BPpELYTkh5QlCH
zYX9sgEWgc0bR5iM+7ETkoS051/Ywuyv5/mv/YyPCSDlzNfyRHDHE1uAC6/tCUpMng00z39M1mH4
RJL5VWCaD6lSl3l9WOy5DfZgZI1oD0Fwwr9+wDwxauc2MxswZcmIUhV7l9fELfwILy0LyFkiVXVK
D88tbPhOLm5TmNNxlTwgiHy2RNOCMM1XH4S6Vo3IRWZv1TW3nUOWFgtFO+GzX5lWWgzz5KJzyPgM
jsz3E1Ql+PncM061AtUKSpGiiv1e3jf0AtjpDvAgI7P8tyPvTy0Y5Vr2heN9SZ52yIAYweKvKnEM
q9YYRgLGieT6xnkmPVwSg8F3vqVb7NorCZxeGl42i231gXdtWTNT6mtuZvHG6E/HYrHz/GitoXNz
HihI1+6lYeN8ugdWRrPH4GD5hhz+yVhB/CRkPwACxSGXbZLqD8368Fb1I4f3tMQiRwCJX2Wpah7/
IpNx7q/4bVsaftPEvHR3hCe3oS+fHqYgEYUXUpMmzI1yRndFw4LIdPKwvbkRK+vNcKuZRgnzokuQ
f2erjt1FbF8YXOSKw9gOgF9CZ9RW2Dz4gLmowQzOSfD/3jRkPZ0aq/a+yjtDjYt2Aq6n9MfR0sRw
Bmiek57tQCARcUVSkFUIyIZZgGXWkPDWVU2q2b+yminDvfDOM37WvQ88WXCJ5vdfryjfGoiX7z9a
HZkrq09hwbqhL1lZZmtybNVV4FG92CAoTxa8sbtW4HAgLdz0CsVaKsKT4iZXxzi9RhaKxb/xgTzo
DUGlncCf7E5CeoDWF0JPyvR2QzSHSCpLlEEmg6ViW+ADYjsGgWiLQJ0zcLOH1Cjq3pbfCTgACEgV
qwIY/KXGeXNOI2pZe93LmU4o9Gny1ijlSPB2r+5mxFcdBMzKu/hjDUGN1KWnxtvfYQ1Gox8cj+Fw
ut5CuxxBrAef5jbf4bvqiLJfTOih3ykoZWfw8upp6Cf66yWPnuXjR74ufRhiulS3IL0ito10PfT7
beWCklJRnc2WOCOs4lynEwRKKIEUDI/P1KNKQT/GHg/OrMQFaHWSOMwOtLogJeh0368M7lQtbdHU
KYLm9ZdtS36yRm7awEdbMTbswRNnc/W6LIAvGg5bcDbVyYL7WKMsobptSR7ntLzAdpD2x9B8Nm47
CdcG30pMAG8H4K3ctnZxrbbE9st35ws93JMRkJmyQgPnH7M4Q4xvre3gH91BOrUt1n63EEyaOyCp
4zHih5gD9ERW6u2cNj6IlgQ9LtPgmajq1/GeTkyfmqbXP3iQQWRtMarJ9WnAFUm0/o+DOxPsyqan
BYuCUlrRMSDB/H4A+u+gAnJDMWeucfmQfCPwhGxNtBNveOvS2kLmKTV2ENq7aFmLvYUlcAY8takx
ky/VSF41wEIUnMle4GME1FivMGTsoClYfXSfEM3C+QKSstp22atIy70iyqGQk+Nki3N8E4TXmsiV
3KusR/N4Co+8n1STlAKM6NZts6HMU898AUkgzpQI7BjcJ/bItaf5KRNeLXmQ3m8wx4BDHIFHHNDu
8KF/9U3WFMlIfy7GH+04W/qHe4WbeJHYzb7BTdalvKw8ZYqYpie23lzNKjquR9k37mrrWtVSpFQ2
7ZOBP2JnkQqR5UzqPpp4kUJNRQuWrsyPzrz+p8kwjuj5QTa7vc/Udgho2vCQVTAev5dzmBEitoyU
rc54VmWoAqUtqy5EQExJlE3zZhvb62G8AjQB1SZsENdq6r585qJZ4YvJ5y4JxI/5bwxpq6KcSTiZ
8h5OyYUIMocNVdbGWWNSzwA4TwdRb2mMTFLdzjHQzJ2WlxDZHtdIxdJV1GfLpYFR0lN7h2XgYkJF
BJxtWU0PRbUP/CNcovBWhY3CnnLWtV7kQJFyodh3zVQQ9jxq5mXfUQa2Z8HJmv4NSQKoOnKuWXF1
epdpIc90GC+HLj6BtVg838UkfiiD9FtOmlhEEPMK9dsPV8OOIlzF0YpwGrgBMghFtMZ9qHk/JZxk
SDlejWTzwb+ciwAIxvCdq09WhiLv9ELyEBBDAjB/gCxqrtcA527va3Eh12O4yb5jvsKWu2VQq4Cv
ExgYHWdLTWYhuDbYxNQ6LIkFoB12exeZgvmkQVi4X3zN6LivlaYJqZrlkPSQ340nHkay3zEJtR0S
ygv0Eqv3ff0eF9rb4I2QJuRoDCJxfitzttekvSIH8aWak8oblReel8A1ujJc6J733+2W1+75KrnD
6esfHMD//sRZWZr0i2Tgm5AgMnppH3io3RelByh7xIxT0E54/h59vkz+U1QfUo06ypLjlwyM4MzA
DaOf8k0hMFFvIWlTzfvUe78rnztvzPT8LvXvzOMuKBm7mo5DAlQ1jbuxl/S8cqG0Fk0E58Gv2j4M
lxPO2nD1Cx+gfgSGskxzo7rGNND+UXK81WVn0YAylc2oNBb4GnU8YW5tzDCVjzwV2WkAkHGAqn9a
lwviMnzqLp9H/TBnW7shs+OawMpGooICRRj6KyXd1j8k8ra95BY9A8dEZ77he1QXuUtzsSoeGkjt
Yn738IGHRArrzzEx/dFj1H1ZNXxkGOFDetQzEx3abU//BkId3BK7XUtLr3Iix1m4W8JWoRqAt1f6
dq/nc8Cx2rZEUEo0yPoth6J8IWqZ1wLS/Ta6g6i+H6PKsp8NIXwRJmKVMVXWFs8g67vE6xWIJT+T
QrXRhpBmuQ7UH92QVuicBqP7UD4PxObIUSCtarUfw8PqDqM30yxm3zVjhN0MCCRy8C566JABRv0r
e9rruW5D7d3hHPceUr8CrPGy/HFlu6o97GkSgRU/O7SPYAEtjKKS5a3HTa9OKhFT8BYyRA57+Uu7
x/vmrhpR+wFsmslebrH55jyZX6s8/LxEJpu3Az2NCz7tJ6RdThfMh3/sWu5r4cr7MNED9wRTOiPz
//UGY8hQGWE+K4bYgtlfzutOXSC/0IV5zFKkpmmcHWP8vcfzjMmbcdOBwl5+Ud4i6ZzVoSdhrn4J
7XLug11qFv0mwb8eeLU4HmeLj0bOnMfV0f+RJMISrEnccqwQgDTbBl4BQoH/RlrWGIhK5pd+LKzT
+o9KH/jKA3i4IaFTI/QpDdYUjH1yLCsnh8hlsu6o41N56S7T16AicwuG08SzLYXxVYcZ96T8L29/
RQpDaY6X0tYxFKGHYBHmzJPyK14fZzVzyeQ1oAHS46u/Hhz1Oxo529tUeYkHWMRWMDcW5aqJwo5l
e9b53tfIEjo8/tryfGrKHpYvcxDdAkxeHkslW1wE38RhhywvzNiHdekE2G3K9gW/oAcyDTdFjZEd
65PaUclxgU6zd16oC/z5BHJlvDKmCJzLq2xnmqHDJDC7rRIjja7gGeb2evRGS74q3YY16P9x3TZq
WqBy1p1+5TfAn9c+uqoQVIOa6JMWusCqV/fnceQHZrz6lm+sD7w0lW1CiB9r3VxiTvyM0UGxKfLE
5XCEkxGhJqq3VmDuyd6REtoQ/toMaz8C9W18ercLriX9Ne24PXdxMfm/aY4QlgJ2agvOltDm2G9g
K9MYcmlkAQsuQsjpzoTbzB4AvCPTaOPp7F+t2+QCpA6/GU3ZYW9QXXdnIb60DdB5EHnE1vrwSkpX
a68TuAXZL099sWSFDnrXwmsRwG5mWuvmV8YfbtNxJvcPXeyRJZbeh0+b2510CEvslY43aCd3v+xK
MG43Umv+Ro2Tp8GeTmLRGchgTNOcLJEpDrLqu+maosXfS/mlpYrRPP43jVf1M3tq255UhVhvFwEo
oec59MHUcVnJGtkrYD5xY0KflR+CgP/keengn9TGJIQqr7FWB/fr31RUWK3S30MnspZ4LZK0DSRb
TatCGLjYKn66MswMrl0FJt64VXlufVxSVWctrKbnnxpTDX7SyMGaAOtk36jRi1Qj+T5oAAU+qXZo
91NUWhEJ9bi+e/kbiAotUrlHmg3S2U+gu69yuRsn9fPI4/pHlBLbUjSIM9/nyk2UVuC/4HSMCYtQ
xVxDgnI6VrzPSuByUYieEIu3zUNDHuofva8gnQ/0bz6ppBjtFo9Qo13LoRAGeX9g8HFZHE1hkjEe
GWzMkXYOnZNklYXVcnQo61ecx3RZPpYVaGnoVX2uwlmgO6dd97oR5vl4HWwqyetfWKXIHsws/THJ
E5zKi9SmILTKlIq/eezdWtBJYvTJbIK+/FB10A2BwnrPrYEjCMasWLfuqWkuCb7r52Gf2u9pZOPh
MLdrjRflZbAka8bpogUBVVKEJW4PxnaUld0NROBlRYvZfR29LVqjAa4x37dU1U0qstrZeHZrl50N
B1OqwmXepqh8XIS3K7qQ39DG1QN8nTKH7PgwYOtrURGen4IDXDDClb7boctrVM1P2jmfHgrOhNNt
Z+tC/aOoJ5xicdfAZG5XTYjzCdPsxILmuWf84qE5s9vyO2WUflCM+1/kJNiT5Ms5ZbTs1fUOB9xm
/B5AGAcwgxAKv2zLZtlgcddiuwDGnpJMa9qkYzj99eoixfaBGShyJLqR9Lm+8V3Br0WZ6MHxK3cI
E2kdkjefmc8oePm0YwCqkJaP7cqrz71U7UKfujzYlfvanskshyiyaZUPFSM4uRS/dWIPqp8j3GXS
iYPY2fVI9PFIHr30xoFHT3wYdplhtnZ0BOuAKQUzOjjwuBEVSJPVN7iyMdR7+qaEp7nXCy0KB+4g
L0yNr64ZYuqiaJO+TY/XOqdqn4xeKuVroj9ewFwNvvuQP3GgQXlpRE8fl0UWXiGXVcH5IuGq6v1J
/FJvC4NZ927Vggu6beeVoOGnsPmcbY1jN3DD/IbhhCu/03aN3Azkuzm1oLeZr2neCy19aRtGicXq
xkyFCBv9yFxDwl1NGRaZ5dBRvTZXBaMxPuvD0r0o25M22i87OhYYh6CZD0kXdbs+ypxW94P2lSez
5dsDPN6wGo/QocFTcnc88TjYfl5oQjsN1YJSH8NGtOaKCXYanGDdGnClRwC9KNgiBV+tXlLPSAbC
CIMu9/30XvcYwFGhYN6dE3zQ0aDoMtQ4u/DxNa9mhK0fEkXV5v92ul2RF0KYM/kHMY/vFz7VCtgk
Ga5nnS9G8eZtEWuWSH7AT0s5JGeSub7QGO11a1kxKQHrSnelCI1SSGrAqXuIW6zBTYeyzRI6anpU
TattGUs0X0r/SLVHesW2qxoEU+E6ecfgwNEM/svefvm7T6eLpUoDqZmP5NZMtmh01q5nGF5bcErj
KlnmxwGbOUhpTXzaxdkEBq0g/Wq4oXEfFUuSLMhNypiwsn+gCZ7yFB2PUBLidAcUdY+a9V7X3Sco
6xBtISASyfOt3isHA/SzmwibgW7SR39slsDlhA0u4ORl0JcQj6tBQ5oqBpRUajULE6xWZVu4iEyK
tce3u5CANO0tntEMrNelaFVy1w9GPTSPY9lGEs7kXdY1eYP49+l/D3iVSmCe5P2Or1JY7/bk4Jfv
XV44CXjQof6Es7oz7ELjOB3KMqIH9gjrmX4BTbaJj47uI5tgUSEEK9U3Kg6MpqDPfN1QqhYxp5Wb
8OyXKT9J24pphP2XsK+x34ev4lgvifv6OUH4du81WTGYBaVY3HDk1y44az1bqA4M3L+w/DD6cz6D
Epbjxz1m4P16+Py/iG9mdQ3CGzcZPEw6Py7Ccm2oIj+UhQfL4JGBqwZX32csc0/5x/zLKuJ//FDT
CAlHaykQq07Ird6iD5wwOhzNSK4qMMmK6JcKd/G+2JTF3H5p9MiR+2EA9abLKNK6Dnlin0jtojbj
5HS/MA/mxLfC8lWsVQF5RKV2T9Fhop6S3AfFJ3mgM+NJ4Qvv/BBVrlMYtovmq7jWYEwCuWpW/k8b
+h8UzPK74PZiWVwoc1yT0ResPAmTLabmyM8gjIBe8FkNU97Bn7T1aBNtWSGqOSpkxFEutYuO/oga
U4l4PkRXgl8JHivpxh37ZXanK++ML/fegWP1QHzvReEmTDZGmaLxAY4b14TVGx//4rPpu1HkXI8J
TLEMBM1rezw1HnYI0pEFnaUfSaO3UudTu6fd8UQx8/n7TuUgJcqTQ2ddZQn00nl2LZlM/BJMQs9H
8gV4SGXTu6At1447CloI4PnhxOImwFw/9xUIcxSr47trKm5/fgQ6udhEU9012hlpYYP4WsA1B50V
2wdQZl4RbYxfFqsPbY60ZIsFkC2bEXdtrXSfWU/nEWYJNLwrPrwsSRarXT61rFVUTYrcRQICRWW0
R+7aFDolNHbacj1eHToQec8htYlFQdJzU+eOQHP0Wivcku4ElTGS9wBeXNBJONz1qT2BE5JrFtBe
ksmRx3tDxRfDwiWFefT/I7qLX0yT+8WGi5pnE0lAObKiis75C2gRZo8g8ufTI6b29oQMG9SlOlEi
aXFVHY8fPtd56bLE5LN1F9gK1OWbeYaNAQQ7lWNG9o9+ir8m0K59iutvKgF6MkvsTclge1xhVzh+
61YP27+WhceaMI7rZdsEfnazC+kXyRqkMgTK8H5q9qCliRrVxodbu4p2DBndfcJ6AfFnO5UY2yDy
HcauESeWDd+YKdn2F3TwuZubEvhONp5tTfGSC/cyNJYGLCjejwcXxq0YdpKhXtCS+f/TuHaSE2qU
obJX8LqlSRBAZWH42pKus/DeXq+xTgTNTIaNp5+pX9rVeFoDjw3uYghy6eY7qayajNg72Oj3bRfN
d8/hVG50ezMx1tLxwmyhKDLl/bYy22tXYbxxz1MMLJr8fZrPZlTMwU7xQh0fJJOcr3XgIzBxd8zy
oRIC43A6E1RAPkD6Ed3PEaRnFZUrLeGFkVEPnO8TCRufdCUOb3K/F30NfzUh5Yic4/00HT6x8ySn
ObO7Ruy4po/uyBr76QQ178q66tJ7Kuz6ZsG5rTnIANV7oCBdCs/xeQhPGxe5otPLPc7ye/Ha++uw
JVVNhxVi6Gjb7MFuwhwN+PoE3GNnpD0pWOihwZvTxuQkrQrnplGHI8VtSgZADv+2gAZRQhNZeqPx
a0dNcIwIpy2cBVlNr+f+tcrnMpxItvdPt1n+UGWywEf+P2sSRKwbrlBFsp5TIPSlEcqcIct7QpZ2
Z4cEGB0xXzqga5iDY5aCpTM13+ZD04m3M2brZDObEErChsFPHODSrwMT+vywDmUTB+kSx7+6S92A
t6fOPTv+YUAskluI9IwzdS26nt3hOAQqM89hTLLK1UtkojwjagvcfaXr0tp58tpcbNIHv6rW1b3M
Wrb24K3SFcBOLYB6zCeRi5kwrTTyKRcBUCSzZ+b2v4aLV5QH3yk0Qq5xeoXlIBilofX8V1PsX77o
ursZ4ykhBAR6icw1Gdys0KGlCq4NQtdfOaCpwlFi9T98QDbY0Fu98+yU2x5TDNj2Hqdj5BtD2763
CLQUca2bt+6j19bXZ3oJWgajYwrM32PkP+WG2eMTMbN7EmiTxd3X2EvQV9m6QouRfb1OOvYnMVUZ
nvWwJSGcvxTczX6gPjXj0qUKRuW5umpqaioZVW9P8WZilLqEGhb7Lxw0gf2u3irYAR45vUQqIJhe
ZpQgBkKKN3J0x4fb3sEgBB2RIEejEDywAYwD1MYI6zKdIEkskCCC/ALbqOy6OXQ0LWRA+d3cf8uk
EoJT7vEvaUFUiozmGePwya3RKJLEhiAdKPinMDejZupjTCSzlQ3piRiKH/W9DvFdeKqsydSWQIfW
hUacyW5ImUTazy+cTPavYIelbW6bbjpTTB4zeqXvrY6JGMSPyszOkdzdYWZ6yJujGvM8UbtgJ4xt
QGF9is/ozINXE68I8HdsGkR/oRJJBvPRnrQoZ6W9z2ICb3LtFlNa1Tn7GUg/uOoOV8jNxpy/+t3r
h+7ABQIZ4lkMbgWZ1UeGhttOhm0CxZM3VEcnTeVI311ySF01EQtNPYyMTCVaOIiiU3Q4b878Irvb
qWn1xB1NASVN1WwtOSDH8MjoXQgKgNawrYVv6yiOzT7HhdZ91nx40GQmOQMHs1C7syxErWvjKll2
2FQ0uzUAVZ+/nyIf3PT5EtNyL+m7/JpbxG0TJETSrX/cOm52tHJ4F2kJL5t+apsRFZqKxqVfDmdo
WENPF7iRTEf6A0MyDiqZJJLYDq413ji7Neq0FpCpaFR2MzZP74911oKSluOzlQlOlVLBA49vDGwt
wafMeoxrPlLNn2xhWW+gdU8x62jB6jwLjnn+Joue/hYtZYd7mVaGYhrfdo7A9miubAvurPJamhce
LHfH+/rBkxvCEJfDzSZRT7WIv6hXBcoXUQHFy4f3KhUugu8zjA0V20ERXOXDi3PKb1YDLWYnni1y
NW5PFq0k3Cu72pbbVHioBP+v3uyIJtCrtxF+09XNiv1K1irCkPc5qv76Q3TVb8P+4Nc/zAtJKCiM
X42BHm40lgNmdMHVyb/8N1MHf5sVLr7Cav9fNcUbXS9VbzpB1CoDDR18duc9PDsr8P0hBv/ucjl1
18Xj2sxj78NxzEqfEt+IUDj7hbzcVsYs8eEH3EG6phItH1fMKPSor2CjOWtUngUyD4fda7bK5SK9
T1mqGjanChDSOXBjs3MNIjsBt5LWZFJD7sBb1cEEJcTwM5eeqYjA9niMFdgcsdHiLAFymBICitFO
DlqkiP5XlChFzHhNEvlxHG1PSLNk1OkrevZf2bU1qvwSc1l4dZt3gN9LOTi6JVmM22jTwVBjSki6
Cz2bFiQHcGmLv4qDJV7uDmoiO02o3w9O1VWwJXvFg791K4dw8HSXLnizGVKmuS4oKkEw5hvgjp/S
48nJisoogpFtFhppBPrUCppF24GClk1Uc1ianILlPI9gyazFwCgF/2F+Al6WoaawvEXhOXUZIncO
UqgcKvVmwAypr6LoMw0IFKh4+iwfAqyANzUeLrlFanbq3V4CSDzgkLy+4MkWHc9ypcQrf202WBAa
/Z8C3M73z4BNIm5xpTgcDBs2N2JqULUWl6J5EZfx9LXa6oEyZwDKBw76Rw7Ve1GUUFV9aCwZH3Yp
X2+pGaE4mnChnvJ41pDaOnGg34FLcRrKNsUE0+CKpeParztziYY15aw2JzEZqAaxHqu1qLXt+9kk
xAvX5mIuGnsWmuwpIVvUsPr1JVGbqQ37RUMlSvEaMgkQi1rjiqQpuAMPHNYoQ1ZkNUC1xmr1ohve
tj8D1vEqG5aL5w5xOYmsrNvraNqclzE47JNfLuVVICTXZToX0jprnwqGBNx3zt2s9XIvKSuidWcx
12wGAP2kaWY0yLvHFKJtsx7E30MC7wont5c6Se3/8xUVkB20iVL9Cb9PaQ8AIfKcWlb99tQNcH4x
c4+kQmrcxXKR9yx6AJ3BrlB34R2Ge64TN4kRiZbmNh/Uk5XP7hRRRldR7ovFdG85gUd/uOn+h9X8
UTC07DpuT79kp1ClhefovLhJfivnDRP4sbQ1Jehk23SsgnKFNIP/wfD5b0YW1mxrZvlpsfVLOgEJ
Xsis3lgCYmzwHqw3mLkr9/UKMSOls/cizF1kkycKZN7tfXUrbBRFegX6w85XuCMn0zh0javMJt8e
cxpMQzDAZ9shI1BA7XtrcVuSwezVBehyjrYwIQzgQY8g6sayNa+QwPXI4xN+rv7zF2+chHDesCtV
5uPNa/rBPYDgVqJjoDavGh46DEwBI3x5UuECSvnTptoTmdRrtmabgZPDexXTLIuu8D8L2pFe7Pgv
+nU3FPNFUcgF9fw/QS0gZrD+myfX2+5ib9U7ZYR4hxaGmqCPxZtg1n3NXu+acDXOShwLzEwrA6ZS
xINajScEPbc1V09GaWhTvyu9J9om8UMZVptBXMOeg/zw4RbeTYeiEaKSm4rn0bou2RZtF4LawHTJ
bZsJfTv3tVKFkEabuJ3aZz5FyKWNq9zZTl7Sk363WjaiijUJeX4qhVkObK2yD8VWCntjs8kkO7I5
GPIfcIGyJcAoqrEBQpij+g95MMwWHmPyXd5EhsLLOZdx92mTvEzbWW+Nwu0vkJL89d9yRulLrf/6
0D4gvn6QE0HhRmEiDThdhF0ioKHzUUEfDJ5KgrSUKBdWwSimgDuZGBe/LEUii2HgvtNtvCb8dmJo
uSLf9og37GShVdw81ft74eN9cKNJc7/DfMEGJs9wDBliy5wGugiI4o+rGhugHRKZHEQtU1TyZsB2
UYWITnpQKP26KR69MQaXkr3hudZFeiRv3Iy0uoEejjpaw7gSR2ltME550BGEyaHK4N+6T4Gcdplh
24xehSYD8H+jcDQwocEnUpIIrtcq3dqPk1As1vxt7oBsBrAzoKyRqSqN0ezaRRe5yoDaQ5TqDtjt
gsiNSSIUGzjv8JP1VHqYG7Mth3+gOOgF1XilAzoaixfqFafFcg97EuYfd1Svn8qax0Kw7kEQU//k
q1KizACTzxKafX8a1dRqrKwlp4n87iLQv5igOJozbqKriBztgZ5mwc+jItO58MKKyaxNiext+LSf
F2LPSM4APYP0QLqZ8Wd+scEhJuF1OYVvllsDMFokwicbJ04rKqIX/D8maiqsnrsw/Wl8zI0sQ53Q
oe63z0y3HlDb3unanEXVR2iEZHLm1S2ucIqyCIGv6pE2nMrn0hvwWLcidmektgncdcwbv6cP6gPe
lQh4Q8m+XrAf7fefbNFpR+ZldbwdWlOUFrNVXFD4Rfi3UivvsiVEZzUXswQycaeNeBJgEVUK6u6l
qEigyC8NgewVqLuUdBceNNAbHdpsRRwaLO4G5U366e6nP2gtvHdp6OuCsa8iSf1ejdT/B1At3H54
da7CKVxay2toQyjPLsGK3ZlJjkWfCteg/Sfvh6RRQYRbf04qb+Rlz42W7FZ4EbTC3/E+uVfUQjn8
0qJxt9xAec8gB5QGc8+uEVn9U0r0RVmz7qikDwQVfydbJUJQkoW5oFwFRmEBGvqGytsNqojKcITl
Lke49S12XThQRoXtA2ddThHDSRSgah2F0Dto5s2z7ibHlxhiXGRCq1K9KpRW1HDR0n0pnqAzSpoR
yYRHmt67VezJIBH7KUEO/tOt6SkCBqQh23BM30Q52lCCYHbeN6h1+TGrMLajYE3cf8fpqIpc6dbQ
fsqbLY0sWd0d6YmTnDZGZTWZ0/pO+rAcogopF6tdhcCRZSJpLDd7oHaLHRJo6emO74Gg1QLOX3MX
JV7+uQCcrwHH2QBDY1GoyR3w9flvHKae9riP9YtTawZmT6P31nbT29GCQ75ehMokCKvBAthBnCKj
VG0s1W0BbdBh2OcINeIACMbjcauhV4gO84V/ORdEVe6CT8t1QbmwCgeCk6+T5a4W0I4gkMyTD26R
TLGSfg8KyAz4zcuS/zcY6r6+YHV6XIUCdC1wEGN+Iv5w01uYe6qFOc+eFXN8cn738nT7mZOdfZIw
dzs3Av2kFhhmf/aiGhqPSvvbNP9TLJE+OJ6UGtxJwQ+HAO8G2S4moZfHUqttqCfTvARiwX5sZGKK
qMVLt3NTW8yEL20EegU68izXEk3TaNESkTF5O4BI7qT8gbHpe8NcYKaqvJ5hie2KkZ638b2XN2CW
PPfRdj/WPhU85hx6Se9TlqqdQf0Hl54eJNxvcHw6o+U7rnLldJOidc1KGb8F65U9vhdi70W9unLN
XnkQbbwOjPgTWyz6q6inh/CMva33CYIr8mRhTgzmAmP6myNYjETsPNSrcLA/0E4kzSPX+sVWqIiV
2J4UAQi9fHh70Y9Rc3IprQ4PB5cu2ndeVNTBI4/SJXsqGy9rpV/iFBeQmT9epMbctXwb7v05ciWD
vkiC6011hapDwF/uqCOLniS8rmbF0tZHFgkvOcfHh1Cy9OA7F+LWrHW3ZaJz/3zv2mbm3t+Jiqr1
IohcWzKMOkjgW9QuNUFPSr14zGBrqCCGufFi6g5DKVFSDNP9Zs66sWeqznxwmw+m9ZgCVBy4lRYX
R66bv4d8LlX+IQFr7KGBHQWME/qgUE57JPYZ9q/IDSm+OFt0IXxGSBJkg308JQU1qbd29saItyU/
P00/xJFDgVV55itJue8Wlui+pRSzQ48NgU2nkNU8jGOp9CHTo9nQNGnD/OxJt9DzG6+b5mv7MfMg
s4K+LD04HF0DAxO1aiisXJipx/+VUOEYierIg3wxdTLlHB9PWTkfBjYLfZHSIw3sTuHwlMmaetWE
JJQ+tQiLkMroxF9vEWc9SkWcaGS2N1ZPV2fMpnY6GA0wMSy7V60w8hfVLbRJdXlm5RuByYF4dGoH
sq5w8qM4g3KMbzlcN7gOhxO+S02imfjxmWyFFp/dTkpvvw9DHH44w5UX1ZfRZgfmUCbZPr5ga7xK
ygkkuVx3/ZHIGyU16uhJngVu60KBrz+rI1fBulq8ABuUZ38/83OTI2HjE0axHB3soSgmhjNs5J36
DJeXyfrSoujzA4SSfyZnXt1/EgjJzPG942fLfCYDZ7W0JJYLQR/j37NLVvRWmg2GRTKdiTe9FwUE
JKOjYHxCj/5MZ98dilrXO8NHMjB+8DDTHG/gp1wwR5CUlEEhLOaA7ehKsNM+Foa9X5nN/Dfcej6r
KsvpN+FjNXPjRb9URjmMM2vBAAJTYXvEadwgV+Wk5lRTXL3lOv/RGhh3sL6gEfFpPUVBfoDtB0fX
kncKvQ+dIQoJLWgk7r7U2rj0p0l4n+nWoteWGIMSseyh7bVrTE6IcBkLp3EO9+vTBXnOEl54KRl2
+xneEnHG0pAXak23FHXSKvsADyMBlATzd09AxJ/AdwbLx5z1xa6wPsXed3GG8aTp45/lW2doajQq
Y/bFB1ZthY+M7lDMjYBN/XFKmJ47sVteTCbcdVVbujWbZKAHlaU/tvZ8fJ43VClYEv/AjTvPDYen
O9IAYq9vTHqHvowDu5x/aMuXCZhwu7xMMPJY7STh9c4CRWbAnBhkzVgbyoqh3cEgwnzkey1M4ooQ
9GQI4qGxS+CUkVrpouGJSDWCNr9lEhghQF9hlO/XklL0osa2ZW+/CQ8eN5cxmT2I1I72/p0TAQkO
hIpOu/XMf7+QvNv6VV0AbjffhZh2zWzfRRvBvgQu0uy56uPie+4CEMd29f5GY7hhpyrRy35U8T/K
xH+DiHiATGjUm9dgDnBCMTQHOCCJu0PlfWZ1CDLyVSilTtWWAKHPY3vqvMURL7ctfQLiVh/3hcCP
8WoXM6BncAEY4bPeS6KVU0ih/RKBrw0nRMeofn7kRWVobjHcWvATnoJKuofqFTmD2lPJqjgk1eET
ukwuRSQXaAYYe/4BUWcdfqdoLmzam5tjXRR6eWJIuFUQkeqZwOOwwtf0dke+AyImWHBrOMBJZrk5
zFDVgssNBiCbsVaY/QMePyVGANcfFrQDdxJ6wFZTxp/5nxmAVSuLVdjoapJTbhI3Ua3sX9DcYG9P
gcTdUaaVl1d0tEbBlMow//AvB+v6aVw42k4jCly/rs8OyzXFrsTli9PAttmQmRCF6FcaMRIbOA9+
BfY/fI41J70NbW/3+S7+ecfYTm/dXhjm2uwKyVsD+ZzIc8G94Law7ajC6pWxwn2q4h9FKxrzvtyU
R3BuyzmQgLv9gWhR7R02hpKyXQIz8Mu0mHQcaYiouFmUecO/QAOnYENn0ukLCBn4Ds2CcxGapLb4
M2JrI9WutEXFyfOBGtJAfHoG4RG7ULqkF//cs6wAaHH8cHPcQQstoLNwyF2S+y7WvsL5CidC5KKs
patDWRmRiiWEaIj73nYVwYLnaU3KkfNso1OYyJuUw0NNeSbbbzuHxuDfpS+rL4xieCk02IWUcp18
bYIu6LYyMRUdET5yOp3ujShXTnVabNaNnp5KbMcLzeJ0FWsu+uoTfuAZK1RGfaPIYaoqzBLmXq7w
tjCPU3Dqy9tOcGajpXANZubpgH4Rj/zOiV1V+58vL3vb6CY0zhvFv/ADH9aKBesA3f+mRfku49rI
GDMr/uN/Gy6YhSzY0XHvIBzZEUhzIbQfN7VZMCnCuLx1Yd6GPKDwIu5NuWPnk6EYOLADYXdKqnd/
+7bjNotLRaPd2AbdaFYkSZ9p2rdIdpvB4uOB3HdRcD7f1dBittrOX3tyuDNT9HPcXtyG4l43bEBU
eY0Dou8+w0pvbHVvR94g0ttBBZqp4gGtYxTEWWVzsugDsdhOW9AZOEFIhuB3ATflKES41Pp6PLd7
y7+VRDbvkE1R019WVWgTIdHexGh27Dh8Uo+JeycU2jcFHB2Q2keVGQWsdMeKcPYBTxnDKjPe5J31
5s9Iw23Noh/TbDuVIkiitZBY7uyMmIaOhDeOd+Iqv+4DoDmk2H88pGBrLdDHApuk3HGG1aABN/1X
a2QXKy4JeJuuznmiN/WPt90ewLBPUEnNh5UWVNm8GaP3uJeMajILFwUO3JKVNYw9Bj/56J2F+bkd
vRCDf3k+7iIKv0OAJT/+A7dg7UFP4z5Y3h+EKIm+yv680bLNsXcZaurVuegqVfUY8d9eSHK2r1y0
2Bc6sdXWOs1NqCmO8tbTE/H3ulN3GV5uEAGubk2lzrSyZzS8XfJlx6jh3P1hMlUMbc0sJLXplNB2
TZUPhMqyv1AZCeUeGnwoFxaRVBy3GNNUxHOsqsPEmg4rbv76cjh1gwzlYKbrl70MXFKUmnC4u0gp
qnLMnY4z8QWZVN+8F4pEbADjD6Lx4e1DT97RD/XOw54eXfnBaDGppucP0WakfYGJX8RC/F9W4Qcn
aqzY3GAaaZikXYwPdNaQOkV+S5CTZukJZODLqf0DvHdWDMdo4JWmQH/8bTGbLzHGvO9lqSBaTZMX
XIBFS087ZpaLtP8diiP25Q/YnTiep6c9h1i6FTydpgYWgysbcvFxD3LS9VxE1ne16ujz7jDfyL7x
riKGW+7YCCsfec3cSB48MgRB3HsH0018hQTRiO0N7XjKmxU1KRRWmsltZqHtBMdiLdDg2hi4eR/p
a0nOmpxcMmgY+064dR/6t6G5BHen+jF6T5DWP2Iu4diG4RbcFKjSQ+oxT0IQUGLFTECNcGYXI9rK
N1FS1b8j9u9mB61//XcBgn1EdYkIAT5PbBfftD4QMyCh+g0ejHYHmAMn9nTOm65BjUFU5/O2peIW
zFH0l11qdtjN7RLUMESR2jE6BMAdprS4/UzGOb0p2ogDwfcpR+xMBe3h+ULTaTuXXKxOM1PyiWHW
3hzoEUNykPoXrdETmtnGRu1Q3yJDiApBZ1YgoHtSwies8Kv9Ji7NdkeAFndGUz6KW14sYi8C5/60
cbZLFG1TCUYV6XSgakWFf8dK2poUzjhN8WWitK3FMcvSz0EliwahocaPkdNpauqojqIrUx1uBfQR
BdbCIfQLYgF/JdlZWqAfyBAydDqu7YlbCXsU/6DrSMMejlqFfSaY7r5Rr9Ijod68Po7/Qw5siPQS
pwl8FsSyNOJKOErNbQ1puii7c/H0CKNCCui8xy6Xka7EXfG9Cvw569QMSIcmz4rRNW6zhi8onrcB
yjCqAbkMKG5vyQxwVcKXuvxhnwP80JgVQmOZR2RGIcFkGLtKaxTftOmlCARJkGuI911cEuUTPbqQ
qtyhW42JN9gPIUpW4a77HdNnfrg7ZyH4ba3QvkXsJ4OF5nqGlCRTk1b50qU3v74ZTZHvu+6SiNpO
iivQ6FMXTtP6x23e6CtI0vTLVbm3qbZv5mIqNPt2A8CjQIKMmyigtDpehuWeVrkIQcADRYTDMDxu
xm33Qka27nrKpLzlnq3Xt+4lbVyIvPakK1Q5k0wNX91KLuiIoT3Pjhbtd1HdyLB6CjnXkJyEzZa6
paG1a30zPN/9s6LS/M8ajBd+74PhQQwQPlTPn4QgrjKyOPd3TWrv3h9WusABwoEY/c5s4Fqyil/2
V0hRJCOpyR/5FXl3LjHQBcYd/1eZyFT0mZt/9bzplSvDd0L3pmiDAcyBVqX/pbrAGyKVUObtk6y3
vB5T8UOkxjAsAYIAB4hlXpGl01GT4/JwWlanSXv8+TbLlkpd8wWs11S8Ft4D5qPckv+9XeHNmuUg
IKoXNh+1aRL+c6USWGCnd3PSyke7NohLNYohjNgCKQLiWrf9v79ZNSRlUjOf2OiW7OnTfp8mZcoE
3/X3Pzn7vtrWdzmFoYYeh4JiuZDXHAkuAtfMcr77OQPkLjf8C+8btDGxHLhg3jFefWqUUJ1nBHNC
vdTB2u6WKwziPRzBTjwhkoX/mlsWxWiUX5e2cqUNoimHsmQv0gZM0K2b3iir22NUEePpK61LaBkq
fDrzgBEwFflrghbDT08DN3VVD15Y5LySBcGXVj4mcswJ19QUYph/BTQkETCZlHvgkMJCukkYDIEZ
fRWNy4z0mjP0qq3GWrxSvn+e0PD5fFyDHqV7yrj6O8n7TZEp5IcsPkbLhPjszqtWG/Pzr5McqFJp
z71BO9rGosqjQdZheGWGg7AIjjRqBav5dMWxbQqmlYIfpbtuBx+++qur978sMRQMcZqkgJIxYTKt
BGkC+Dbnvi9LOI6ZUYR1yMmL9olktQp6L9uTVW7nghgWbtvoSAuM1IX76I2hc1k0+UoIKtXZB889
OSxywgHZiLBRaNWKvQdRgv/O3mT54nqkFuFrkhbjC7mBzW/feu+ZljfPVJ8KjTxVUTqwF4M8hZQW
wazGODmoT5K5o7Z2zm1ug7bBp/ozAHofr1Sw3cjn7LHZxTLUPNDj3e71trhkeHd1UsAOamJHSFjX
Bu3c/88sCPvMBdeWuaXN8kzCUlj23ggpgh+7S5yDFOBkEdrAQRqQ7RmsPYDotbA+HWhKrSLou4me
8fhBRm0JgwVnIuRd5dMbq5eZpUptBFAReIw2YmlgMbOU5NYi4MJ1ItWnnXdzjn/DRI4/Ett242wm
zY65Tk9OIgB+qtBN1UmnkpXnZVh47yXQ/XpJJTPGjFtTrTG1rgNGzS8B6n8KOWfFZg8vdjdhFMoV
P/kR5NhorVzFICKenyPZJTEchGHBo4uKQNEWxLo4HAdxD96EUWVVTPe3Vq0eXoAFEOKR4ngPAe5C
IkMd4oVnLCkZbq6cl5D4ZkRgzOXKPcg6xjXzJx47qFrQMwVvAcSecpwM5M/j/1k0ArXC3qRs+w9i
9o1QDT3MZOATxrIZCMcvxz2/luzCW3eVHU82GeBNt6DsSI8m5X9/Y02unFsMHj0qlMVmTdEUP0U4
DwLeEv8qXDo8+EtamAgLomHChFfe9B+7GrKHf26Af+bBhkPDvC27FuXCl20wFecbSO+S3CgvJZSx
TROS8zYHDF8HpP8ixrmBCCD8EmKFznl3HTGrK+Xm1nr0EFSxQ2aVH7hVOd2H8HMDyq9chq2cG79h
6Aa7GQp7Npo/hQe6njcD3xoY29dDJWm59ejjAq5nLDV3+7wNLvN37yER5Ls4erTtkXKJPBAWC/W8
6iQd6/Vcd0XFYuvMNkfR1KEIw/y6tSsL6T+vOWcAzYjSgNmPPTYaPNwPteOQmZbdC6Qi0QLJUQds
4f4tk7JvID1fSew2WXtu3wiz0+of7yFENhuqFj5uo5O1AOqXYkk56sMIPEd2ASCDQErppowNM0Ud
bTA8S/LWAvSfUTMk0qC9BmuZ1LDcZ/1hbAfaUBeHr+mOlvE5hCy0sUtXQ91ebjzCTUHyhTe0ABHq
eCoKXLYUv/y6zOePnU+MzJYzBN9ehisesnbICC5qq0LnLhw03bhzQEtzq4S1kAXAkEVR3TebVxTU
tjeYQOzFTzPb27nHx4xe5KfWjoN6+rFeBA4+Cij5upcUF/U+ZzccEI/fs29/HtaEbgvTf5sIXR1p
4oKi6AELZweowHlOb83rNsYQGh+tGtz19hRKY0WfkXcSUrrFr1PBkRBEidisbMOXbQmVxF578exN
rZgHnJ3yewAiij+BEdroomE43LJ61x+kmq35xbE8cSSzvr4ZU+tVe2YcEtb+qRj2/6kHj5mnWGKZ
ImPZbZNfuz+qtKnpN7cs6WoH0ccWMJIZz6BwI5Os59z9vas47IuED35//b+W6Sb0+sCe99wri90t
dkXgIk7lQ9SICpUWoZ3X4tFHcbQnQwYhS43ILqAyaokP4cN/s6F06GN6mbgulAQFiqVFYY2P3nKT
luZMNKuzpScRg3U9VbzgTACCACrWauT2mcBjZkWkaZi6ZnxCQdS3R3O19CI8Ny26866u4qTpJHfL
bsrN2D66lexi5hE5Jl6JGs2Wb5CZ7HFWYCC9E0I4xn6R+mkU+Qx8dbM6IO2IQBCmu4zStC33d14H
timMEcBn8tzsD8biA0gKhiA8A/Zp5R3Sn8EeaafDmT/rTGVHhdKV6P0SkrveJ3Q7lCSyzdBNVYf3
MCd3sZd4nBRRqZAdbbj7F/3aZC2eo9HBAn164GTeN3/pZXesIvh3Y7CBLrl6lvGBqGUAQLGdej2n
VMNZeqtIMr3+UdnCDOT3XNb3FEJ2gsRHssgUbMMydyUvmH+xGUT2UFXhMfTlBEvyRB59d+kchmgB
o9bJ9+Gvhpx8+qBeoUM3tXT7g+aVSHqzo/rEV4ocJPkA8bvwB0iim5hR6QPGoPmg8gQjTWuFwm2J
YK9HmFAF/oP6/+S3Qq8vyzt9SPNTggq95XWbhwBsTaa0YEGFSvnsj0Mh7tXQeN11rDLXm3yLNz0z
FdcuMmgxfxcWa0rr0WoZNyEUtePBtSZYTCl3zn4EivuKk17Sl4CAStMv7t2qSbV07gEMKwBdZemS
7pSGR/AT3I5DMC5NNSYF5lNyxYTNlBiOSLpQfz5KFFsPAtUSsjEu1KscROpFYHN2L8BOEsBW6cVs
SvQJhtQxHIvOTePuRvtwPvTEd8BY9kvX20iDU551MYS0FPi+Pdz96GnVYBhfBQc17kPy2apW4fNS
LgxSkL7jLkDBGqD/cq0O08iSK8SUWS6CJtFtCrhqD1Bv5LKthCMeW3OQpn4UQ0JY4RhTp23bo7tm
bOgnpUkpeR2ipsOmHYhCA4IYg/s5GJ3CWk9n6MDHO1kIt02cZN/rSlmviZ8lGqY0LKconB2/TbWq
ISDdawkpmhJLR5WRmGyLLeyIE8bfV9ErR7zoIoub4JfJxyuDb49JhUwer61YKqDj3+Vt7hWKU4kj
2s0m9WGJscBChR6mvXbzHRuO4BUeopxzlDak0cAvp6BzLjjUDbyadFBiosLn9GiDd+p8jyzDIE7w
M25xEJhycPwoIQpkmQvI/V5YTNmqSoq3ZtPB+u3zyUmkM/8ASnxKiOKRx/yfCPJUy6j72OWf84+q
evjvFS2oEkQ6/+kdtGbDpYAhbA4dGgo552+ppg/qS8GUZVm47IwzlhdCxrDA7Ld0AGbUO+IVHePD
czM2rE9JFUDY4ftdXxKmkM25oPzUMVGPEysOOEP1NR0lWZcpGv5z1/TpzC+44GnLW7ezTuVhRbHv
JtX5mAAF73HSY2Pnb5bsumufYZPh4WzQDEUM20ZmwpFVzaGRrkeZnt4ETISVBp5YFD6xDjj8sCb6
lb6ZyMmSnDH++zJWcaF8yGppWf6wCMkYD+i9DAuqMHnQYApRUe0G3n6I6g4akCKp0ebdhYEAt8bY
UNMU4CpFL6TsqfPESpt5LjjyVJBaIsdKtiEkqjE5+YFeP3Bol5TRYV+mIoqVUadhelLdexFZrJeJ
pwByQIDG89LkPwlnx5xXvknRIml105/Qh7bNIViVvfRuu7Td5eNXYFz2Z7gRM2RccrPS6vGF9iYE
9LwEvnN031MC8Q2FlKtemPWDCQOaxJDeiBN0qO5WTn6G/lwWzKyBvrt4BFEE3ZkZTmnn5Ho22CY0
+AI2FRAJweyV/X1t99FuCPStxTSMYVts18NpHGnnaGNOUwTmKJhlxywQATcth9itaeuoDZi649ci
bmTvrLcLhQBH6Wi2X73ufE2rT3pcQHtOUAMHPQp2bBsFOZ00S+2obM0FBzg5IKtPaMCSDserC9ls
t3Z0bVvWMrPnJlyOmMTZy7Y5R05N48+8Lr211mxczqfdWcp4xrIirdal7i4L7km7UFO3TP+jF80Y
9iWVZANIo12xeIIXnmsvdNq/9Jr0DrN1s0IfDmKZHo9vh0maZG+LrJLedc4Lxrlmbqg9Sdt3C2de
nA0BKBfCOizpMTy84QxEM24ztRYQpsuyUplvyXWGQjQNnxPJyUfNsmuugYsl2UFGuGNi0OgIB9Bk
V09laY3G7146KFOFS/dFYcVe+CHfgCVjGxsO6NAeT7LS8USpNXAnLFpgCvaLfB3LBcYlEWie+oww
duGx72mg34IB3ClxoQDzw3GHwRKGNCHTaeAmfVEEod27GV3Ft3vEYr2Pzo+2HkCNKnSETnotXW9v
vvllS0xn/7geKJzW0YMSUMPA0zytpDshGCCI5UYoUPdwMH9iW7nRp28PYjScOx7/qkOg7uncPWJV
RKT7u85Th4QOsl8lMkHroKOVHsOHfyCsv5N4KJnMixb6hppKuv5AZklgkMU41h1uYV//tcnPixEN
fODYfieQBGechIXQXnXYHVT5nZxsyRCrHDEIlOrZr7rVCOV73873AXb6j5i0+YW0Kz1ilS9MuH2/
GZDomtv630eb03Y5rLkySgf48+m5Pz26834pkdFT/WL/j8rfy2rwHBSoNHP7+loqOvLFqBU3dOmg
Y/q4Y7pMCg+5/UwEIidJK1DE88DoAha6M8gPuNZbMnizts5Y9fG0zUAoXRDNTkehf84mavBjpIMi
35HSI8nx1txX4lap4e9gh/PkuweDKw+akK2i4BpTSGBo5zeJiExkmy8UdAe3maFueMLcqHMnzw6X
F3YyOoqk1NesZvncHnhF6xaDvQA/4uVb1lP0LdRKc8nAtce28sZzNLOnRfLkQdCOflgD0SJQQFhF
qqcDcBvsI/MAHp8wEA41pg4YGkfc081nQnEgYMPRr+zFSge5Dnj9ry77J/SvTWE0ZBgW4OjysOEM
kyXI/NmwSC8LPeV1vjOlCsc7e9TOVRoNhTJDctZ86m6OA0nejC4reP0RCpLcn9GwFlnwde9qcKjv
xH1Xzk2yxIqAoGu1iKF5vfpodCNNHKmExtMLeCd1HoUfcRzYZytrN5CZtPx+/zMFX454rh6f4Vw/
trf9SI12nZa/hgZyvR2aCXpXG4bOFfUu4A1UvSlJjP83sG/IW0uI3KnXnKYCVEe/8TL4uaQ9ulMT
uDUaCSJey/iZC6Bfnx4Boo1q2uyiFoWkTPtPFC1Kl2XIfyZ9xs+Hl66fUGEmb7GHfdyaDeOu/chC
M8KrIQh6sgHP8vYkXkRd8QfiEVLz+eYuRIIj6eRLwF3IjAq89vKbZB5FcEY94I6HEJEpfiKPottG
ipiEYBoFON82YUQUPiY4cDSpjBHjwfSA03FHfr+iemzlQf/mzIVMa1/aC5UiqFNgF+HIQBFFaH36
wYqKe+AOUiP/VTqC/oV8YVzPzkYPrOKik6GTqrgqs6rUmnHK6jWx7lsO53nukHmj1WC9RgdP6W5S
wnTJZ2PWxz9Kz+8snUxY2eUs5soIMkzFcfA7rKFhdtOGCqINcd65QwHRmxYsr174FrHWYLXloO9u
xFIxGEwWcLHIOLlZe5WPFik+GlH1B8bjLWQ3l4X8B/FZypOoRRsgTWZuS3k9bAvjIxpTGpBAcMCF
ayB8rQOUkuMipjckpyuDW4PaGEztUnOE79cIoumt4puY/jNlB8ti9bWQEg0x41ZE7VQqCv2h8LE8
rFYWj1rMw4I8kkiHrgJSQ7Qu2TjCpMuvLctHj9xEChrkvCHVjPWFrNBrDJn5PrV1zJOzCeyljtkI
1ty8nb+iI97Ztm4k/oFnGcpUd0/2y8TtsFj6ikFvaIVsgg42fiBykwMUW0NUDg2zJkwuwZg61O1H
S3VyGh4uS/JF9qroE73HORUc+auYqDFqIbvHc6zUp3BJUx/2qoBZxw2zcOxJZJk8v5mUY17tyQ0D
W5OsOH/3oFfndr+6+3GKXM0icSzjl81/wdDP42FxK8rbhlhf8vJKWgt7C8npZRl5GHiHvVuMPnd7
719zayu53R4IjPRkWM83aPXVenSYkKLtOVNUtGsaj2+SVq/dEZIx0EdyPIMZO+mhfJc/8LkidlG2
sbiQEPmL18VgzebE23wInugBHKgmuaYBay8gTnO9qcK16cvlVauGHaEwATVLCjl6KqlNc7ammA0d
reTa23udNN9KoQeJu2jGSnuNS+x57Eq5Qd+miv5SBWG64mecKHZjQB+75+e9nKxU9HQhahCiIwK0
naTM0X6BbSCq+sB47YFzcsMUGW3/xE+9yVxMb+i4nWwHNtqiIa8upRgwPoS0sfOb8F5+0wap/ElV
PArPKM037rO7ulYAW2jAk3uqc1Yb6xld9ZXPnt4oRLPbG+lyLAcaILjHKzZ2gRSYjTpzN32xnqd8
ykBY6/TlRzIu3rUKU9k2Ql5Jdsw6kEQerhwWevFsJCLLiRiQLqbr/rCsMkFeraHrV5worJT4R7MF
Q+FoKtGHVCmTzDbojupo2wjK0Qb3sPAKOjeqy5ScZLu/bxu1IFm/eEHTNAJC67euvg294B9VztW0
1WKjIRACPh7qgnwEDDFsBl4+6KOk4ff+P1U2r1cvK8sRhhsw1QRekTWYKYGq2p5qk6vcZwoLSjCG
4XtulweSVbnvLxm/INHH6G89k1d0IzzKY4MjbaabmjYXdaT3o6R4N4PGpDuXLjbxJcOThV8db7VA
hJnvnhTMl/EZ4VoQWJ6EqAfQeZwpMSQhO3dV9d2BrjI5OskpcJ5WPF72xW/CSphkvU7c1qNdHhEf
+K2erpFzmMGmH6y2IiAkg90xS2tOUMZrcW28LTc6UPf5EVqAQI6hfvUStKZIVwGOcEvrdv9RFkjf
Uf+sPXIMravnHy15wf/a/FIWyB4qt+ggGP/W5VLZc9idRRD8bfmL5GA4rDvoVRlqj4Z//6S+g72H
IDjjXC2P4HJOFDU37MZwpAa30u9eA8oCrXL2Sq6tNgFfFqeKrSEfLA81x75RcHT6PTgFlK7sVIGl
5JSpQTtAnSZjh8WETA50w2oirEab0uuP/i91M4n1DRabIeNbeaCAEPS2/W0irsFWWaYp+yCn423f
L+a/rq2hau/zP8W8hrmTvpVdCoo0eS4gWMGjRRa2GtZnXsJy8cA62+Vv3Z5CVuameYB9UHh1jLGi
T74M46LdOVMOaIGTIKub/5kSoOxKfwynDigFZSFG7YWk0l4YY3hdZlk38YCLhE/3p1E4y0lfy5R3
Sn+fPs+fZKCXAcxINeJUr0LKWXZ3mYKI7ShYPukZ8ta5JWZ6IJpKjyv0bRJu9/1HOc0dlPl6EMj+
2zBbN6UKbPEbeu0da2PhlnfPkQwlDWzqYJKlFHSi04U/l1jC1uW3k6lpNXyX9zkmlSnGhvCu1iOM
BfdrkP1hFgAlW1/N5w9aIBReup0M7foHmbFII6gLCXQfJQeAdKU+au7T2X5x7wtjvY5UlB9zgE/2
GZ5TyBvYm+D2wnGH49h6fcOVIcZ8HiDfnR18HhIiyGkOTey4OFVHxhBTjIdua3J5k+S+bi4qKd0c
uliScZZpQlPXRtd+ID0T9BWCVV9lTeTU1ZJNepy3qZ8yiAdZ9FHCCAdvM61vqtjJw029XzgOifU5
i5AxQA+iVVGUBuJ+p/e7RfoeoQ/9+7yW3PxTIOOfCFOIWoVIdBPuSL9pHSYduGePzTl5vpBfVTmN
veLBKBWAdK2LAnAfVKNDx4dBYiTpireWTvLyncJuhc/Hz82vwY/fZDSafAn1yhxxRXtB/NeUR1iT
gpFisPIh86FxjauACuiVRhDiiaV5sD8RbIrUfHK+jHeEb2VQibLayyUyxx7VsF6e/IH6C3kFRePr
mAG3vkOHeguYDnu/6/1AxEs/pgbRKo5CVeELX7PcembCS+QHVv1YN8x91W5/cgrJ+F+f9XZPf/wD
5q4AeHwzGCHykFD+utnOXJs0qlKWTNsAXodOMofiw8EI3Jh+M+5Lsb+ZNGTCpFY32lCBQUm979Re
zq1uo6LGOU52laBT4P+R+j6PlM8UJ0RGuAESndAsBxULzEy528yu50g46LRNrG+H0DbXuAXj/lMe
Emui7Oe9CCJJEwjRVF//pG+pwJZwUUGSJVT4geAE1uU2zp+Q77pIHZt+TAKIZ6DA/fbzilS2NhSC
7OP4iOYsajXIruIKmO011YYRc+6BQ49QS8ZJWPSzLqVolrTmugz6BlrdoPQXsW3KVvWWaT2+dF+t
KLvok9gkPiDNuUrbPTUKOGG/p6jlDWNsf/CLAtayHqzZ8CVbAcMSPObLt6pjgXyhsXcJ7sXVcIGI
8JGilY4+/5V7A8wS+ydbp6nNBnWFJ6mYOq+fQ4253ynOv1jCTTrqAQmkI9mB/lI1MCxhaOkLXhYt
Bps87KomVv5KolRmMYNo20Z3SYtlyGcGJgGkSLQFlEayhn8+C3QTmdvgxqzt8qgPTpTwr6oBjGAr
NgMKWE26yJev1seaxldAPmJ0Yk6c/8j4mhQ0a6rxWE/nsLRvjVkRNVOVQoHGprDNQxx2H8PN7L4F
m9DKxNmxmgzFK4jEmWazq2qSX0nzzPiDtbH2F3pS/zG6Wj05Ir1ysVUY5qO7jSs17oHAdRVlSwFq
6gmaGXWprn2vLcIlpkXIclVj3zi5/U/N1Zcbp45XxIrPIKryx8x23un/5debEYAswznbXRfMYH8h
jeVc/B49wcS11ffWJN1ot1X72zlXfReML7VZxe8sLX+myk3emVeOIEmwyglgmIldThxN6L12FH65
lPWpTeViy+kFF1sRH5SrrveE0v4XTBPtZd3CHm32hd7CoCmr7SnODLNOluRwjcUJbOmTtme+zvJ4
dWqHMjf1v2ztbEwKR/vgitaZynD/gIncyZU62p39yCcwH6r/bgQnfvHHxtuKUh2vTTq7wW0+TFXF
UIXmH3woZjlzPhrqPsbroMoEyFxTHIXvWYcK3rysGa+FlfhRVQPpncWEcdh37VlMElnQCvUCuz7O
Uk9B5a62Kjwn4wgTMMBZRB9zcE7krAyYzDqKECPPFPJsAAI6NwZUbequc5xBo2pHZAXMvEaIpxSo
B+x6GyDW5iYIyfnvHWZtLn3B2tqRbel3WBYsQOc/Sxe728RIpVBVucKqGW3XZE+7Wdg0k2mXCGBN
cFTjzGLVzaAS7DBVCp2sScOT6cs9tAFA/C7/LCUmXUAPNZKGIcNs6uMqKpjxopI/u5+lFghRDO1k
NMzVpp6g6RXrWf7h5NaymRnDcnPs1MFIwpmfzDSZSylGsWfeBs4DL257XCsaRl7ndB70Rmi4GA9F
D5UtF6beL6IrOj4HaR0Xp0hZvEo+0DxrjTgWa18T/RMjeWCqxFOS3D/KsDikLbx5XwffnzkUmHpP
JFD5eJOKbBNkhHohgIwgdbvAPSgGjh+qFEUgfj09+dXsmvrktSuA270rS52ADOJwHtHoGTED9CT6
HrCHAB4N5sPsx7GBJGS5CMND2Ob+2q8dS0h7kmJNDPo0ceT2fpvHM5znwziMLgTVtughs7uVkla6
JWuMdcOCmo8AHh/HYKv11Auxfnn3MAy6G4CCva2qNn/jtUs9uAJ+aSw/9/djo7wFtaNOdEUAhvDs
IJpAk/l5J+NaEBkf4cGxlEGw3bfCEK80s8mAamb802oRzEeMBf4xn4XTIGwmflaHPps72hiIlWyz
+q4Z6gcXpsNO+poUsDHPr8DOShVz0i1FA3eWMSBcfWaRbrOicF/ZNYaxyoOlfcWwJTfhVeDmoyk0
OBdw/W7lziGwojhYgKWP0DHE+DYYMx1RO1GaEirQHxuPTyojgpFIGfYENOpgnl6Tr99lsrYPh8QC
dIVOi5Cqg3l6t723uAsE3NX5h0xxk1GAQg8gjWdeYlR5FQm6DRQAsuX1HkIPnX673rj2ULFpDKi6
CW+D8NWF0tsH+Ba0JuKcgxUlILBIHc5jMPH61eMJoe5yrrhcrbhHJFvCoVmFWfu4BuN8T2Qm2z+m
E/yaGUwzk6zqIZ3tP27Z8yCtV/J+LD2wexEAsufc9cQaP6IdTlmx012+uxY6jTQ+Jv3kpWM+QqYl
B+zud+I0wPqvrTlruDudtsFNO+/aGRULs1ohN8vxWG8L4bJF7xM2jqT6t0ngdimHn8jn18xYxPr+
Oad3tHFVE89AKREYvJ/6Bts97iaOVrJFyysPOOcvdJCPwVAWTPMSjzY/G2GkOzU7niteR5fLDaVi
uungaiEUazctkKGipt10Dx2Cuyn8idifRJqP8mZhtRKWMtRSoRFmpaCW/cudaHvhdM8ztK6uUWXn
LY9/sduBNDyqCWzjNA4JvftwCyIx5LLLdGRG+iJ6+b596eyn9PmQOWy8Xlej6E64izA7Enk4eHrN
jB2kyyOdA9kMdl3W59dbJdSQN/A1T+Q9dq0m5FQRF5PWo5F4mjbj5Io2Yph8ZRIBLxtQagFVXdfo
pbjBNR8Xj4dvCeqqQRA3E1TShe8r7w1VhpUYY27c0huAOW5VdaD08axJt3b6vaUu5YuaKE2zbv+h
lz+SwrQen2stRs1fEpAUeCmDpvPu+zeqf47CbTO/oVJIElZHupKgXh8n5oBJAlOhfXhRXqVI3LuQ
V2aODreh0fuWxCjBT0DIGhTpCrRMKErhe69UMSEbj6kS7ZH0lKbpvRZTRBSRcpWJPtdZn/mRqDlt
pi+5Sm0FWxqkBrk43NIb0ugtZYiYzXO3X+caLLLKAdXHYgG96+YmzDfiUIF2pZJu+vvONFAc2pDo
F0gmXdNMw87/xI5HHZQDRbP+cH48e4c2KejxYpF380ZcJU/hVaveP7xZEnbOX5WQHj1lSEO8bSwY
Zm5iqSQCrnpJQ9azoYqh6DwP0Bqg/ZHGnabTaFFWtoDUw7FIGmfzpQSBuaPrSOi1CX0pSJ4nGq1V
o7LeKCvrsou+5jdflNdbt2BxU7pUfYQnoQUuy8evNyQtHrkBg48bvUf9GGeL1DA6vSr9oUR7wIKF
cy6I8oLyYOTHa5phrlXwAIpWlzZ1LnpmNACMMEXSr1+10PGm9ieeypDHyJobJ2OPdokA3M/5RiB5
24w2TFiGPc8gpYceJNLor5xKWUIJfh6mA3lceosiKs+DlFb1Zlj1UTffq9K3/jJ5MT1yOkHd3YMG
8rlBXqfPYs2hIbAGZJ+H/gE7jVuZWf1K3UPEbcyWPRyutbHStbDSzSPG6rlJWw/bmjRMDW/Uk/Co
ZsYOPztt0nS/v6acuuQt27coJlebl6kXNZ+N/rzfOdsTbZAiivtTdzDTmULvlfW94tzXB4Y2kqOZ
PXOEDHMdgcao0GCxNZKw1smRbEH5tFKcuID1UqRGprS6fhWCR5uaB/G4oVBjJ0g9MkpDXY+LrwCP
J+vqIKLoDVunedK/ODVNA+HMzsqIyjFK/SrOLltyMI/uV3sm2BIo158pbqHuH4fMsKbG47eV+AHr
BVrC3TWagSIF51L6hJWrMAqrpnz4GSWffOyR2IMhPSN02xT9K9S32iVh6fmh9uV6QNUeMNcnHG2O
1oNIQ2jG/vjT1zZ8HcRsLNd+DuBf+Yw5fo/EcShvZzVU0uEJbrrBe3YmtlpCOkBq8sYo7Mz6NmTe
iNQjmrLmZ0BCifELVbzzPI9VbnDwBayjOfKmMcfh0GpYyglDNGg/uGZ4WLAIr+B8mWeQfqqeDFSO
mbmaWZAGoROT2NofsUIso65W3KXhTomkaTEoOqh6E5KM6Ze5zWwgRXA+vm0eEfbnjIePD2iJLi2t
8ea0T5WRdAuLzFoxK2tS2GU2H4dPjUUhQeAtOShw8J6mN0Qkehcz6eRY28vzWgYoKnbm36kAnkj8
NRWRIbn07d4/uHLKjCP96MHQSLePvCEQeyA53CeLCcr9kii4/pg+SxcZfHYM/p/CKdix8EFYnMay
yTJOJfxWMGHWj+2z3nu7n/9pVj1k9ww6yrxUve+JO9m17umNXTIpD0FS565Rn4rD1HsDUuGvIg1O
k1uDzKjjI67KCHmMPLO9DCctrU/VwwH9X0AmlPmwQjEKGOv7mZ8Ktiw+rDB355vyml+zuWxgBDP5
xUSxhP6JX82HavYvl6C3OMfGYAGfr6WaFMfjyRU2k+hdelT3UH3M82DMNcLzQy58LC+S7ugjh6Q1
mo1eiGNWPKnub78g6PTntHW3IDstQeA2SztKXZUJ1GgfeACDj307+NyR4rPbN5dWep3FOJODtm2P
fgEnxkwXclIyA7uiy3j9sX/ilL3R+NjqTAY4IxEp5+OQbztU/qW0wtwIz9ErHidwgxGiKD4c1zs8
o5O3F0l4c1Zj7Tzy5Wk/qpPrqwnzFUoVq7dLsFb22hwFxv9r/+KAfPDlM+M0dy9HPvyrIZBuAf7w
Yt3VcCGbvEGRijBcs9hvO/pya1nvIJWv0UlfDGikdoukt4tI3WF4UjPACVrAH0hbgac0JhpByqRF
7UtbLu1XACIZ4JCTCiMKRmw2WFGsqHPridhKLJeEdF/2mjjErTRKRtgesvbGpFyucC5GbLZ7cbqa
FHQDk0k7A6bdxPxN1YLAQaZ4Yv+er6M4xjkL/Ppwt6Hzg/iy73uBqMGV6p1I8a4l3cA34zhAG1ln
XVG7x9R2Bn7vUZ6FRLxvOQKfb6LcGp0BgKYqUGDP6AcqvecS5SxQo2X+iXjLu2GVxR//hqJG1ehj
KZIbzSoV1oesrHfIOgGfUgX79PNPCh5VOiMUkg5u5KpIOVdW7LNl1K5pJITaRYNDN7sBP0SQZtWf
YW5FPq1BQshCdJIDlPuCrpLAT48ryvFIi7E5vuNDUu1jDgzs/rj7SHjKEJaCxSafTKQQ+c+2QO7Q
uPn0cpzmYZoEqsU9JNPUlevDx4FbZ023TMfJg3UHrLyIUCZxFp9jCnkj7DGKhs7AV9xnuF7RVgF7
2wrCYik6N85BBYk0Hda6M0Mj+sqjnW5eBu78ts+9BfMBs7cr1Hu7Cbf7/Z5XPn5PCpcCrNfgCBP5
p5Kuer9aFKsa+j48tm+K8gE/KIhIfhM3kejZ4J2lwBnyHnMIJY1O3m6OvO3jtVyzhnf4M92wCtQK
QJWdNr0O4spfdUfymPNcwnbNO45LjOjoG7oKxdMhMpVTTchPmpwZQiw2VtwZjlW1gskq9DVouXbE
zKXfD53nrCL3dsvXs8qc8tjM6rzpyD3Qveyq9/BsRaXQWcVHTUhnzshqZJe9uZ3Mqyq6HMMxgNLe
vttd62Uck4R6ruUt8dSOYyM7KfuBKi6ImexITvrFzMvL9ihpi3DCsJIFt63CWkM7aHNwbwO6t8JS
49bP4rLrSw5Au8FELJrTXCOx6CEg2OlWVrJGMfnrm5ZC//QpMPmUJ0/nIeLCEKrSA427MPknjU3f
KC1llBnBrXXOy6KaSQHKnmVxhqsEQXuzkF/mo12jObN/XRP7mz6246a1FuUtAuNrlgrLiJwTH7+L
FbJwlDPXt8uITPxg6wy+f+mLDk4mDhtcBRj3KMXlkHIhZUhG6f78AAlx/0+B94Umulf0+sn3oXYT
8jfXDtp1+ZhEMQwJ3zd6sWITo55Wx28qkfvN7b1Wc+LOi/EcpwF/d30FO1yL0WGiOsfMnPF7YxxV
8QJ/XhrCjGL+5JBPC0x5Grpp2wdSWBuhdMn5DtTFZXIiKfWqeLxyiB38DsmIRXQYAFmlPAZVg4t1
YKq7Gr889k+2JapNgNLHOpNhu/qJyRmrFkSJYT+bcXPSUPRYaqZ2RGZmLz05c25JbXqtuaz2i4Th
+qGz5cXRfZPf71BVq2A8llxF4yudlFj6JXspSJue2+YMTOh4wZWCdoNn/z6tNtdyv57SLBe5vwVG
/5+AogJylLDfWzc8Ji9c4vCxOInZ8/RVC2NZyKJEXF/zquyJOAe19RBb8yvwIokXcTxr9sNjKGmN
uomHkxVBaSabKY8yEczmFCkDvxzPVRJaYx68/ELXoJDeLV4/KcH3gjPdyM0Wd0gqqfW/EOW+HPw3
f5eGpgqq+Oe4vfpTWY+zR1UW+EBx88KTFOK3Oeu7gPuRSjYjQJelqmtiloiOeeFOWCGOadgYSXXv
PkcJ46KK7jK7Af849YWWRZ6BEAB7mIcrF+dqn4fSs+NKkILKrHK25mPFJfVnVPJ+I3MUC5Kx2inx
kVpDkPhL7EoAy1MyKl2JdUrVrGfbusydn8Ub23HnZZ/Nx7HJOJiZHHb7mainHFZ/v85eb4lFZtKJ
uUQp7ieZ5yym0ab/alKk++2hbmppHfB24Cpggz/FpIfVyaGipikA/bw/habSmclS1O/JG8MdpTUI
0EaOuwef0v2LYFDmwnz818/PLh4mUXqbOHDIe9gBtw1adygKomgwewVz4PJf5G9m3Ydwl9QTnpeM
5DVSJPoKDthrzUEb46ozjonXBfRWJhlAjYQM7LbBkfwVX5RA9UOnDbb92YmNsV6y33yfk/L3emn9
FHgHiJc9fPj2B0IkpMEs5wkVWKLCpSgXpDpDbvyjIyxBjfThfSQQ38Cei2/EomE/rI9pL2P5nGgH
GQpwgK2eOQPbyChoRacDa4LubhFCIeKSuS34ZjJc+VNcv22r+gMECMyQW3f1GrsruSWvX2qq9y5o
C2chG48U7laFeHstgDcHKRypydB6eLmZgq53HANnpKF4/wpqMNulzBfAcfXwwMNAPqPZkOLP6vmU
j1v8KubGr9ikWsxK0DRuj4lZ/Cfzd15PE7x8Kkkt3ZH69qzznyp6wgO1MU5f9C4fbbu4esUeUFwx
kQTS0D6QpZ79nl9gqVwYyG/8Dax0wn9VKAwbGFXBwWwA42AHJlTJTwqeFLpnbVUmGpYcpPfO5HSV
aIc5ELUs2JrcppMbp1QTirbxXYxTH408fsnb5y/agNYuY9HxDWYIXCjbUQ+et+Zy9bbCd/VY7qVY
VE1xV/KMbpQQpLrvzI45nkjzlSD6KkSU1GfgLWBnfz6IuSfYZdqnHRrMxlP0NYIA5zwTUmwTkefe
BcZr1LHZ7q3RVgXeuMakZ1Jo6DNyjMD+0PQhs28KVxIGQktSACMx3LZVtOakRlarTEXhYl5g+qSJ
YpBcX93CTD02WL9H+foiPI4QK8Wzw8+EWdkOZouzKwluN/GkWI5r4OADSXQTfMerpU48pPul1d6G
jqtELnCCjB8L/gSW89DeYYBt0FNd0+l71+PmLdZSOibXcKxCLd+o4joENCHnoCzl353jk9IAJlNH
gjwmdr08e44tSsu1h4Z/ZJ5jv3toKh6uV+khmPji/clU+mpBwH6n9jZyqkkh2nV2GMWqnfSS6Nwc
iassvy3ZqGOn0cbRQXuUbYXcsB/Ktmo8Kv/X+4mw1bbgtvE9bD+lmZ7kBHQKdsZHw8vNaNGSPsQl
1G9EWB7oLD5vQmM9VCU8TdWQReo+55bbjrkK3Sy7jv3y6agq+T6D0jgxgzYJ0JnQRUzH0d0nHl6v
EZIoiFTq90udEKSsrM0/M1kIO/bli0HYMbtnJr0Sloc17CNZF22UC669DPZzXmkng4r3RLFE3BSP
UHtXMCvHRuTSO4HDgkVuwXkgyIDGqGzQm1NvqwFYIjqsVPSD0LZlKuT0WQch+stiJPHWuefRB+8U
P+kl3XDMdmhZG5zX9RrNY5vdjyNPzyK3RLc1IdCQNkhz8iRIQdy7QfFlzV5reDNGZaaMoL3yhXtI
HzN5fM25dt3uW45kIuUjIrnsFGAXXMjvK3GZR6CLvBlglWjVrbo7jEgcLj7fmFjdRCz0Ciy8o1vq
mHfAztukp5cJWxfjfmfztX6TgfeHC/0ofSy+KM+cEUdZrIdj7NDTjF8VDNNtRt61Tg2ePk7Y5Gdj
Y73Zv9fBdSB9ohZ5kEutwtmP6sf149ifxCMrem6jc30xuyuLD0EpxD0WmsfWYlpmKW90D/8e+5pP
Wajc5SWP1z1BnEYgiEF58e4KvBo8a3NNVxRqKqDe0cvJOlX/pavC+KemMGYSor2dTuI8I2r+jW83
GmEzul4g6qbOJCcT4rEdl3MCEL4cw93V6267thqV1oHwG0AyoUjlccV2O1d5Upov509AnVDQuRv6
ohXDWOIZADzDrcbhWA+09YBb61vZnN67WNDctNiHQBKmXEE8Vn0S6rckQNoGbk9nCHieB04mXRoC
ieMdEUp2RxaSZKjdGf6+bKLo6YLBTFnmDipZs1si8uIwQSEERuhAuq76VRArbQ66yYoF4jg1rm6g
Tbd3uIO/SIiYmavUyKLorWdvqC/JrwssBHOV61Sp0PJh82MIJ3dCktrI5HxTtTFojr3TxzNpp+wr
30N+G/GdLVXX8bnW1uTglMc3nFyKQ9FsZJszOoCXcT6WtyD/PhQgEX7gc7v3QzBUuCbKRwxWXpIf
tyEETsuJ441FTZdJCkgfcPRyDpg31as6FpupueWXYL0btFc36y2UyYd9zz5PiYWGCGKTU3xryQZG
DSsPYnH6Np9P3HA+8KV+PC9UeWfRQORyuTJGR0rWfL5LKUTmP9PLCLJx+Je+1vZxYLOBoZq9rLgF
uCcRC+DOGJbba/1MsXsw+mu/wudZqi6zrOAZXdrHHbqiU5qcQa0YGD0mQPoysI0mCoXhvoJKH3tt
kILiLYTfRlWgw3KFxeNOgwb6/0pnMMYTsv95q0m2tvD4krS8UoUsCBGfXbaRSSxfn+D2N14nYXd2
VyylFNPoF5b9w/2fdvpDSHSsCQ6+dvluefiGFXYo/fmIfRB91oBcX6c5oDWtg0TTaaTlPX9lIP9M
BqWNWAE0dma8WtZJvZw7U+tvxSMOriom2KSbYP2I8XAo2GTRpa4F8kJJWYo41KnGQ5+D/qmD3rQ3
t7YzAoIQOeZs/cs/jlL6xj6lmmRYGk1pulHYz3xFciXO3sJ3Kn5RKeQQ3/QqRph29MrvUgzcKJDz
lU6YmlpMPnhJjEL5XQnALXmHLuvX+1MTIAfpKqXBO9K9SqDM+FE5AT0TPT6gLzNwlm2foh4aEacy
opeRb6JYT60UkxfdBYqTIMuelnSVS+xGWnWe3kNHv4dechZqqdRaNULRPApNximGVUlp+AcbLItx
PPurbtDRXNifnTvg+OerCFGr/oADkQm/UvigMgMUj+leRt7+P+jFUTJhvjrZg7+JDYh6L9n1F49i
QGHZwoHNCDtTJoabbknok3JxNs15m5WQLA/LVQYCduTDkfDEtWYwbBaJ0Z+TReC8NfWS+yC39DU7
ht8DuugITpHaGqe05Gyz56td8hBOpjsjuGdZ/958AnBtJ6DAOJtewxotuRW7632M8tt6hQfXJJlY
Ju0jHYidqc8A+j8g/n0F3rOQite43ESga3OffZ0/PA3bDXwSgofMK7C7aFmAZYw01ySH2+7ljjiE
NVX+mc/QJjPKpiuzuVsf/x9CAxyQ1SkcULJLETN/VvA66c/HojL6ct7ibngqQj5/W6gfdxwxQMMA
whx7oBI9OtAgYg55PwADqiKmGL4EnqikBveWQx3V77T1Dt8L1/Tv1vN75yuinhjWFVG/FoosdRFF
6ouzn/4ZrLeDxQ8SjSCaGP+wRPZaFFUQFOElb6E8YlXECrnnP8qqk9VYp38xEB4LKybabeyknM+e
6HxKp/UwfZGbtCAH6fa+MztrG/YBReyhuiAsfui/7t2JcgZOQ7DMg9D1SXPBjJ04t3ph4UXfoEkJ
jHGrj+1ACMHG08VDjSuwA1w/07I8rEXKjEaCrt2Y02NnDWZkDwqjYM6xH5zhXufpgBlY4m2Dysmg
PSEV2azn9ttOxlEwMgMMS5fYY71NcwUgcwLVxag5yuwjR1R5wS0BR73Ca+ol6iHpu4TYheMu2Twx
vGRLbpV/mkhBh034Pv1wTgrQP5TTHuZlcfKbS1yFCeCVBzFoQ97RhU01AbWxSUHt1hDXlS4ZBxQm
WnmDVOn2h6f0Y1Sh+vSpB3SO1ygSaIeJ2G6LUC9+V0+jXPOw09UJaeIVhJeT0fSxRMsJEhN60Pzo
SnDgoXmFdFPr/AQmn1/YWmo0bZacNAEsVAsFH30o3wjqmzz8IIbepFhYPy5R7FwnhpA/gl1b4qck
feEEFvsMHNF0anxPDWujgTAOrRtAumAGmMXxhRd8meGIBqI+4JOQeb0o4h8QwIDYCyIL9A1CdZRn
FlyRpPcCRA9lrgxDKS9BAs6ImQVL/AX3Yt/SqamAmEZgWQZIVb5wGwN2ghKwQOe5G2wF1wx2m1xY
a/3LtsojAJgwSXKib+d7WMQMZ1Hvzqo3/DH4Fe+sq3QZBJJmIiU2GCzmmDP/ct+4/LBywikGL/iD
SiS8VIJ5dpEYonACbcyduCW74rOVsu/valj6HeGAHcIjFXkjpk9CAQHb5aA6BqBcMOP0X9JB8+j1
VK+O/9mT4HV6BSQ6W8yKNcAmRM6QyGrwJKV82C8Vw8OLRUTZZjFopYOe6gw/GO676IX8372CHvds
xWD6UFVk0LpentkWfWC1T3CsxMFMi1C41qKZxlmYD6lFOYk76IpOx1z4bygz3t9z3raw6SvvAyeR
/7WEsMO7FjL6sDS5aiVOGiNxxcsqAhpzq81FZvuVletZgjYIL9VBy8v52BRw5oZR4aaj2FA61ufk
o2wUH6jmL7+pRNO5UxTeu2hyMcUDndannv3zG1j6yhU0Q8CICyx0XSpfJ08/HND2nH3NmcbSWbpQ
86vo5CReqywj5PqBGgKOF8VUGWtxrOJBqYAxNERhAi7Me2/FZFNwS/fwG+1WnbRnTNHV1SHacL0q
Vk9Knbt05qGq2giulDzK6DndcZWzzgS5P1cyexYBQgXVox6snaufQ/Irh0J5LnYCQBqiv6A87sSO
BO4lKDbwunSRG7pOB2DZonSA4v0bhSTdSuQaxGRqde7yiexz/KtJk+NiPbeuk/LqN+42j2pFjMjf
6i/wlRdkHk79hzsIzyPD79wGAv/8MD7Ik4pIypsw5yUkAActX8khmz4lsxvS3x754MR01q/pRwaI
6ujm2sx36RhUJH1r3cb+YVVsG0Qz484uZsZxUhHZTT866HlWV+Kc8TfxyvKvndd9QXPQFcR4oMKA
Ek3978DKgDvD0gN4UuBgYT7OpsgvgpuRRY5oOFl+WWzTy9jtrASLdeaOeU9nSM0kezvG5HkzRmhm
X+B71hRdHlUHl2dEAcv6HJ8eKuigrY7ILKzs75gn3pTmv+OLi+D0sQwvft9U7cNiQWvULLix0x7f
OfSx8k6jM7GsbEO0iKK4jYzUJuSlFvcDIaXRXtpWBqj0xYyjLa282q7IGRlVAN+ijPqczoZCLRa9
bePVpLYwAusTapBpDrbn2KRbzkT9VYhHN159SsQa8Gv3RXDBBPdwRxQGic8t4amU4bHywPiQKlBT
jrG2wCBJkhMrtkBymyeH5XzCNFW9/qN9SeX2pZQ/KaaHLC23TJQcyG+d6jAYp8zRDv2h37NWU0/+
9FxpcZl9zOF31QjO4fSdQlpcPvs+9fAoCBDC0gOKjqP/pAhbVOfLAdZVHfdmlt0DTJQH4kJ5AhbN
F+PHf1VYWv9eWXDU3PAtuwKLpdXOfH9rN8msYSfzYky0EEwkP+rtsLvGEtgjVHltltXN11Fjsvog
brwsm+jV/eDClnJoUrnHQIaWxQ3bSn5ZQaTCz/U2pPw8XXz1BWnFo5Ze+D5rYNEbjWUleVfiQXH1
7ltVDG4uO647X8g5KfTVd8febiqma7Tq03zHJtIBQyBfEVcWUrVrX3Vji5HmA1ph0NspxUcfcWCW
Ez6eKCeuyems2MeUY2Fvizo+FARl7G6A6/ZgSQzVGIdKYmxS21ms3YZzfz446u1VYWIPvSRAgQTM
rKF9PpZh4QUCqkFvLX7WP+SAuOKmsKvh0CxpPmNNqz/hqtSb24b5XO9gZgHgBW8JfKoMzM2nO7cc
Wtlyiiz38a4PTj2Nq2cookZo/PAF0ByRTShi5x3xer5ab64ky6sU1YzBHtywTxyL0dJI7AsplYWT
qz2vcA2UeLfnwkR5NtqVJ0Im7AjTHoxx1OwA3MBSilO+49F8OZHicb1gl19d63T+F2n6/KTeInR3
d1DDWapxj691u0Vk80E9SC4KNw1tAKrpb2d8nVUPhvhzdYvxVLk/aHSKHmFu/oC1JO/aljx0tvr+
tuNRe7duLDcT9A0EQhsTGIRlHopZ7yeplUVJeYWrXIlL2i67k798RibZR05IoxWEtL3gYecut8g8
FzP+pStSxt41JeQr7QUPe6itENJB9I2bYxUcX+xb8bF6ulJHTCyhnzJZuSRSrR7KqOSQuZx4ICaD
KD4lodBaRJXRYsgh+KpgN9dkOVmx0ts4oVmcTAeV4vwco+R8kBTO1i7H/C4KNPbIDWXh4qOZkCum
bD27NIeoseYcBdFgpbkTzLuapGC3Dhl/XiVpdKiubSwCCXw+IZMoGJYNGlcgVZJI/S6gLa5Lb+cQ
SXhD4J8LhtBGR+fdtcFVXvaz7RZIEQRGFfT/BULQy4QxWnDle94RySsCGVoRkN/urhH27sbGjWS+
h9+umJ2YgYDxQ60C7xoZDz/zX0iN340y1KxUrWvKI7BkDz5clSH5enaNx8jjeSCa+HaDkRpWEJ9N
k/j5TpBIx54Q14oWaQMj03x+vNhlMGM16hSAIRMBcHVyXAvV2JmN/km8VnceYPxiFiTjoIg8KMbH
DKkxqABLY7fst6V8tAajOnzJ2zFyMlhVOnkqe01jak2WYsj3GhjebNTSAY9wca52BDYt8sWfQJbY
KD5mr1m5hINfF4BdA3v4WwcAUbsT4zba0Fe3GUFvh9RWglkc0AnNT8RuFDcSVEY6GuNhU6GKVA/P
17PpZ1WJy/hqnYPrgmfmQfnw3asqb0O3sEtEtZ3elT/y0OgdUN0IaBuFUiSAsd4MHzBP/TV2G4xh
4i+9gLkP6kvfBIwongz0X4it8NtiH9yLHZ6ng1XF2J2TNYoZkD4iICUQha4VB2v4fy6ADnbpzY+f
LIrwgpktziEahXzUV8n4CPx4OVmOKvLPAUf+65D+nYDMwDp0u3qVHeffkAc8JcyHRLa2WA42Fm7h
saO1RfB90QGeBSLcKl3rPvNuAEWkAw3pbn7CfBT4xAs9YLlfAQ4bRMXA7t3TlIZnHL7FwnC1HtQs
ebWfb2aped41xxAd2T6qBzqTzAe6259GIH8aIAOsSSxyyA/RU3ZdkkBWameV6mdHNgcXm9WzaSUt
tR4HZ6DwxlcZsUW2Mh9/332qT3yYpHYmnJOxEL1SlCGV0s5hfRrk0BVgLXiBrqPxgjfuNYq3wkva
8vwrW2VkVbrhNTgX9SKLeiF5mEAIgU7jOen9maVJQHUSxOO0b35cpb2A7DO7QaVNksBOYuqIX3f7
K2en2dt/Gy47aJ+hnTlSBWJbCDevXO/lqp3Lu2JSdemq29JZz3aq/FUtVfypSGyadPEP/tLzWATC
PIQkUNO1nc49Oo0ltlPJWoeY0tuCgb54M6ymbejNV82M9TfWUI68Fdxuqm9WlSZpSKqsqtNTpS+z
5Kfa1pHLdr80Yo4QykrOSHiU/u/83tp3ql0SvNA7R4YxrMeyO/fMTsboBr2dka1qqk2h5WBCOuW8
j1nx/Ow34ZYpJTQz6Vr3IKX74bgSRq7Lqx+vLIdXf60tIacvAeLMuuy0AoBNe3gDNGg5n6xJkn6y
zM3dHmLXMy5irX77ic8nOVJWsYtUjtjzxd652CvfSezW3f6a+yfXBmy6cWk8gJ+MAAzSPa5weiyN
uX/e3o23mC8ZVBTCIsbCydBzS9X/7hiTkWOkz+rKeNPzS9i0Ya0X/t2k7N5FNQNJ0GElWn2iG1QD
VLrOan+3SJFlGrZf4EA09zR1F5r0GQpAxlYhOaZ63oNTQ4FFMKIhNUq7DcsR9FI6H1SEX5fhXr4r
hR76w0CTwus1jzSB+9Q+sVfFXN7xOhpDVq2aYAM2t27x9seMDsCk844qjBrf6/gCg2ohNk7HYi6x
aySqNQBYpYpabK+kwdPysbrenuFxDtqIMfkWR6Lj81BGULr2aCd3BPWWtRC9jFR1kP74mCu/BKzq
CrcP8+S8X6bH6QfmpyX7BlwOAFcL1eeBpMYdNBsI3iSvrtvG/+Vi0wsrxzOKOJg2euqO/QvOob+K
v2aM1ZPNI9+9FYllVgK2LzxLxqtagzkchNgPbejURhhId55jJrWK2RhreCQvZQpqffwPpjOslU//
jrtEh9+WV3Qt7i7dvEa4soPkQgAhK5DE5bWW3U7EV6iTvk55KLTSr7rbFrPleTWMxkTiFN0mofoD
VMCoopMBmGm+kj/AoNNZSEm4cl/7T0bv0fmXkuH4QAdSB6/39X5PfvhZfmJSMnpkpzfJBGkzlF4s
RGQojNzyYqPrWEO0MB3omPhIBuPSvOKQ4is80bDqvrcmz4M1pUedEwAlI84E/OTvm5duQs9kDd0L
6YrbDHB8Vzlb3tFexHToGddGtLqqXEHFVUUbDGeNRWi9jxUwGyUMnX047zuzexCLJu7u0U8tb2Xw
wDSNUFFz5ZM1GSKWN2yF7PBZ+qpsuM3lN2FfVO9laPHIPTMxq6DiQk0M6szg6Y8JNklzFwhdlbz/
tWQTApbLmpHGaShNoYXNWD8iVxy78QE8BkOc0IWuupKw7PZtRyBC8Jl2v62lMgbVnuV8ToLclzPZ
ERX9o9/Uq2WqXH6GQAbjJH4K3CRdCa2Vh8PJGULsYhoWjISVWG5N/epq9+pFHVnljnNsa/ZAmkn5
pHlrlzZd0WgpHxuqOQitwYbJqDjFx+7e9t++Bcc3dono/6GbECkeLT4QHkJHYtoVZcCRZqN+U3Zn
oQ6f2zS1h9lFAn07e/uaKf2pIAypvWquppJ39vTdu5xpGqzSahWbVXvvGFfDkbkNiCShgcgzR61d
s7czSGl1rgT9MiXoYEbOQgeI3rKfy5elEGHcGDxso2MSz6M7crwisCxG7fTkcttquCharqRz+UXT
d6iTckf53Emk4VywK0YZiUeLze6cmrFVweVznl+GqRh/Le0Q3nHqTh6HpHDiYVmzYrA3dyFy81Te
w/W5e115QUW1UJJz3rZHz/arsanzXvXGRw5uQEnkJ1EMKxsl+Gjqnf4eOnv7ImmOz+HwMgiwSB5/
NIcQPADv5VV4zy1ATUvDwSnAHVCnu9pUa+Dqu696toc0UhKtdgYGeyY9ZCv3wa6PWX4gpeh8m/p0
8PwfP22yK1Tp7SYM8xSs+A3M8oJZ66us24R0Ltl+4PXhPm9tC0wHpd7v/S7GADD3FR9dO1Mtixvy
Veo4nlsMeEkx4yIQIeog37Sz4cLofF43ef7716YlGyVlhcuLtmt9oBmDhKUWjq1Kw2Rov5PXNtax
FfhT5PVt8c/NdGdBwYLmlEFLPtOX2RFiAx+O6mGdMf9NKLXJjTbTH+RK3N4hAu33w/4sGMgJ/dnH
mMOTyns8WuCCG8NzCXL1QuGd95pJi5VU1osF2Xkam3SKBWf/aoVXPA9qUQ+ShE2LJE5WZD4QDgL6
SGeWCtVxTnWOI/XiZfIah/n2qzO24fDqwzaJfkzKDHl8860/qJ8UmdGXeYz096XUyHK+9l0ZuFtA
6uNGnY3/iy3Y79nqbwwylLXDYghZ/9yv9Ns3ighFgk37aPnYG13ez9QV1tTcoz3l4bnACilWep2l
m4SPQm+7iLKA8lMakXTRDT122ig3r7TQQ+eiW89xHpTUtZwHxN5iVA6i/tkeaIH4p28G/hm8L5c9
qna6blxMOxxO1LjX/Ayhojujq3Tlefxn7+jztfWkv/Bb44HlBmxSFlkG2fSUSjsV0LDixzzlPyZB
0LDEFdjfVNweP4sTccqnQyhZfOwLA3DTJZI84EWylSXqZ1AZlIIsqXKhC1sPdz79e//lhvHimuKc
tRSDQi6cG3bYBL6AbnMhiC1bQUxmOHieWA8zo346lz8RbP/SwuePB0L0EYGx1McgalS1LsBIlAOA
HIS4k1eCrMRh6uermrdEsuGZeVRQAfizqY3pbUVcL8u8l0ccuom7UBPBaKibM244SN5Ik1preYwR
fbvqB6OW8AG6frzG+Gsc9MS1owLv7nJY0GSyBY0R2zcj6pFt3j6G7W4ggRDbjFGYnpNO7hy9ETJA
lV48apsyrgEG190HvOgCM0y9I5WvliRJMzEWmSSvZ39C+4fWRTT6V1ZpTzx/WmHcgU/T23rNK+il
0WYDuaodxevuxHG+O+bVp4/ZQOoc/uJOFy+Xgqv3vJ7DScup71970Oe6wVkPGqzKJlJXxJBk8Z8+
Y82OcOFDQEwH8e2Wp7ycq9Sifm+3roqKFziY21Ki7WcXkZfR7MGJ+juCYB15KyQfI5MFXD/iODS2
WSFjj7KT8f1nYsnMRdW00ryP6WcL63E9gIING9vnHLpxkH5Nnsza3rptxrr9FSPzNyIuM2x413rN
xHxrT8GMJvNix//CI7SQoKDDh0Cs7rBWNnebXnoe7VrTItYl614ovMLXhS/QjmLClEH1HHklBbj/
M3hf9STULZgjnzQJDHbKdKuNUuNQdeed7pTiWzSznrcMtJCThVUOQ8SKucTCZJTetKv0+mZtPmrK
7WBACnoOvlvcm54np6kjsrTj/xYhaf7BDFeVCj/CA9A+6gdrx2SYwjToSHRDuQYaWFoCo654cxU3
xs3wCrabRl0lYMG3JbXXBqDlWuBkFH9wzneW9ZJ2QMwFWj8gGXhCYogzRUF9WbnP45Ilvq7o/qsh
MHXRIRE/qf8wWA0hMk6XfTdrzAMTpevJCvVk6twm703rU+RS3QTee4M4Pzrg2QqZLzk1KrYcPZGs
FH7E6zx+vFOj/GYC594/zaH97pZikkWZidyvhantax1oGezc3T5VM7BY8j5uwI4qqegL5T2lB5IU
XNt49FlMuDdExPe+LuYhVgav+tjtIrw64OHaEvvkqF+Yh9umq+sNtY6xTGfJV+XMm7izHn/mVlpp
PJsJOybjwWNF8aYjQtiyH1LLXePRmJMKh/6KrkWmbhbr4H1T9zfHsd9YrbQOpQ9o8A9VMUUReUg3
i65QWvWaoI8y6xtsg1GFBcnx4eLtKFY//ijAAp6EqaufGFEW2Gec5ld+G5R24jm5XYE04Iro8hpD
aqDqv6bfOsJUPUOkHedpcKShcDZ33ol2NX24A0wGbdJdZYnhYZLYBBH6gX35Q3kdBuYRsljCSQey
GlZw/w/0O9ln+y+8AFM2A840tJErLYwwLqSrX897dsnafVm3auz/eGrvMAw6mA2LQdh2VrYjfLrN
gImev5u8viH9qNIeJPJL3wJ4g78acRApVher6qEg8PTs/j/AoUWezcKuX/1QsuEFTEtcAqIQ4Ogl
XlO0uZSmFhw7ORI/Oa2YwiJA644RBxznlcQlEjKIwrBVWf0yJuRjJU8AL2Iv5XvBs+aPbP3KJYBJ
FUIMohZTvtfcrfBv1ntNm/5yo+zog7CzKsfkjLWcHu31BNVuvhaK2Dm1KiVtGqBVeG3gqGTc2PaL
v8BfUgvwnHk0DboHsi10w9LM+BxXIGrLBSXHNOOln0ri3rqm7Oa34wyy3Gpn5sqR/ID0qpf/p0v+
B910Tw10HbhoUkB22vm1+Q6pJ5aUWW4YAaDFKigER6Tr+okRy2Y8YBygTQ4s7ZD6rQEB/4bEnz21
rhx3bMIfL3536faBwwSqq7Bm4DecNZZ/7H3d7iga3Z4SKMjGfm/pKCK2wWTEnYT2QgZixY7yxVsQ
NOmqjbQJUpR6rTwkQwilFCc+WvBzptoozaZPjZryuuE5C0AJsBqYFUMwFEhWqg2Yr9k/t/5uvX+z
087Ns4qee8H0RLcdgany8e0LYEkGT0H1AbWaxj8uyqMxS6JTan/AAQrAyJan7IhefNAOrGVwAh2I
LwFFEXmwWhU10QajO3IhiB5YWwzWqkbO2ejHjDp/pXRVT4vGDRGR+/FzDrj+/W62JNcfKTuvekQI
xD3OO38SkZ/yNkD9QNeLJFadYTbP3H9E2vzFnRbKo3lrU9sCf5cA25zNQfZeP89hxGLx+MyPfmj4
H415yML4QixGfuDufLeciEoHF2vGAUHZJ3qCYXaJP3C31Mn+fdFcDdI09VW2DCfEga2zwSsPloF0
a8CNHqRBvhbygZdXdu2Xw+XKxnte/sP3svHrKjck5DJBlq9PDEh7xMwgrq/ixsnQaAoj5vX9mdik
vKcDYZdp+YeHoYDJBHfPJG3W6Z8+vRbMFZHDcvlRnRgJkMG1jwCXOeXB9D+63xIxZz8gEA0TXM0k
rsX/dP3Aoybn3AE9nxhTOqehKpQ+fvpadBAxfAaLj0PiGjhSgfwMo2G0NoTvTy+sHwcy4f49YNV9
nbwf3yX3zIQ4XbiqaKMdq9zVVFV7sbxAUeoNAQea3ZmkQ1A3Yz+zakh0fQAw6hokXHoA3HfTWCEm
uVnGLVZ5IMh4SIkF9W105xjsARG2JiCkx1weKTDqeSQ56mHe+++ig/QJHWg+HI0GG1cakYeBdajZ
oJfT/H/hNsXRbvhKZ1BrbxoGNpncfRlSmP2OqzKiwqkWyo1TqMq2+nqc3oJktfR31Gu/hoTtOuJ1
nKY5hO3ho90BNKwn9kUDaEGx9fZJTtmCImJXbm7lszvkTU6R2rQmC01y1TeIHbX3XU/qRSbbDbE8
/0IPapL9/7PRX/JhGDdBRswSejyKc8wjeaMehI2SaKWfkhIWiv+ozqn9N0c+e9BpyeWMTv7Veex8
ETk58iauA6KjXAP7zrf1lgxkt+gxvvg57C7FEo0Qg0EScgmSoItjD93FnWCIOtWTgJX2MCDIz+L7
Y/ly0r7ZN72euMlp7MTGmgsfam5HpHU12TXGM4L2k3xdaL7X+JhQcBFil6WfUn6D3AOB9dd/EhDV
JZnU3Z80NfVbo9a7B0rsBZMVb3u6wNb6hwsHrH8N3P28PjWxNcHH4w6J7ToDls0nQ7+aRR4vdJo0
l/BVWYHayYAtzQ1VzzRK7Gasr2+TH+/LgPNTyhkdGjJYObZuxLwC2Jh2pGHegHyOklbuwlOhkk43
+6s8X0u98ho92IJG6h9T8uiJwSe9kJxXG6TqkTUxUCPbzI7cXSBQeiqGn5u6qS7MoWNTcas7qcSl
u53XAdD0j9evC/UTaCpt0gAxBmzeoNayFBshTqQZdJpacrktR4yiqduPAEfZsFQwirq0DgDnJQ2U
Obn+hlCiWOn4uc9wLNNWbLy1Ba6ZVDD11wjABg8jdxUhHfhIxPJo4F9+ur6dvUOA8lfktMllW6RK
QxM7BJe/+H4Uo9Y6ttYrewYK1a0USAd+IXS1IUhE+9K38evBoE+h6/Nd9uAvXYOPE7Eh58IEt5t7
rSRCosSBm5VCH+cPtTAlbaJyIyPUoMDpoT6zvbDO857CzdvAC3JPCwGku/c6Z0U4wOYSRLOQQgd6
PxNf+VQkpvIMTZfrgs5qMTzkDfcfGrEqp794ET2VZezun65R9XDXZSPaeHfhLblWezu7Y6XZH8Ot
FFjGwk+03klVBJ6ORsraiaJTMz01aMaiNormBoODJVSh4mnFsobNalW7aoVCZWurxViw/dtgUyE+
4zimu/sSctCNo9I3f9v+sWeuZEs+9MD67Lyb2Q7R8qf2/pPCSYY7v9H19gbc08vj3OTi3WKNsDPe
4MsAOhWFinDqtUAApO9R/piyB1lpwhxakX0qEKvRpf+QK/OAmcn6iDOkvTRFVN+Y6MnYn2ViiEeg
hi1uWWtOgZayHBNyEZjVjkk9zzNzZpL1l18jIG+zfE7rNVfUQQO0nQUMsvIpX9h7mGOpW6S2zoAk
DxPuJ6+gCcNZ612ezFhYsfp+LqJ6pQzTdq1V3PovwfTvPqsd0Ak1ejs/hTnaQpjqSq4N/RYdoQoN
elO1o4+SyhvtZfI6rqwPwJ247Fd4EMDaJORFSDOca9eMbZIpzlElEqVK1ZuCzMj4ywDZ0Wu3Q6Cc
QOb5Am1YHU9/t5ePUH47Z5fz/3WAnfE6s49jArZl55ac58vO9gvt/7to5dwmD3LrBU2LAKpNOaIX
ci+RPH+oVJN2l+K1TgyTthylSdB4pd3Rsn+u0hjp57yLBt0ZLihpCSRIjjCar48KBNV+JkMnVgwE
EvwieVoKdAFxaS7X2w3ZA4A9B02163tr8ZhYkC94tL9krKckJOkBJ5Nr0eyryTV2PVE3Ngopk1QP
rDS5Tix9tmR8FR5XhA+lbgn+52GTPfS8TDEdzdUjJXybc3UlGg70E9tX9KIb4Xq6dsQ2ozLoCBoJ
HgASUUiyatThVFXPbRmTSoXjD46n7Zfx5wdFuleROmAoiWGdrc29VJi+eU2k+gyyV+SL5F//iNAg
Jrsg7jz0TSYnGV1mf3l2m1d0dOP/GK7NIsqJL+z1XbK0ovanR+6odmuplwmb1MWUktdkDMHEfeC8
otXOVovCqcSd/rLQjuKLEIEL1mrDcu5Ay5L67nUVfXNf2cPSmBmTwhgAvWlcF0mhRVod7zEY0QDz
CacOltvWx+e5mEH9PfNvbGpob7C+zQ+zlyCFBHvcTsruSHwYJ5s1yxKGtF5+EHcQvSOTQgrIOE4d
4572kiY+7+Wz4bpMN0LEJVfstGK5q0J+SRALnL2MshF5anf2Mp9cUZNYk+i6FjUA84ZzrqVH+9gS
AZsYbrV7XlkrgW9TF6vf3K6FMT7TcbJJ53sVRqdz+LnGrnfzrfsynytZ5aG7Ly5+sFj7TnTghwMx
zLZtRRtD1Lhy2TfuJkuWgFIqoQjcN6rP3AWrGmqAjuuNE3+nNfrYP7KPfR5x52up/mcrphBOecgY
xoHn/Db8oU7IQgrxX1mFj55AYx6yb6PAJTKccj/Zq6hQ8HVEIsFaoq2D66M7VBL3U+wAL2+kORuA
bZQdmvqnV2g4Q8lqj+ylBGQx8W23thxAnA2/pqqQF24V/kLRyvvcs/R4+l/aFBOIN9Ygf6g5dWwf
gZUiS2gYFE31fXZD/RGt8ChzQ08S6060U36qw6jXgbCnECrQWl+Muh9OsoWERVWO4w49N3+knvOX
GSxculLaTWXEUqiHOmPuK65sNY56z01WbtQQWcRDHMqvtYbNctt0NSp7lgb8YlmAEfdnnzs4ImiC
dO71cSVtpCZdC13w9SWxbrl8pKIAz5xA4EQdmiQYiSYydK5NkcXVKok2INJIrv3GVH/Tv77O9dJH
TkvztLCWElPqTGosLGSM4hY/+4r4O72i0oAI8mDYF/Y62YY9YX2dqTZ5Uc4LFyjiqmPFPKStXeTg
POmlPy9f+Rag5eKB6DZYJRCpwZmpWMQrYfEb3/BK+ztXWIUa//YOQuLY6suH9g+/7ctQXDD9h+XQ
Ki6sRpFwVxHy5szAqfS2fWXmZA7BC5erHF1sGlpJO1gSbgJ2XIBDez1Vtw8Xqx+KiI6Iy+7v9xRg
hqdoqEpxZpNbXPFbEGq8aBbdvB4U6LIu/ANnDI3JEozvqFdr5cmYl+RA7fJ0OUZNvIvb7sQgBkWa
JxKXq+vfyZGLpt745ftaLQc5nxqTYcOS6oWgT4Bge4tqpnaB7omqLF75LqoBbqNb3yRk/cJiFU1B
rO2Zsz5OkgQYZPKamoADhNNBCldd2uWWCJ/e2LuXb8YueNURH2QNyOa2q1eZqThpduEWgIGhqWyQ
4Hans4szeO1VGN0Z9cFTYhwixGDnQl1ugXzGdq3eC0pCdOb32MAd2MmMhs3czYqhWBRbD5mbWi10
CZk/EA59UYxpOZk1KUUussOgHsEx6ZSR1MR3RI4tb9bDUSoj8oSR2n4gQD6sGkUBF1yoAqDa9aiE
Zrzyy61LkupHEroWTt7fYnzMFRSfq91Rbw9gILFgEPYJ1jLXnfLhInRafI2u2bMDADikxegcsDcR
dKKn+RPHSo0iA7Gu0cibNdWg8/Xn2ysnlxLVu2Bo3sapTLfEKg6SvoMOelAKPq0Cg4K7Z7xIqArG
4J0P7OTUHUGhhyqdzif7oko9wG6mbIKauscNCgC3p57iMHvcrLOcBICWRZn7uT5jyXBhffQj4GvE
JQhE7qUY9JxpcVOF1X9cVg0yHp4U3+kB3U51gccZoWQNkhxxOX4HSHwtcNJ1UxT7gUR/olZVruVS
2kfSf+C1g/F/hEpLIWtYHNNV0P2MIU9+6y4MsCt7xu5ccOTXz6P9t+bLxRSoCrbIotCONX7vlbpG
mOLI2LROkRTN4ko2bBthGZRr3SCNtTHRzXt1R4xJ2IJtH4xZE4dd3b2iLVhmo2kpaXnTBoJfoiLk
mEqI4Ri4yV0/Ysknn8GG0mmjaJRjpNONKkVvU1R+8199I2f5XqZDD+YnffLefYt6wT2uAOs51Elj
kP3bzKnymd5KgZ06JvE67Lo+evNfwT2ByeF9/OULsB1P/MlBS12tONOn0ebySUE8eiYFsBDhrcQp
bl7CHLwQrDK7fgMshG/aZmZLjlQjVbNd/SsRzGosnSJv88NbLEAe2MP5oROz+O+4MFbZ4VWuxLIr
pO4PBP8UkV9mN423RWx2m/ji60FOx6sgI/LSiyIxcwEeDbn2v45xpnUlMHMwaQM5EacEsXd67hzz
s8SSNA6RLQb8TX6/mRLYJPJb0uKsLLOS66r9566gyWGD9y3fogzUf8CWO1PZ0x6OdZfHYEGBWLQ+
ygp3tSiQiA3v5ArslCSvM9hLdM7o70Veg9hQuWKik1Wk9ykKwXrPSgbo+NNrmMoJ6tkmrJrIC1Gr
07OdkWNPXJeIN6xCc1Jj2c2WhRrooBOfQMf26rPY/i5UrCQRxpv9hFcH1nc6Huj5Z+NmQdjZdOv1
tu3b0kcV6byjEGdDAT4JQXjJ171fYVqBAvmKohgCdpnpfbrpLvVpvcKh3I7Yvxu/DZ2X43H8XEaE
wiqf0ajwgJeVSlZ0XA1rtt7Cgj4Qa7zMfpdSG+cO/2AFQXP/S34DFJTWJAqqOOwUnHufmbPHylwr
aj86OpdT0KRRgbQTZShERgj/xR/z63wsqgVMqThqu9GbLkRMfPfMhtfYv3IIS68+R8pe7p1AVbAR
LkuDCMdnBq2HyWJwIPjgvD6fPIOXrRnzw6cwrs4CvJjYf63P0qgMxdtFwwTkBc68GwPECe4RleV1
8J+Yi/TT3c+t/gar2boiDeJc5Eo6KJ6EPfVTQaKcNqlFyX1OmGBuZBWsINKszMRFm67npiXJVdY1
u4ENbJbsMbfRJ5R+ztSCs/eN0gLDIG9HvDc78f5c/BJoZSt4WRAukPThj1trxV2S6PCUAYEAdRu3
/5Hy6mzEfChUN17XvcTsi//Z3bGPFHlUBweXjtNqXDNO47ytIE8Ont5XiaiVJ2G8++ekr7XuMXsV
SnTeMfVJE/hrRGpzW3sG5r1OlihknoON5G91yFOsmccFm198jyUpaZyrCHxKOrVXIsNNXgQcphTt
aoRaIw6WyOLwIElBDQZKd49GYYN+/Ycvlm8tngwC3sKV7cFCVeZVQYZlHUIvIWAlkcyom8EsS8Xz
GUS38Maq3q3/Q/wAwD/EZ9Os08+055wMzlO0b4Du8uKnubU1FM7ND9eGFLaEgg+AuAr2Zd/0TYgP
MCK1H81XDO+wN8id4ysQyPrV40yw3RUym4zpvmzUmjVA6QKF+iou+8/5Gk8hQgQyKbHPEs0vdd7L
jmjASmuZ1nHdkZ2toe/AQt9tfezfSni0WGNIfZ8kuhPnkWwp15XGgU0iMm1SX9eZ3FKY35kHxLAG
avDUbMukCDvFJNmvltHkVjCQF2kItOIvpGuFihNuCyt8IpUb+USg0qXkUM5yWcmGWzuLZ5rrUjEu
4xvyVmIPpFZZNsS5AKHhmWK2zAbW+eNTuz9SfjrEbdpqy2CKrW5KtGCdKVhIrS+gcpuDgmjXO8YU
EDCNmjkjvg+kLzVrQf3Iit1RnKcT7Cv+T4G+FgHq1O2E2c2jNOLIHFiodeWSBBupWheU8iSqaLZl
m6TsunaqF0EVEgEb5+B5LMhgWMG2lkiF8RKzhD4mdxiMFiE/brVnqS6X4CLCK0B6X8qmx82Jn6C7
ucXOGaXFELsClY83CyozXttu/qw2mdKPLkkEtHQpKUois4oQRPCsjwcF7t1EHEaRGOip7vdSo6LY
Pr4s9dWxycBFwp8Vy9ogN2IhbucB16sb0/0oYLlIL5fOWCS8dp6oNl86/D+DogH4ufnT51UR40HD
yZWPMaTwQHhQwAF1TYuIJzYghQ5w33Gd4N8IAEpCkNlwqAVQpEb0sF9SL1o4EY4AudibtZtGPwvR
nm3xfC2e9KlQxcQq+wmogAF8cUVmtFqk50tlGvLPAtWRsxtt7Y90q8xjiSNTygCGO8s6IisW6pLc
YSnZsARO5XKrY5Hrs/44YCn1PBO5ELJfV4VomJT3Zuv0Byh14wxVdgeQUjYb0Y/bCG+So1jQGoMk
TcWqYKbHW+0EHYsmsOw+na+buWXEPp+h4lXbfCS8cwSxOJZ1tjChC/snoU5hvOOe7gvU2nHtqrJP
TB0b6OXtRsQu+9a07YhpwcefuRyV9p19IdHKeSXrPl3XgQaCDpWbDZUu89owx88H0ZlxoVEYjrz5
05bfpdPN7Z0Gr3eHX6EwMWMvcsvPrpivyB1nt9qq7YpzuMMiZE4aWbJm4n1xvznFQ0YNXdpdtILo
3HXb5yu1IKiWbLI04u+AHABsyVmrFaoCt9qwUaBOC4ZKlEzV7NyFiHLpeAkgiulfZ+DEAhGnSIeu
eb3PEMoJ2KWvQfiTN2OxvkME3lXACWX5oS2JxdFVn3I5ajTDqasAW8hxprZ5l4D9yqQ6OqAJ4bmk
kfaUMTlKsMlglGWZ9pnkdtW1F9189iWFFYgDRJKR5gl8n2dpeNvu1ErTqgoG3S1SIFFJe2RctH7X
+8WVYI8Iecbizc7pUliqYyT7+XZxRU3pRSdTEux8iBvAFxeILj587suHlyquIubgFa7oj9d9QzHg
azaJ0TczeGH+gYIZ7CDEA1yrIon7SNpP1aIywN7T0nDSs8dBL7WbK4e4Wi7lTnO4XJC36wfTqUms
vRdTTMIzlJeyrVpunJlplZNPhROUj+m2XJuaXTq4b+otkmsAn7nYG56RPayrRP0enQy1VDrudNxE
NEedlrC62TO3ly8apEs8GBCmGluk7PQkJ7dW+GYwE+5WvqIl+kVHxtJwPWTZFiwuycfoYqayXqib
BB/TJeELb64BrVEvUkUjdZ4py6rIVWXqBZJYfq3p3FWuZILruqlVNW5eIpjaMEazeuwFPRPlNpEt
rCXl8sSL0SfxXFD/xin/FfMw3oPkTIu23KIg4dvdk4FiaNznP11016P6p/PDl91FuI9ufPpVHABB
VsegrU0TLKsFfZkMsPSCQA6LIRrbDiKxwBWk3JsAUVdhG80nGTbHr3udzJ4mMP4/E7fz5m3j4221
rKQI3o2wJ7M7VbCf8Db0WyxTuhL4OYDwfta6u9mLeUBhXQ3pvbRIpt+HSscRicw1/585E/ad6zAp
RM3nOdhtG1U8N9VKZ9A9G2xQY229S/JdwhVXRplV4kxckgudPIdbkd2Efb7mL2/hp+gOxVi0e3rG
7Cxz/1N5ltlgQg73reWqyNxTMUSwAcKQhMOtgtBfu5iahkmBuZR62mFSvzbHvCAiVc7iPWOQOSQu
+NETXV3/rjPgOMoCOoypnHcI7lGIdJ5xpYQ2L/AnD90oFHg/SDF+/ZeltARCwvhui3IsGMZEKCVK
PO3//2b/WvtSdS2R7wGIhIHYgYeFwmdqTnV9L3QlT/BIrA2C0vZF7MXVcfWMA2MucDCWPla2YsMi
QNradO0Mi7aM90qtpgZI6PbbRypVe/8eRdbJWqKeQAek1tmHgFAYhvH75FFkSZG4sueOq+Zxu0tO
vZTcfZgnzU/5dNla2Rl/M/S6cw1gouxfQWLwpzbQhZHXjn/9Ma4fnp+OmCBjTwW2hbCzLldASsSl
yfUTWcjjXZ6JJaKpKYWo3Z3bmgB9aEzzQMWzDYdLXJ6kIOn1jzoptjgw160LAvIA1TvWf2Pu86Ri
anpxLbW7ej1JCmfZ2tqFEwDG/Axo+hwhmhbqHO4Ze4zXrewQVz38y1t5nap2511ckd4MYimTdsWh
F2vhkjnFrolMpleKx7Tlg1tdqUKgYxvrt9mxLh7ZmjLYWoYZvvvDiqrek/Wv2crd+Yx5r6/H4Xgl
nqhf49xul3lqSfgyYKWIq6fyT9OeQp06P93XB+Oh2mqgXlvmtwJiW4oJs+QnUi9cgxzHLZEXjlv3
7Ef2CuLnLjtMEL0VICJlhWCVfA3PhArSKT7+Gf5fDkRGywIMVlPyS/UYdyZv+YffdU3S81uEIs2w
QY/HHCjwFS7CIAhKk+sYjQ2k/NipxZ1/rAoGHcxEhbWCxlDdLX8d4MTJfEkNmV3kh1vy9Ruz5kG0
IZG+xSVIEDcM6nUggfs4o6HqQC7pORIIR/0T+wBHUA1DdcYFOngOFBbpdUjb5IpgkuFum68WZj7v
X8fZ8nDoOGGNDWQfj2MYzE95WLY7zKmh2wgzkGRGZr7hR9sUJeEO2RsA7qmaWucovWKR3MGKK8CK
KCIfUKTMoOKMmypFK14yB/4NeYxn2d/tw3Kh5Ystb1WpAh78G49+YZfssCesP4jPe16/SzGqwmjA
NeF5tXBertZAGp8eeNpiDdFiZIzMSuYhRypVkw/k+vEzYCxDhM2AmlPR/dzHuDAs2+rJaQUZQhqr
mk5W5TVnVRHFDn+2eobhD/RE74gFEFcIeNH4bt+LLzoYFH+p96XrpxUHMsATxlH75CPc/k43nSTw
YQC0H+49rXA7gipngqhi4P2gNvsmowH0I04R15cfkxYPXeCG152OEKkcrCUA9qfh3aHx7vYEW+U5
OrV8b4XUI8f14CsKahO+jYXdAtyV3FHervuiYvQyHEaXq9lBuFYNrEF1wQvG/Y050PAmhcVnOEYW
MV13gpaz45JOBmku7nqh7OtlCCmIXT8FHqCngWJpSzWNmaC367piqOtb1OvemJvMYFbElQSUbi9p
eJkzRhBTwm2zbbkclAgv4/s7lxlmrl4HvNTNE1bA0bxISePWiuskNJpQBkZVO3Td6gkpwZOCoaQ0
sbHIe2ZL1QRzabBLq3chNwxcG7bLTNePZCffRyfC8owQbw7YZ1HPPXGorf3/XGEO2Cpa7ir1zqwI
9BPy0G/oBUkc+CzofmHQQW2od5VFADIA54kgpUM4A8YzZ9EO4HFd2Ptum3FGbRhMPxsy1CUvZYnS
/9DEuOg+JU3pJwAIzcgLD440m6lWIWtyEZ2y37q0/f8wReP+0u4bgo3vUkJetwHGFXpsC4JF+ZXK
0zZd39MCt16Jy82vSWN/7UVnXViAo7m9SFyISJNUuGkoMIA+3XyxG7ggIaRTOtS8e0bV+rNIV7w6
OutPSj6R3nBLO7QhMZnityKoeQhoIC2PZfCbpHGCSbc/b/+xGuLaEHQUOdhrXDQ6Vjwk2XTKW8Ml
rdZqpA+xnMv0c27TMLX4uVZuvFgLddiXAVI8JYPc8VhblYcX+nwLY94FVGvH9a/dlU5mW9riyqCY
jp4IRroO4xW9PhoUK7ApcDUlLWccIOU3mhPvyVBn2tGqgyPgxKeOu0eB5Ao9+Npja5/KJa4Pa3vA
bWq0j8KhYQm0oul/8qbzEiK/S+9ACX6a773cahCCKIIwLPhsG7MlYihMevFMJ2ujsQfjX9LmxB+E
gUQ69dcom9cfHX4VsKiSC/JEbd8ojUe5VtYZA6i604olAELmNFd+TmbwELx/43R6LbEkHQb65S8d
+l03iAOGZB5SYHD6d53lDrl76hYNZj4i7/2rdKQ61ifoKZWCqTnSgegTJZXlo3gMS/lm53F94sCs
/XgugdHKuMPy+YJXvlR/vUKvavjO3buJU9hyu3xp7Yg6WybuQEo0KE3DDloFJLHtyuaehBNM0car
GMKRLl8rccanJa6b4Z3gfwb5EhFqpgOP87uy/PeoKhQHhlw+AjFQmQCrR5DmhO33+1fAxyiZcLDr
zW/BGS594wjqwUqR6OlgEdiVpVKjvOmWlpKZ9rlOJVdBU0QEDBX5wmWvdLbB16sqbRGA8kjVO9Xz
ifTeSjHGrSEJSbc9cIWlj1QM5OmldHTXTWsKI8D7kI6ls4lyF+T5cyJCh/sF0tsXCfSJ0Kj2qh9u
Fkfv/1s0UdiND1CoU0zaDKfZTq4KgbqsKniVlmJ/fvfgdslqLhRQIFkKDOA7PH6YlF7Ei2yzwAKM
5pXLExaJ7sxXldVLrc0+35Jys5fVs8fYpYEB1vedtinif80zPPxIKxxrxo+gktaxmWzph4wh05qR
YS9LQUojeGIThKzNu63dlXOuMv3t6cF4nmDpEv9t+qwUYMS6IDNPo5MT1YMBpk+atIwA72QjMp7A
OcHoacSOxdGWWkd2HpR1BsISQi3NESyRZAlm8hBX2VrFY4Ipg3Ldd4SFItlDB2gRlTDjvy/zJJdz
YQPTXyUja8VPUzORWEO9E6WzbpvHKsAxy4zAuvxxYWqZuRtiN8tTXzB4bEtYNr2kGwvdVFWGrCl3
xE6E6d78zgPG12qMMnJskSc1qgv6+ZJq/x51gW5hLl7g3jkid6IZLKU4bBxUJbfmu3hY9hk1jfNM
nsWeptJxUU/NWerzRBaKACMZf6NFDpj3uM+8CddzzCtF0xtWtx4fE8HPK6rIfGgBEXkYXL28T20D
Dg6PnbSxMVKC/FLI2IA3Hj9O+EIgOEcaX0FbspdKF5OOis2NSww3zI4VAIZxxtdjlZo2DlHO4bkP
MP7T+bIEE+QAA0oFDn7b+K81RMXcXI4TJv3t+5yU3dxIaRWYytYSgwGPLd65QOSye0/OUmg7yExx
UFYmpXkklRo19VGx80wPh4bx/hurMK0bjTRt3xNC3f0Wk6ou9wfXgQVZV7wotwMrmnNrLjIKBZga
AdE92hrd4sta+1AtjC0ao8Z1UzswS8TBhxqS0xiRWG/zxd+JqOozBW2tmzKv6vrIdYFuWkUrLOzk
KdydWonn+vv/8eQDzZCrokyCoGXCwh4pPvfspjNmISwQRkFdmWP1inggR8GS/xQv1qEnni27Pfyu
6frv3Qtw2zF5nvCG7HqZ/a1nJhfhZNGHdS45Ni7sssf7S0IAc2phkiMk7LoUk0k18h/2wgdWhX3B
hiqnvVZ+lpKQgEnBVavT2fChCtxL5GlmUy591L+jaSi/rFkyZfSfThdLoz7UBd3xVkIdjy/ZttQ1
fhUgf6NjjjQt534x5Yy0ZKYZs4Idxs/lrGsZ1DBkQMSWcr3vWvT/ULoNAg+yS148S+OhlaPtiVAU
TS+NbkU5cEIK4svc6NEn9btCelvuwzoy1SUJK/TAOuAT8rNEbYrrBr0typ4dNaVw6idZRqg/F+hA
ec4Ds2sChXQKb9eTYQ0LNjutYpJtJZnVt9xwdi/tF/VTlISFAdoLqkWZY3jKlTHtdmDOOFLPZod2
hwW+dsH+QEiYJPh1JGjZEcayDH9YBGHfKyoCZ5Pkcj9iY4urMuQV31GIw3RIglF2EFpNsok01yoO
s1m7MRvQqUq9SmN2N7qR++CfDxvr0YTRkFd94UmHJAAxsWGI3X8DQJhed7xILW5/PeiNUHcKmuIA
TnWwHrbQIdJhGINLHDzKAPZA+g6ivAiIbJ1m/3mF6pnVzkOOlewF3e6yHXV+CQxfjAyhnVdoqqGK
z9vgTGMvunaVVGoAvpjITnOQVewR6v+w1Vi3S5V3Q1y4K3yeO11t4/C2IYycw7cACu2aGn6xkB84
A80IbD0AK4jJVfUk4taYrK+ai0RQftHe9tAcSxaLGRw5I5OJLp53ZLGNAU26PQ7kkYmY9zaSxAR+
WjQSRZy7qp68whaNB6EW+J83HhTSfWnsN+OElZ0GGaPY9rucJBMpoyCmXC6mvjZHjtNgpKwSaz6F
KTyvEsDatYOhXgn8PC7tz4NWMT/Dz5iionn6kc3TsbxBlGUcd2EY3uShwQVsxbUamWE8K6t7k0RE
fWwKkeXL0MOdW1HQbHt0pcXWiogoJWFHxAWVhR4zq3y9dMHbpZpVASXVbpmxWqOclEM6dK1udsoI
liUxGYMxt1L/eTbVO8y+fer+ptypiVusvXcdf7ATFbdiew2ZPQ22hla5s+IBuKujeVPKLHCXKKZm
H8zBq/+KgcpIhE2Mx3cahPFOU7n0Azuscd1+jpTLM59zgSoZplSApMLTbvpGp3SeB2A1xAFQN8un
JNXpzF7VQfQq911vRUw8+AHGhV0XdV1My/o3T3YfXaQVeqkPPHS7a+AjHhCvw80/rpU30NHxfm2D
NgOKYApQV2yHc/alebwI618acdBAQOlCKUk7apLe8k1QFBO4kAyFYsiD/h7iIoRxvFayKtSPMd0j
/BfQY+FvNRrhd7o63AoiC4wMLvsaxA/W2MENyTtDiBbKjdKy4PEBAF8NDpELe7KO+E8YrsalVcmo
4uo9q4YZrbTBE1wHHPpcEwKHY8r6GGcGBQIBhwqnuYxj8iXpX3UhEOhT3WOln+QrJ9vk5LLLFfz8
sWfw8IqUGYdzvMzi4ZOYt5vCcB+ek8aTbEBEtwrd6042UPBfYouTTTTByDclYg9CS0XnIiM8Tv9i
zi4zfvUxpPV42VveeychFu2WSoYIKy35H0TDYislCvSLP54K+6c3YkeYehWH/R4RHa9C70ylv3DL
delan6k+iqTNiUoz6IB/i2853cp4VMlr1hCEHhAkTRjvgXsXUXwUQ/xZIjYXIY/xlWgYOdP45Xpi
flzBebQczEt/n9/eKyV0Fu/JtiFhkdsWy3T8LqYi4y8s/kBovLuQQa6Rir50mULp0HQgI4xzhgTJ
hZVTzPCqHkktoh+QP4Az2gDnfZ+1d7X8eJXNdGVwt445cRGX3TY1Qj11DtyRz/ZiTeP2KreMF+VV
isuwxwEZPUdFB2RSVyhJEwuLPOtS4Kc1iuUELOJn2l1v6aWqOx5hmh3NMJY4H/vlyHj82fxWhldO
GSAU3tADHz7Bk95iLR7oruaeHR7+LGnvYSqvkA865YJx1JLdFbfFIbk35zJIQuaqZKsZJ9c1p8+h
mpcrdwL41AXJJeuSXMZxqndmyrMbaqHOXz15C5BuUSq1ipj0KnA3/D4uxCOWMdhRGkRtZZSo+zoZ
+TqainL/4IZAEuCOx105Eq7w2JdNKeZZYS9F2X0mI3Q2dU9vlc87r1oH2ewS2Ls9GF2uxsnUjaKb
i6czJE6l+skuZCs3QqhiQEHEyK5AxCNjU2h7KpUfSuWiuyf42hqG19ddnmuS/jdNqf5j4biuwb84
tT/sXQyEB07iRcqviPhzHYMPXnchcdKhAXPHSdSjtO19CRoVo+bar6r4Nn8cVbxAaBfXAEzGXaUo
Vrc7BEzd4P+WCk7bzrVMbhhLr23hAbyDssvzcp2JIvpWxrJ3X+GA87tWmOLpmDcb9+BjrtcHETlO
AIt4KUDRodSeWsqIilt55cJl+zykmuhynZp0R16AQBiP+w48zFs1pXYOY1RjaFhPY9MSZ+wS/w8x
7y4nD0VwWY659AoRxDd/cufXs0HPE9eKpZVSozMsh6gbTOO8xGPqtJz+p+zEfk61aKBfFeWjWuOw
wHN3NAs5/Vlsq8s1QTZ7qaDVOvzOSMs4+6Te8CVcigcB7JQUGUVEsUt4wiiSsOinqlOEYWIut03b
7kR8us7GGenZihJjS7XTHZWxdcMQ2JabHZRDQs23D9j12RQNWIC3JXYgD0JxEpJ0n8s6v96J8Y3v
xYTtO+aM3En0VM2Hou9cBQ0aEm+wYo/hn76zh+jC52kTcKvC0pKT75PnXL5Qt1sNME2qADCPocuv
pN+IVJtQS/EySrO9dcjRbKQmlAsVtuGEqgSnRMt1ylbSrGIJDfuJj5ySwlrNnb8eF3v0h80CoeAs
wGWtLE7TxMeyM5TItZKgz/19/33jOifCtfDeGTG+JlDaFMZHJFwZz+k5NNAH7ThNz/vuYMy8hDNQ
o8z7Hw9jj0RwIbo3sRjcyWLrO3YfwKx5/tnTnIhpMB3UTS0WIOXEnlL5gdrOXime7AXvOrEopojd
o9+2uVSxHrPZEw5Ch382FvAz+SOqhNyxePLF0+BgyW4vITxSrMmry4CjBeWRKCDnSZMWdNXc2FlQ
/NB+BEX+XTy+agc1vwNHVScPfvTBUQ4ENvP8hv+CBvogoYhcAHUO7QfvI9/2x+2AiPrKFX4QNvxG
WC0eH2bgc27oJnzlJQPdBLCbRwtGI/qqDRvMNSTUhU4C//gtdkOvM2MdiF4uh+nHadFdcFw8BJBq
0t03/9y7CPa12MyaF5S9/xOJ5dIzCHsECL5++v7+SP7PJQGq1iskUo8E27YhID37R9B0eUoYjphy
u3rGZ6KhjrYu6OLQw5RlVFzjLEMsTol1gWea/qUBPMRllwUoKMa+ePQy9Q/+4U1TP926ywD0Knh9
+R/p+X5yxs5wRd9mVueQOdrZquoT2vVUBIarFd5W+08+AeWKXltCOAwCAAIKgs0h8gpGA6czDlrL
sPHQ9sC3O9SdqCt1pKjL0E2z7pLtZhug/S8EmrEwCkWhM8Ec51F3MNCoN+E+9zpnOKIS7YPkL7MK
t0XQkAVadFo3JcjeXqLD0J9mcwl5GyjFNTjGkQL6UK3e8YgVQPkQo7KvV+rS36NiFKyEgwiyhtbH
wLRFW/1+jUUVcEbk1f/k8pocDvHkVunlPDi+q6PzaIDM/f3nHrbqXmaeFH3tnujD3Y8hMLwwaqa/
lYy9ysMOoYgT/ZQf4aS6sgniBoMLrX6tP2DhmbbpmAOWB1gbiGxB2cLre39HNEb0+NwvVVYfNnyI
8LzBCbOD/3lgv6z+YYC14KrL6L7zqqOelcQqJnnpjMO7CFNihANS5HEdTkLz0Qyrw2rAh60P2052
JvJCZWn58+taXwMFKbDrR3n3gQRbw71MG0/sBdrD7JLop2UAxJE1TS2xKPdQ67yAcDzEkyR+VGks
lWaN3EzdX3wTKLJ/frZ2i+H4fwzu2jPTi78vn/sEtEoHO1cDSeNTWWkDYwfADhC2OpEBZXK0uNo6
zYGR1fwEGf034aV1wSKJ44z8yY4Noy6V5qetO+vnigrSFGz9Lnu639egmNp88PYHQT2T4/htZ5NT
R3iD0hBThfLKS7BGDjYkFK4DnOSWjhCMNDZxF6hej0di2UWZokNm2xFKgwBvygo1EASTeKAMxogL
JM9tuCmXEA7Vj3TO+fcCuD4iDoEwRkz+d66mgXkZ09eZnxXne81xJgsjnBNZfnhMn+P1K6XhqDpC
cyM7Op693ek4UfEbGf10EETyy/wW3cgsnCdn/Sfgy/RN10v4hP6rXcq9yP3q/IpDuTVr5XNl1cEN
GOBnCfNb8JN8KRosjybW9fQWeCgF6w7bwyLw234nVkaJZ2S/0TuFIJFUpPEL4YbsDLUOO0Lwa8E8
c16LVPTvKfwFjvLBopGk1Z5kIzASW3wIl2o1kOyQvsvqr7qtIxq8vsQ7eqfohSvOuFyvAXx66NPl
zhIwDHI9y3yX5776pvd3FSPWHV0eDOm4iG4ETlBY7gThvwSxhxmMNy7CTzDjjoxnxtGxqDU9+2C4
SOGnDH0U/MEhZyLVmu8Eqq9z6Acx2jPUNAadEmCzAkP2LsMNHTJJih0yqBgnpaNJfQD3mJYT6a2t
iDiVKeGvp/NBpRSI0E8kDNOaw1RZqzaEbzhb+6MoSHl+sZWBL9e1H65rFAED12IyRhPa1uMYC5HG
uARX78TWs8vH5mHN6dmjnuKjXLCxYXdz55AE0Xi7jYxrpK5j+EmvCsBXt9pvtDGlIKPqWgmsrf1b
fh5H88bZH3JfHAadyBK5R+msgvKxcN8w1L/ULQAK2IhxrSQy1ln0QmvVLpuuEH4f7N93cUgpxazi
aj5eQqSMRe08/e/5ay6WMB4SXtjX93cdLSiCZUMt3wh1IPlpLe/ZNsORl5R5Og68FOkmTlFILVEI
4Z3qiAn53lstQbIU8BK2OA45SCCxR09FPev7lokfmXcjC6NRKOdciU/rLdovVlNFOid3A2YlHIH7
QClw0cmvC231qOOWrDQ+k8ASKiXJrw3dHacThitBp5LsG2dtw+vzlSpRGrovUWK0W+xOcQbMAIKp
v1/wmCqvwixOo+tcFNCMolB74+w51x1lpagO5akVPN6B4Se/9Z4tZaGesBqCwwaENtB86/L5ZCPK
YgBsFN9KNBLhw+EPq5SQxbhAH/z+hv2+CWMRgkkL756XO+7v1cZcTTYC0G4AA1mjf7TLhEqNo12v
JXcKYO+QHS4vz/V29UfmkIwIZ2CcKfKdzqoyxGuTFVC/snvnvy7O8wSbTlOt0TSb4x9KQ2w3ZUy2
2RJ84GD42WsPGKH/ZzfWV9/udHSXgG0I1CPLVN5gZuRtbA3O0q3Pk4D0riXDvJXyCs8NYcw/OdYC
CD0BOuvukz2NPncSYmpKPRIAHV2cet+kaY2mRwo2pVk1329s3bzY8xPm0JifIMHFMwa1jrkB8WGX
5fg7T2wmND6wT0jRZ/5tKTmVEIoBzyp9V2Hzs5jEPjjj6cNDdrQFatKTyTOvx0IQiSYEG4cowRst
yVZJPq+ncskzGaSCcxaOXjNWommYgkl15deLZu2UpJQaud3XgH95SeJcPz95n1i4RJDyMYd3hCrA
/EYbmoav5rTo7A8zOsmN9MeHT0TyHlwTq4yC+jE/ar6qlxqnE8NN+jJibF+3S8QdLHBBaM63g+yv
BZtWkGxCK7tRNdqjafITIiRRmzSb3dX2RXSezv4HTuvFjAJbE81Vtl+AwZPGKr1B2KERzcaDJZYa
cM9Kxh3o7bkgIPijxiqw325oxr575Ioqk6jPyqkkrRATFBD4PoZtIafMP0nEu6TZDTz9DLhtULfg
DRNbaSC2TC9asH7vL86k6nxDzZ0M2GY0o0nhtjt9N7q3mg3pewd8cSwEwCi6VX6M+4M42khczhUy
WPvX1uunUCyyQLDSIXrw8MHTn7KU2jp/yN/uzBHLG/WxjPZ+1+ootnD23DCeYWaclIggl2jvTBrV
EiolFuU7MUDOnoQwV1nRx3gzRFZi/UMvgqX+1yivFbO5Ea4hxkC/Za+QdpusJa/heQxwZ8BHAQU7
XvhPcW/qiTeBLVnuMHDooNaayazuayCBZu1Gezw4kJ7XW4CU7NFuvejvaklmmIdDUQxFCtJJCqS+
2+z4E4qpJmiuBuEY18Xa/xIy8WIjYjB6ZF8aA3RrfYPS+byur4tO4Ex2o5oPoI3OKDVK+uTGDzCD
LLj3TaRkgK+wBV+Y08DpTSvRuSFe15RS3ZdiNjbqb/L3i1mlyT9LuPIEVn83zxQIHiLgu88YyB7W
p021raAr5Jf+fDYdV85g1lg/UpOC9LOmjBTlD54b9crK/YpsfB1C9WwG2W6optoGXqdttkirEwR/
yFrhYKtVGky8S4QsgI17gGRpzxVbyCvlK3rrvbQvIF3BivY1Q0hKy38pfHPoySQvHRpAJDxxIHXI
sWO1Q0k4heZ+nNkAMWzRUBrdmhSLysXuHFwfu98No6vSazI1y8UVd3ktBfuB+Z59NSgObWfAdctH
9koquaW+eVx90uy6bQOy+tuVTWzj/Shj8ehspdxigH0Ip6Qnj1nZuaTkRQWaPg9QsEtKtMXqoXTf
ZUFkLbYNA/XKCfoNstLXg3NGWG3myZRFGcmo3Q9/K2Gaj3mzbqgGRh45yER3mLHhBuXKdS6+e7OM
DRVpYeXS/ZebV9qdU1+s3UlV68feMvveAJ2Ksw/YjrGCUJr9ZNS1CvkYk5RA+HpKpZn3gahDTh+r
hENXEoRCpyw2QUhcXMOXR3ZlCcM8WnmXLA5DHcE4BVSwU+JSzfotuXjaJ+UXuKtqn3ZU4E/r3Edu
MwGR9AXmHvh0Jkssns6yGh9RQSzEB2TMn7CXbQlLnQ7rBMp/2HNH9lXT2BlUjbdeYRGVl/N/9WSH
RxfOYyxXEOSOk/FHXTf1KJ6N3nJcT2uGFEdwBh2iIN7PNXmdsz118qj1Zt6XuCT1vaKukv3u9Mj0
p2fsCzv0pf9ZYrBup6xm6EEdimBp3vdZoM2kGQzy0c0Lq2cr8/bdogETC6x/6nve3BRQV8l8DPdC
0ZNTZPupkfwmNk4NiNzc+00WJLfU+eRmtxrG+XtkatEjPCnD8LqkXrhR/FT51I/sKUNSnkmLlagV
2R1a1JhHHtFlWrW/NBIn9iKQ5YIRPtr8g2YREHthin4FhorrgGNI0yZdGZfzAUgtSxBOJ5uHgOnT
+0KqVlDW9dEebhbZZgsiCXey6/brU6zJmLZ70bHTbh3s+DUFyQl5hYeZxZPv1xQDLwHdehmqjcKU
VYCWJqDJ0BBXkG+Fc24149+BrIwu+DA0FMbbwQmUld4vizb1YxtL6V2HYIyQJ18r//sFmmnnY3jP
Ef4QqczRb/v1PBybJf9ytcMky/LCPOrZPyaohc/8C69W4S4rMdAO/PudupYm3mq3kfu3Ru3t7bfH
/kRrcsANTlnqPcWbeP3NcmmSwvCSnIWxo5qw7Kn6j5Z+0hmIF+f44ypDNvEVQe/duu02V3b35Nmw
9c0UGgoWKFiBANVGfMtPSkyuvvtA9mL6koNjOZJj2rim1U+PcFL/jbQdL9/ZdCnDkULzGd0GAp6C
y+CMKkEnXWZV9bGiXKuVXYrBcNrhp5j9ANEZrQhIIfnKEBIpy8iU8ymi9FqoYjUthowIVg2dMGUn
OZaSjTUrF8JuI/CJC+Vp+coblh5Df1ElyAxEwzHgwKhigVJHdxtyBjpIHJxKjpG8hAbWOm06SvIK
WFabJh5BaqxFwpMU6oIfRa1LZSh6OyPHAesElQ3XnMPvIrOKClmXXYHHkXkO7iVBSU2dxOwx4xEg
gej4774rC1PytMPkump5J+Pa6bZ2S+5jzoXUmNwXmaM8j1zdsP0lZCGEqhZzr7CVZCoG96uCnUkB
TTQG2aNhjidCvYACXrO/h9quNb24sCDD1yUlhQFWNJJ+aavDezDVyPS2aZQOPKWn4N+gaUvF4fSj
+vr02yfLgUXdhSe7H4pY01uAQ6OCSfI8wdLCLUpmVTsc/wK7HaOV9lJQc/iHmLsUMeI1rAAOd5Wo
bg6VS0qeM4TzY4xAO/Ppc8sr/rsOuT3U4CLAwKcnQpO1axeud/EzC4547Si8liPb9rW75VfVjQhP
BF3q5i+6Bk5lcf0Net6cor4Y4+YPBSk3tL9lVBjSsfMiFrmn4lQGanB56qvCNoflg3YZf7IMgZXv
QH4yJOI63qNDoTHccEcJHS+k9FPmUlQJbk5j113ZtrPCqhGUgIUYGJ8ee7QfugkK/4aa7mkgmhM0
8e1YFXqulIHPxcc01hSFV6QXOoVGxn9/uZf2DVG12u5XAYckICnoUZLHSgn8zEI/Pt1YGCg8eEhT
UVuhHKWptWYbCKQtEmW3HCMaD/6zlCrSh4sXErp9wE3iZNsEu5DwTLLE6e8DowrzPPq4qZ9iHR0u
rnqu7bPT6pQJ+jURepIYPvY6e6BD/2V374Ao0j35lQx/ZQ3ZbU9e6jG7bE6jMMivX1rir1IIWwZW
wgFfPJRjzzcRhLbFYz631CJIX5pBs4u7ddGNrDf7w9P3inZ9IKRbhZbuAKqJEQqxitR5zzHF61Q9
MejrsGJ5a8yDgInCGeaB3VoxbkPxgBA/p0Zre3Di6FRS/q42H5s5bEOPDADA8cIWHuETpuJfJU7S
Mgl2oxq1IT6Zsl6Xz6TI1frbSy4cBCp4+qZ+vmiWuVX6NqcTbOdLAluWk2ndUAPSBQrP1JSO8gZA
72UNEqBsgS2aCNyvHUb272q5Wv8ZClxlyJHL1ELE4xfuFFtJHGDUUYEqcHmDigCiHsSk2IDVuJrM
m4JSFcL1d8TFEQEfsLWRQnaU+S7fNoPevcJKFwbO6AkbCcXcVlfcbzBBj+elIwCB+FHC5ac+ABqI
875rxzJ39g6yCWusoVbomEDnQxn31Cz+AmA9yzFH6dpS99w7Mxiw5io5dJL2GSsmzUksptKUTVhb
124/PPPfz+p3rX5Ff5+Vkfqt62d9cOW2X6OCY8Sdte1pxUAC6aSo2M6sDX3qrp8UGvWtjRNfqHEN
2wQXyKpUPSa/arOnb1sxEAgHDuPEqRtgHXGPJ44oHzQEhNepMv4O2th3S5dXLq5s+ppOONtVlcV5
/hja8eggiIHb/rtbkQTB39+i2pVyoIHWWtMz2gNrpmPl5m7J6Aryeu3wlzEvafMuh1uF9eQWQVCb
+tHhjw5AA7RN7soUjx1ZlUCjp7BsOOdPYZkBwbtN46t8eWRDDC6/1DTmRU6ETjQhX7gqctYkrMoV
87p1kNVuOW1sa5BHG30xcHu6mf8a1+93eStomgNYt9hjQCtf4IaikKSwu6CoIAjB65bd0esjADPt
PHnTUeuNdAlQ3YLB5R2j/OSQT1RhxNHNdTfVInn2Mvlw1s3/sSA+rb3YiUvTaGPfiQJGiHCAcPAa
sU14MENrYI6tDd3My9+EKZW8f9oImytgTBNH7LSnCct9d7NQJ1c9fIoFQVNHYqUpQUX2YO9706Zk
SuW5Up4/d6NRL/xt3FSCfv9AT4yrTKUGzRdrFQo8nVk8HeJNpJsEbNqD7wLQwP464vniDagG+ZRA
6mUz4gGjfvFVxHpk3JkaIptteOm4acfdXKqYPhBQzXJKB+g3tARTrf03KYD49P2Z9nLjRX6+b7vl
BMPmruqyW6cQ1X8J5/e+rP26KrgKHnQbu46VCAk22UGAvqQf5PX5c41+ShbgezPFhqM4KM8Wn7GX
L7FI6RZmXjPsnLM0xDozF3DeTMWn8SqUu2a/yev/dvf+Zvz+VHbmTCrWEnyeTud084TlELvgn89p
pdYZ1UTPxk7jPRFGaBtw2O4mO5/KZSIHvJmeBctDSRPNahNdty7gUPoZX7fuMzC72u1G0BeA/wTn
I1xwclNgKKVyQtoQe1njUNtALk+HZQ5k8SthpZwmC3HY8CnuC9ndw9A9NcWyDz2HY6R9p3zf+qCL
rXcMCuipsHJnosaNHkyriTWOxM9ThGK6YDlFiV0XPF9wy5EBH3ublhKsZtFjgzYC2Ofzm4BZM4M6
c2EHb2IyDe7kfzPEm/7Z5c4JHof4aUpGCgYnvi3sBugYPjOFUxbl8mAUnX2Qy4Irh3aD8lp3b5iy
n4gUwvKq3nPGAYHkpsFQ8+TYVwBiawf9lyLjXDW18QSq0GUnOMDwQdnOzpNh9OurH869mA5nKW40
+0BwXaqJKj5optmmKCAKYNDocRbQA7QPyN9+5NXsTcw8d7HViJLVB+BaWmIi7Ym99EflsPWQUibR
l0h07TIgN/Tu8ZFpdn5EDedzBz2JQSX+d7FGIlmt8X7rfZPuK1i68YU+ZeGUSGELsqXIDCNS4q4+
3I9v3egzsQzH5x6bhHdeH/qfrMBX7PjFku/G44Xzfbdf7De7Vw6zKIW4IUREW0wpuVQsScqefVNZ
R3ZMih4rxzIQbj2f2OSCjbMXXVDflcv6+M9HNgTJVRxeiS5Dxa1esXuWM+UUJFXdbEvT9Azs8EbE
aUvbfnXBSYtSjb3pjK1Y8DlaRM+rqvTgc843nH3L08lZ0StoICHV8rna48mnSNoy98qO+5EX6GHf
wy9kVQQhlSR2YwSzhWuTSeKowzR+CdDX5/wi25PGr0pwu2RwFmILX784UYp7zpJSwswObF1mfF/X
+qgDv7iSnNxbQjV266K8n4774WxCnWBOLn8NkvzE27wku/Upnm7RCC3y2IkD8XK1XmrRqzCUuRg0
1rxXH5Xj06bgFzlBYl++L6fXBUXgVzoA+WJFLnWU23MQsMxGATSLuZSvpN+HKuIWI7EU2IlGshj9
g4Bb2cxNbrKw30cODY7gdtAPmSZRN3xHGlq2TCA8zJ2wz1uYreZ9l6z6hsVbOklcMexRMayc/mWW
djFVVBt/ogceiHg9kGP648wCimvFOwhhvAzf5kepvBoESdRRDE8wNUOfk/Dra2Q5BZ4IRAj8jQAY
+ZbkWFZcKMDxP9QAnYNdB93A4H4dEPsuGYG9mIhpTXJ7E0/A0qXuor5oVBZSXBUM+WcBuHmuBsfy
wuts0JCiruYmOlqJ95jv7qNxRwjAoXDJ7wdewyB3F8CMYsPHWCglwCqw2JvlMxsNlKSmfGBUmAWR
d4Wj9Y8EqJzVilLOkXy0nORdJi35J/Vpq9eOCb4ghNYAZ5/w0n8+sLffYst36HJgF84KgoYVlSlM
tgLtTjq3lNBM01WJLLpp2o0CdVVr3ynIuMTSSJcf3rCooig5ui28now6VNOUx+SCbCceFSCGlEB2
hkRgMYr06sAqw0Y0DyO42dtM3tMkYGe+CeZhLnEoroMUxJ/2+PGhNC2x8Bq2DFQNUgqHIfco/FBB
NxAjXAj4Ey8KKSsFRoiv1O2C3z5dS3ARMXRVUxyBC4wBfazW1G8zasuDTwMKbOD7eez3mz2EdWvF
+he0LqnWEW8ZOauhG3+NIpf2ok3cSUg1uH36ts7eU/VnMqxfAMFp2V0p/zh772U21vRNgflPe1Hx
X42/yIlGvbgY+qJK9xMECXuMxHhF9RHFJxISsvKK3bWNkX+H5urlML+nCzyFTF9GkqXodLnFsoAT
FwWNu2PSgTFxfwCz7OefU8fjvNqgDPJDyd0Bao8elakBuhgx3nHpPk14E2fWEoknP1wpzt36N/P7
NTt8yCjL2p5FPv5Cn28L4EVFH6sIvHZIIyysOsXRnh3DoGtTa3awD8nlCfO8w2at//hgC9kgAkGp
OeIIEecJOeOzz17wWRCB414FhZd/86+Otevn09AyfT/0IWxvWgfCWrCPr37NJ3lkOFt5b7NDngIH
JqWMUMtkoGL3NslaQpA+5b1zQ+n9LBf+qbGH80TozG9La+VT4FaPlP0Vam/s4uUPLJJ+YR2y8Osq
U1IZjyZNLt6XWGA/yygRndMQyT6BK71k4Hge2SfbBMJtPgMZv11uF/pDtxcH6A9N33lt2Bg3X2zO
UrQQXHdLz1xS3gb6jzQaPEHV8pI9iOBhsEiwqXyFkRfNn6DwqOxx0jw7MHfydrqR7X/lMLUGL88c
RGYc975IepMSQLd/4Vi9MCgu2YNQZ88RQA9uzpJqFEF8i3bglG0AUHS3Gu2C37Awl2/UTJkaawsk
0UbZFrPLNeG/qaS0bfcLIwImO4JmNc7Pqn0zRZiuyCvNfa9GkdT/1F4y6PufKz7Ec9/CGXJZsmeO
wcwM5hkEthhYCmB8m/nDHF+J6utWdDEWXGmAGw/ksAjwKq54KfKasrwlQa6XYARpyf7oP4qffSIm
ePibYXCZofmadV9lWnDiAf0+TzQI2RwL0KP3bF+wmeHTzIkAuM/JJdJckktfwwF5tdvdpRXuFIpZ
hcOGa4ig9DLbH91O8Q5PJsJuSZvPBxRezcHdCn1ll8RjkdKLncjLIcOxoMONEmFVdufWEvInnFf6
fprrW5i3+SAohVQQqfjYHoqoqjuAzcG1ownxrcYXualPxyLnJ9TV1G7/uZaCvx+j+XUZITSp7uEL
Z0RVmnMnvLeYRAOrwk8Y3dxpUT6+kZ7WpdFBXfHHwEPRNtCZ7CbRE9XNB2l18ZTfX9SWEX+wzUCQ
OLKs8s8zaG+diZczpqMY8Df9lgA/OLs0696F3oJdKV2EzeCvGGzR4QHiP6lec9II0jjvTOtnkKJi
nZL187xCu9glF6xJ/ojReqkdCZ3z6bY5MlADIOgTmc4IZ75bUmp4PJ+9hizbDz5ym6fjXgA5j4kp
dZrQidxiokwf+0pyUKjVFPkYwK9J3DMNG5cNMHX7H/8WJcajTs17OlemR4MsIMMsFsYYGfGxYmO1
SpD1Jwzlwc3pz/FGLBcbDF7Ttr8zO/bf2k4fF64v9vTUMO0ZWr4Nvxl9G1e5O1whOdjEGWh7So+h
yv3i3WzRwY7DFW9oBpv339pjR56N2vxQFKvaPfYs9ubcOKXGSzBdDjFJCHqgZmD9z88JPQSrcQZ8
/OAyEvFndNTGPG7yUGmPEGDP5mq0iBSEoPIyUYYfU+PQYk9nR7WYFBGGz24W9A8t5pYe0CguS9V1
+4Y+ocPpJLa+KvfQOxTu9Tl55J+tJzdg/KDCUy3qjsUSeFaEBKJAWrkbznjzpMtWpcK9yaxQeD+G
n6LKmQx5a/cmmYFMsGeUA3pnPfNDffKtTbWodsLrrcgpQPWw9EGyQ3NSGHDhgC2OjOSptcJXriIY
rrofhXb4MtVJsBlmLQdW8D2tCYiZSR7DMI6oVyD7K2RmV1Y+JEQQzTWsauXmMngYbDNc8CKVXSpo
0R6Vij+Ke7yBCw6S/fbobsar27ov8v8pRotv7YW/vaEHif7MxlSVHaNrJRRC6cctUocaEH9TYx3N
kuI8G38WC1R32RThUU+OoQ+J8UWs8bcMZAn15l6U99rZLPMxAoS00cLOIZdGt+eMC/TIWb2tq1yd
SW2Z/3YKefZFtMeiq75uhP2ThFjzlNlJA5k7T0FQP+kVc519F504SYqaYM6hpR2nVuVmPyAkfEQ1
jBFfLOcmbvlan4cL9DS0FQxGuKBly/WgaZVTZ/iD5pT1gro7VOFUnk1mTXS7I2FiUt/SgOU7W07g
dGGMRYy9iJ7YQb22sfB90yCjVJgWqMswcaNecsNnkjugRsKcNmTzfQTNiAZvNrToHV1S9FKb5uSb
H69d7lkW67oK9+VAJc7gi7Axt8gh7mc/zlk/nuEfEvNKdHMUdCcnhiCH9d9WBb9L8xH3srTsFY0V
aeDQqeOU+4vIBOcW+tcCi89o3eYkWvT3DPLTSaZzWB8EmGibtyE8tWJLNV7nBoD4384EMAYh7iyl
xENLzLbO5Cis4XchXwYr24tVzbqzW9hN18AH1Dz46FeNbIeXnByxALUf/f4OXqfUM6zLfyVoApTi
N5pKkOjbZiICs3LoIR6ldJkhHS5/nxjlZPrKnerymSLMzDNOIncuVKoAL3DRrGWRDH6mK66TZU8Z
vhuDYu72nroOidwixMrAS4GSXxRC1eXhusRs3z55HEMjDI18Bnkgqa7Vv2PFS1ymClsfvwysRl47
iy39SCFApCQHLoMUx8UGS/BDzeZ+u8jzi9nZkUkoHK4FGjmMbKOryk4eJm6KBCfPbl3WExnM0wCL
SoGhr8ZhdLUWPnALe7zlxyFsXGjJu8Vs/G2yY4loTcCr1r7aeFu1162vZQJO7KITaNv1xLNR0kZT
w6YvEGcaEnfm5qjKoTJhUQU4RO6yyD+TY6XzHAv7XXVKSaCV+ksSFvSsBsT5P2SCjv9BWxa3ZwIh
Gyy5RJmzRjIuueDvAt5kOmWc0v6DVfmtReQFwN5Ei8o1QqGhV2fJdfumKVslAJYvew2LChYtBgrC
JcbUL21bAXK6RZ+GPwKp2Qb7dE8xDE+p/Tw7X8FVz0QhBYN1p3vdPzlygCfOwV1NX5zlTjlle3lv
0+3B25HmbuqhoUz2UhJpqKSzkWHPoYsA6ToYyeu9d9USmNxxI5ttHvSFzWnexpVienH76BO65QEV
Csd4KVWHK+Sg/8MeGrxMIDYerKPppYQQBUbxuOYrRdBnMEGtcb8aJYsTbu1zNVVUSkRRD7Bit8EW
MMXgYvB19GZMBN2fkJawZOY2JOsKG+KwDdIxQRyeZ1VSqlDHcNnL9DodTGE1rKbMBETpeKinH9xM
IrizzeazZdSAuVxbpT8aZPfTkAbf5Zb2S7IsJOM3YXgVTOGnXneLDofKOFO9qLmBB1q3pd3w6fIO
XdWmYftDEhT/nqvZqKBDd8hRl/NOIgwSavcSpPIX1JnxWcE/FXAnZbPKo+2E6E55zQo9Jh366YFm
gLCtB3w2gog+S/4yHyRuGwcac0J0nTL6/ej2LN4lJaPtwOZngNI7lgtZQKCbH4qv/mUrqoTCs0qJ
OW7F9x8BE3P+4Y4m2lmguqdE2PePx3HBjCx9Wuu7WCeaxK/TbK/70qaYvZ4SKr52doyDW3ZOg/1d
W7DR3TgKEkFegUY2pKa1Bv0bOVGdaP401nYcSg73r5zWiWI8pyuv2mgIxq0RAkGwOltz543NRFU/
mQyk3kJ3xOEcATcQmqd3NNQuI6hW12brEJre1gN4poBL4W+mfLNiZYZ17bO3j/PNDeBmZlXrp04F
fOQ0/AHLpQuFNs/CNoCWE2r0zen/9j7IsPvgXnsqSCkx9/vPylKTNdl6ZMqhqYFDkDBEeV2p0Vkx
f1wikRSgfkuYJxByMDjksdSJ+CRTrxsi0xy2XTk+TdjZQbYwDv/+4nM451bSZGO0pgj9+zhfCqLb
mMaVfSbY85TH8TvwU2EozVBp8MdQFIn8BGlGBygypUlB5ciCtqjKAWyqwiD0uVFEBS9wetU2ctRo
pnIvePE8NcHnSHkPb2AhdWz6lTqpOvjoP6AM8SH/K8WihTeZJ3AkHanFGdCDzUqBdo/L3bbnVW1/
rMFJO4K6UGGoR+Rww6iJFYJTmsSfVsJPOp61nd8pqEYyGde0eCvxG4K5FKVKhznQWj6N4vCwb8a7
EzCF0z2mSUHFlsynLq5CZoJVH58QsCCiAfnR3DtdDu1Rq8R/AZhN6oSDPMODzk5jrIB5JcEf9z8s
bSQ/9JXoinRL0STQl4y0MheyY9kK0pGnnCgtpTeTGB+F1hw4t2qMoYts32q8qcCYzz0HWLp+e7CG
uyvSey26IHjlfz89ubrbbdwXbIy88TkOZeH8+W30+qBIm1TU4mEpdUNo3uKEvJAufixkg9rGN4dV
dj5u3gOgV0RO/eeX7Yo4zAGpba4q6n4LSRr80gI9XsFJme15SRm9h4PCMcorD7OHeL+60CifZqZU
PfmZbxeh/O7cHQy8QtWisiPShETGqzltVdQ5wrr5FQjdnWZp6C+rnUZDnxOE8Ecot40WnWAZpbgW
s6wsaEFBWR7C5xtnlow79JSSLokp9i/WIxfy3gTOYyO9xz4dVgfO3B2bdmz2uKGtL72Q2ZQYP37P
yF0YIHZz495eW/LH+nOGprcagXMA4A39+8rkZntjPuoYH1OSZmQJVWYJd+x1nA9WMeN6nlA3H41N
5oh29jqm+tpu/SCpPb5vDPAOzrghIXQ+wHSgwla+rwX9oLFRRl3Q0AuP1ZvAU8pa3xuCbvx1S4eB
GOxi4Gc6TkkSUdr7oErDi6QXfZMStCh1ZEbhis33P5NpLRIrRt8NbSZdF/9wBLfXXJ22bBeMwDbh
X3TMT2PxXh/cx0xvh4xE1e1qZt2six3BP7GHAjOPGr2h/+nOAiFQ0YyIkr/bxl+ZQcUOgLDqopph
IaLStSU6ur+HpqEQ7irGSsJ+lMUD/WCuhqCDqjHQbwdECU82GZEc/liLN08fbbivsRP7D73FM8N2
hXzbAnaC0OWCJRyqVtimHqo+tknDgn4fm13zr7WPiv/omdT2eIqvZ+dWWFpBv8OLHw/oLugEkZ9Y
EzK41iHd0CK45lUHBAsf+NK9LB+JLWVlAG5UlaU0yvGc5I+RwCEsu4gPaoC6b0q+mrsi2oxp0c7+
V5hl/8HOjS4L6ryWxm0f2B6sWwunZsTIlryRJ5butpNZKeZDW3x30UdI/I6+HR9H06kthUxoyJ2W
PC7fS05+haHaubwGxxoAtC7pLWMquiKMqiS6Rw++grN0XUEw0Tiqxu52q8R93xnJOa0D2OKZtc26
q0vZqMXeee/WFDNNBZFJMuS5KR+p0bZwZ1zt9MsuATFnbfQsqTlWt3T/bWMavs0jm3QMcbawjFnB
hTVnV9T1BTaUy3N+BXpkW7XV6BDE27wcZKS0WkJ6N/Ns9ekG+uAIZdaoEASINeWk23LH7haC+V9K
xeDQVadBCw7l0PvDUDmCYdssg7gu9gqnOJ/HeznDqSRFnxb1hGSYvCfY7d0bsY5/Zb1mk4V4Nte0
aH2K/jf1ecaWVzb/uY6O81H8X57Ck1NeNHgscrqC4cI3MUY2FeTsV9KoUp4CLpzKNB6bn93X6LPi
57kK7DSofLHj07tCKXJL4UDRQhcF7d9d7a4kyfA32pM9pYRoSsjQIBZChzlmu2spxu2z7lB0pMpj
8XXvh2LT/hVVgDns3QUmreEkLkJpNaxANbGeHl/g403uD2nyasvtLymy+fFhJ/YeZxBRaIkZ3VNP
2bSye+PTpSPwJPsJW9hp1gfjedjFaxRbMZqw/kJHJbBJI6zMKem3UrMHsEge7/qVj+8xpdVnq8pt
fvrw69VfVv/bCIbLDnKy31A2sha9VSl8f3JOa8SuHW/kSbsfq00UcuuddJ2Q/pCEFWy0+/thqKMO
GYskTsk/2Nc8tHW1I0wsgSipR0nC768fIWoHJGklufBP+iUQC8Y5xYZXA2kwYwTR97llMfe6Lwbq
LmUUduCHsHIjaiG7dHc4abIrBc78iu1pTh5aPrMkinMLYa1xJfMtbzHnK4P33YLdciuCumbfZbrp
2/yAHsZFkZWJjVYoAl77V/EB60RWx3RaJwwPUQl9t/ZeX1fTKYzfYOQmnvyAVzbat+fmjY+aqKEu
H7i4n+NuQGGyXy6Bst/tc4lXuGLWKkUXXBfgYLmu23MfS2Z+fXkxBdZvhc59wcmr+blP76qroLAr
qiRyYcYCkzfSOkh/R/6IIUBAv5vWUjaaVrxop6JZ6pLtxGe/rwMg9lCT3ZUFI6FPIKCGO+sE9URY
QyZ6f3bo0wajtH88I5PwEiTZQD8dWTWjc6AXqu96LLeZ9/aeo1YzvUG0H7dLRcrtCcNkZe+B6K8h
JCvrnVAWNoJcDdrV4VqteMk2kmtfF8PUuuFDdzxh/cZckJbXajv+VpkpVbO56kAsFHwabdRr26u4
GiNJnoREzjoeKqwn/oXj3hnE4XYMOWpcQtla4TAuJQuartlaVNmCdy/uMCQsK+7PffA3Qd8RhffS
+Awbs5jJeElsCTzdzUvuDg4QECwsHyAyBLPyKxwOBbpyt8nRbB5urZr4NlHtyuv3O2EJKCH9iOU2
46uYlxgOQBPOrkA26OWU50XHT9NZUL/XUXAefe4QDXarYwbHDYQEhWUqqbbDfwyxb5JP3QPaUJ2d
E6LN3fo/l5Bab+EdZrPN8/Wm7Io5LqMdXFIp39tdsaAw4wdis/nqYb2XMqSPiXjtH7JtHVDNa/b4
AjR8B2k96EyrEduUf/8DTk7TL+v421rxMyz/FKtlbZ/L69Oe1k2nX1dKluKHoANRLuS5/+bmYBhm
/emzQIV6NbV6QMiGjoYJFvArrAsS3X5+7zz+HP4aMJYqhCyrb2ZmYPvXXrLT4brzN++xHq/X/hH0
lB1FIBhpTDnGfnsKOCNo7ROSGUHFFTNyMlEpuM6BtOpyoBNqZQnogicYk2kc+nr0K+NcGDp4IFXL
hiMV5+9BjoaAUHLBhwNsFKM6PNg/eOC+VNuMDCnY6MOgk6MpmIvbN/MZWMWIzcyxWcO6zyMRkY09
vZ/F5W4zrS7IhnxgjuUe7YEwGy5f8Fu0jrqUJfpJx3RjUytLTyFO58RnR0kxp2PPXzZd6H+/p9oa
SCZ03Kv6OeBz7pCFdjZS46dGPs5QxNM3lEttGuoKzcp5M+kGVYFXotmVz1GgWPzP09AqE92YmeTk
gWbCSMm8k+cR9uRF7UL8rK6/pWAeh3ECo5/jJVJdNxH0MCkX08H/snlpF0C1N6b6eGLYSTIDyzUM
l58US0AYaGT5QqHe/5u3nbt48cfKVMDwN6h/OGgWc1/GUj19losv/xkeIL0/sQzOtxavx48mQ/Pg
UnUPji2iV+DbKbbxIvUuUlQC50kBE7vAPNgPegg1DzAWGgNm4LoQHq/OlCjENS6O4PmqRf1/61T8
nMRWcZ+9n96zjswI7ihLUJpPkMVdMRdrpfUYcn6xrFkXt1MtZDot2mYJ1CesRaAY1/QLZU8o++Va
2zQSDAiiYzQP6XaX00t5HEtXNzgYql40fnxOOBJS0bdz+/v16egYSgzHio48CK02K+nDV/9dPVU4
CA8oRm/9rgpEN4UzzPeARJ6DGrpnVruvIquQmovoXJmEvDLp50n9G18LOLUV45BZRPLQN8xlJVc2
l/EoVHisGFpRiCs2WbtooE+2XrIydZsaHck1iBNxmq0OHA9VeYVC12o84igx7GltuuvJZVu92kWV
m5/acOOVhJHr42CLl5CB+FmDiWPj4AjOnxDRM/SrsBY/M+0xV4nau3F2xPe50PNh1ufHR7W7UEp6
JzCJS+Hwi6hBQT4lpPG9i8HLpK2SqZmSR1/HkhXpMnT8dI6ReuISsE9yoVqtYs6tc6OaB8we0Pvp
TN40fcv25t3ar4wyF6XrvIIfbtIpfs3HDsbrFVgzt8DSk0CMNYsYQW/Yg4s8BLmBVnqrRburuOfX
MqEkGJxsybxGazWrdyRQqlcTplusTuLrEeWvicL1bk9u07gmnGMEGhT1Gp4qF7BkUZ2gaSwQVoaQ
iyhB1Q10IGl1N4r+Pc+hvG9MTZO9Uz7l9YAXg+HzdABBRLXopQ26+0XJt3Dwayyb5w99cJk8kyyZ
KmE2l6pIoPvO2rq45xzxxu1OfO7mNgFDsxk+rELQ77rgW8SD9jv+wg+ItajpGASmW5IfDYutucho
shD8M8fUnERZRgfMRGpHyP+rLRwXXeyHuVil+pm/iMSof4BtdAncUdBZQLp/8SW2xho2Kfyc5Crd
76e5rMW+IHdtEW31c1HJknqzt+Rp2zl+GYeUNH2dlXXLs+9Fow6qb154LWz9nMRo6uH4eb1WPZat
MksGXYhs8C5KEYvsaqPHgLntmIaYWG+318ixba/Rbz4ts//ekvkFYiCSXhwemd5BWAqLqHAruPOt
XhfgTF6bS123USKoHbbSTOhhkuPYrWb3f65K6xt9Pks1c++rKvei/f66loRpLnK5UGhfFAm1A882
+2cxq5Pg81Pgue5TfsR8paWH4mumsLN8yBVsTBLhw2x7vcqLgkbZ4ltlP/7JSCy+MKNXjeb6bFlc
4yysF2zjVc1UVuk8GhLoQVoiZxE6hAVYd1BagQEOOm/DtP6hPoiKH4UX4ZpYvLkCoASTpPAnQY6P
/2JrKOiVYkdWEL9X95k7Nk0d+xwAGGfbxYFohK00DqBOnp6Ki+ip9QT4aauK7sP0vqZWflMHpyzJ
FTDPoDBwfQmFTUlvew4pN/pqbqZUlsYZBKg5kaE2BgFDdg31LoPiCS1RpH6FXboOk0vnhGLR1WMH
7x253dpdil5j5wF47MH50lmXpEMa1+h13UKc8kcrKPTUESOdbY95jR/q343F5K/m4eWbrYpYqFH8
CZic43ZG8AA4kcBi/PqCfaP1XwxhX2wLoE8cCsM86kPxqTmX8PFh/SlEmML5Cv5MCwo3o3c4jVir
Y2PqEGHhshUrIuTb7oyKXZLnMp5sKc9GAromF5wwN/t9P3aC+fME8MhMXZYLGLX5J4lYIwzV0P/M
vBlE8T5RHIzOX4vdk9ku4YTPOR04QqbyWVJPjBDSSo+qkHAxQA3likfnucgkZm/atqwqZjstO9Sr
O5xiaNS51RyZmW37o/srpEGUX7SsFHccIPAfU8VUHCIoZZbc2KPPrZ4QpZLpJ31IsmhXzuhIlfDb
gtytDxZ7msKwYkR09Wvj25RVPQplORWk0B1WGLYmeJldYs/XcCtNGyllXNUQmQTicsJuKFaxuLSY
fK2r9ydcUsHPRPq9JbbMmlk+WDkA4RLs00nlJlMSarKD4PIA27r21X857wpG+zxcO59kr8S6aAma
m+KP97g91SvHn/7gsontVr+SX5XGWHu/z7CFb2+ZjGBUViQhzXtnNlcASDfmYMYHSO51xw8kzuhC
5IuoHIbegFNLAwZDSbw1m29X/OxdHL5krImQVoENF9DqBRdvDsM8zGJ500gW2BTthPSbP0jyipb9
LpUl9ZmC6bwZY4h7mBevO/HwEN0drcTZxJTpyvh1gs4JIS5tBoUKh2qtac5JZ9gswu1aO+fYru4E
XZPHgGkV1UTgiwePixq/rT3Hd4PFuwlDXs9c6WSLE+uYADtXnMWM0ZFBfX/9N5kUeJrdpPvI/NkH
ITaS4Iq3S+j8nF3+hMl598QWzcJZ+y4c/B9xQaDmZglprXUocdq409fBRoEoXkVKvUGRYGAXbbEY
axGfzBzNpzRXWWmNZ8ihre8cJPJSmCvunlFZPIhczhPrnFuTv2KzacUrU6jPqoDqk0ApW+jyBVy3
AOD9Mt9PZalH/VdyUhPc26k4h4C58GCfDfv0mge+nd8ADLB+PwYTXYzLM2feQdM2w8p6tf/3JDlk
TLWc1KiolLhd8okPXizYUBjxsdTHcICSK55kYT1AIZP3IP2M7u3IrLhDfLq/NaQgc6rK6E/8mfar
73JALat2dPi1XZVupe0cCIPbi7x78YxW02A+LcVsqmz/9SNhsYgDksDC9mxeAOYiunzJU0lELixO
hP3lB1I6+V3x5nWd05xJI8W/qTfxmTVCQfX64KII3JCWRbE/CTuQyFk9Y5t6GziJO7OUGI4kwC/j
+DnVEkKiZ+6g0kST2YKxy4Y7l7yMx8fojCdKhsn7yIJOpnLpiPUu+B7MvCjsmCi3nwOZPTB+4zuP
E30/1Y32J+KK5zMlq4iuqG7IvYmyd02XAnmoD1FS36/4F43bIlMAx22XNV7R0fwjFJv4ujt7IGTj
bwA2Jod+LVjmdddwurK/nRJIjep38A17Ol+mc2ciuTJSTjojBDzVamsVHpcEWakXFHn5/CWVny7H
JREJ1BZ7Lf9fxSh7qKLoK6PUntt3ccYllIoyhjpt8k87dMy8C0TEJxvjwd6avqLT/ttnU/ab9xhx
9YAvWyXbJr/2Y9bJ3mfEOO3wkgFk1NHBppVPhjzEXj5SeVoi79wwwVOtqWM2Fd5Y2jza4mMQNVz1
S2eKmxoP/JOnZxuUCMQUn3AQ/chK2ep1hM3PElwcmAYgxD9QyKSNkmpjfdi5wiM7axuXhlkc+0yj
qdd7J8/YmOh1kt3MVu92bo9oONYFGn3wGtxQ2YGXKW/P3j4wBV+tKOYPiLPhtFivSdDFkrNrSDmn
0VN6fhyCCjFyL+0gngr5RAFbrNww/O6kPHRY5sDbdykIytX56Gg1rsC6cEqHIxJCCPBvZovvJqCP
7hIHw69xfl7R0XaKVWYGddaoOSI9zslZNjTS1hINHSRimFiBtl3jv16Q0CGl4nYZ0qRcxiwAVvTH
n9G/z8Bm6Ttro5ZgSZ/jVmKUSRTftdse7ift6b3ZFEpm6D3UoY5BSSnVjyRflmcZqAcrglfwbIwE
SqERQVY9i1Lp/k6+aVmDb0UOCz6urI6y9IKK1IQPNDF+P66oBpPgjQE8hEerwv76HFOw7K0iddHD
sSpKHCkauUrX1II8EQHg5z5Tqanjp0r+U+IVeo/DtKo35Uz1BOzL6iV9ETJ6M5oy3yaAvqZsW1K4
pfYNuPw629KfAUUe8EhqzDPUM5EVVdlN0ofWT5wVRTys5AP48sxp9CnypnUfAWfEv/fobHs/NUbD
n9ijY8MCaiSSkc8R2wxNgRG/f/jbzXMWcq0uIzCWzL2H5MzPUNfgEpKOMHKKGWomCxhinpPOIno5
ElQfCu7P8Gul+DOjwvayDgbOwWAaWOrnAEdA0BGW0fw0KOPAENKu+3LKsK431LzteJWgiMgOvjlZ
yY6SJZAr+S8NYwNDObKb4G5gPDf0liTvhH9/3F89aevfDSyvCPgENIeM/0OEIrryQTHN0vwJTzVP
76oypxxHhW93JIuD53I8mvlLDvC7teRhn0uk0+buoasHAtFyz0oSqJ17sIAS7abIsQpRb0J6Aiya
bSzX/Q2b9fxHOOjh90ldjf56XuJtPFsZmM5zoUSK8YWSRkmUaJKkunZ6YrOFhSHwkA8vFTXz+yjC
Z2BcD60vozquNB0X3mLdCD0BsPA351Ce4Sp/gnobmvEKGwNuplD/hQpKTuw74P5+4qqPz2qVoWVQ
SgU4k7wIZRSSJmbQxnnRtpy5LXOI2plXE3XOueUPkoOYZgouPjGc8hsYG+08IOsRALjVOWTVEPxB
V1LJXi5EpwhN3TYodAHVYBpKfDhQIlLKaIEfiJdBd/vnSdiEiPotfsP5bt2YKfT/vTilUffiV7A/
vkrrIzTO2l0ebleEUi6vnLryXJolUJRJcVmybCdwH1Wsg8c8jtB4HTcgeahTgvWZaZlS+zPvmoCw
kEqnGy5oXgKiPKXO/tOy1+lPiGG2fa28JGff+o2A2r3c2JXf2ycZSHYdioeZrYaOTHUa2M1guRCb
UCgSjS9unqFiIOEqbNKw7cMpLhd8C2gFvqkWjkGYGvSrZaJ4Vn/3tk6FHfGIq69vRO+KNPFUK1D6
SvTxB2gqkKQIEPcfZxRpftHzAeeiCIoJ8+lFM3j07wO3kP6OiPqd6OS9YFCz15p39H3dXyIlHj9G
GRX9lcbIVpIXy+6tSQAjj6aZRqWdF6CbZsA+E7/Ae4g68vfuqzrA38D9bu2BNzqJEKdisE+CibyI
X5ThoNFH0spPfbkC+r+ZDUO4fkuhctV+4CroTY+QwXyr3GrE7fSzWbMZHwFzn8xQ/vZEOIaKhRyB
nvfBgcuVi9H7gsVHfBL4KjnC0eUl2Q3Bm9VSzwXVDKuluXvXDA8V+bZxqinsRtSJPpwU/GA9uTVY
GHoTxXljfsaTcyUiAxwju4v0lxMmo/Tk3je8tPJnYnvwnyn2aPuJKh/QUK9yU0itctQLQBo5WL+D
uNG9RjxzuiHap0fCh/Sfrb4ri57dSNeDzpENGgakCINomLiQboSitRCDAvX7/VzOPcqKSQrXor6T
1mrsxHLjhU/DY5DlvPX0FgKTRRTJAS5h4/4Y0O/N46imoDIrbrEBYw/oQZcb3lV/0TpA5VcMPlU1
7E5HaqdmVT7/ytjQIq9JYbVSJNkLqyNx7TnFP/CgTcT9C9wrryCqB8JdjdfdgeZfMpmtgV8Pczw3
mDfUou9iTg77KFnYezSGKfsGum2f1zAvwFQigGOMw1FOXJWxGSDF8ARFDPZntBaX6hWmMGIF5sLD
bH/Zl2sv6V53AqWxZwEghFz9+eBlDICDe1tTcoVPxWKj/1J02mpgd2puOhlnGOBahLdpFVeZ9za2
tM4OPpTS6GRymAMkcMTtTTlZZSJhX011Kgj/gjttRp6inypD8xjCGDmWcy2KUUN4fQxkbMaBvKes
7T9dkUtoQitmdOcYSYvIua0eiJ+yDD28DzrCumnMDZ+6CAzkS7g+YMxyVnqrdPcBCIxCVl5S7WGd
D+pip0DFG2p5iPDQZXTeV/8OhQ99nGM4+P7VjN3X9vg4TFbdr3YAHv2B9roVdMQJaSVn4wwDDODa
wBB5XUp/XQ1X5Bm2k4Ss/a/KLh6Kwn/z+7a2iOyW3uWQZ2Xtd2qrfnKmcmgCsomR1kRnu1Fvgbfe
JLA6OWT6+xRRvYT9cXf8qHCnZyCvjsNyOkg8VKaGrMuPBWJKmtJBPxlzvJab19iTDttyeSr+IYUN
CLD8hpTKXylR0/UiNQ445RpJaGv3VpY99xrTqeSynovj7GPuSB4E/M+5AOS7x7ZqNaeiBKYu/pQ1
yPogcoeCmoLnMT6SP21UB7q9FiI97UcOwXn3FPXQX5Vu67c20Ew17o1vZHWVenDFWXBBzgxugA+h
47Hyj+6O8zgWsN16j6tu7z4NrEyYosjADhN1Bvmj7oscv97OhoD8Xi7gP7DSgGwfGKVeWRGZc/rv
Ps0pXVJ7el6oLqvStl9PsyS0kfbq1CLB3Q0/H5YPo5Xyy6M6xLZjDjE8shmNAx1dhQYAL9zz/WW1
Uwm1Qq42tYbNGFGAORbvE96iPn5+E+/hrBy3aNcTQ/kJWuOg2eq22i/Ddxu3nJI8eC/WC8KS6SIh
r45scQaaC9CALQIJiWtDo/m0SvhBQZuKumWSJZXdD0CW+uWVXBvFoNCIVqalvBxDwqfCwpcNNo/G
n8MaRNCpkQ+jl0s6Y92etB8C8c3SOVivB1IrNEBiuOjRCRNOAxokwYQoFHUhUFvgK9lVjw9zm5up
HM458datvvSImlhumMKtsG1DsIg1ATM4OZ6sn8pdx0fYyJwTYw+klyZclfbptYRHny496zYU35cz
PQ448BCrNupcm1JBogJLT+IbNg2amK683gBlkbcbK/4dwGpXx0abqRijoraqweFct2KkjrFVueJb
NEVSQdbaZ2Pf1cgl0YK/hKESSQwYqR3VOBjbz9VF1guTrSq6sygAk4EE5xOK34WVwBpAqApcFeMN
sfqevvzD5N/JqamOgn1J+sYAY8DXFQb2G2SUoGrKWyF76LMKpvRFow/HsEC1To2gYB9Perli2rh0
wOAYu57gKZVAHMstmwVmNu+lRNOEK4AK1l+XXKIlZ2a0TLL7OT1T+p5dyoEFFWn0yWixvC78uzyN
RSLihw4GpKOop4OBc3IQ4gLykQqlXgWWbiWK9N+Pl7qHw7/Y28NvpgMvg2NanIbSsSO7V68eqbll
EA7sz5QFPM9pyYhfMqtgxie9W2uByRvP6leyf2PUGeUEU0s18cycvaj2OGgKByjkXtUiI+fCMO0w
1vLUhkyXqAM7PAuhvpEyzQGwqmoNuGV7+FAF60SgAGFYerZWSuqbxm27YIGV9HcTzuEI/52ncAzc
18vxKGShjaebhXcGHkJn8XmOD6Buu8D8NpykqXuUkERd0Q2cnqgx8f79pw2a8do6phMv+fBkD68C
taVEjfoygv6cf0mTAfDVbIgrV0PIuMEmtV6PU7+U9B1FxUxpdLf842Kcim96Rd2gWuMGnWlgYc/7
7AkeA4WyE8AerqaUarvDlFwmCPysFSdORmsuZ9V4sCwrSVYF6QnkPi6VxN7rutZyzllzFRpDJPkd
00UmNp1fh12auzeZKTXHStB1sdu872zZ47MLy+J3VUJS4oTzRa1NOgkROEBg1JZ0eEp/8KOpj+ea
fEjEpXy6CGKVsglqKGZG9O7Ym2zlXqvTd1ink6xGL0TJ/iCCvYmACJVMuKOYaJCMIP81aXRCeWsi
NezmE5Iwq0ybqkdqVhiZEoglUQum/UQuzVUVjGHfYvGB2VLL5bEiH05nZKTRvSxLAFehAMiY7epj
hPXtx0/RgYXD24vbn4EGbaDoJUCmlKL9eFGvMnVOpn0k0zdWQ+NZOtYaO4P4gjcw+jp1DiquS/uB
1E3LN6yMxdOI9M++GnzU1GWzHQID5Kfz5Hdm20J2lK8BLjxxYsJkPP5iHWWHo7VX7UcfrCsvr7zR
IeBNaDvzqIlf8flWSCCbqQx5Z38eE7XyujIhXdoyt0ckIEsTFNDGZNtugjODVrPOdJLGqBuTqUOJ
redtpZuFd5V/7yb9R/r0XfDq/xtjP/kiypo2mT9HrfQGaroyYFItPbaowkK2W3D2GLjbRMc4OmV3
o1YhLzW6h85/FM6Mw053c6aG7+aq6qNNDPLKe6UPkV5VJjEVrLdmKfIgimUmSo4A/U8fsjaxnOq4
exP3TB/ymtfKrvBay/0ljwQ41xWUqFPGxRNUXmriH4tDDCygGh18IkVVVykT4TOzYndZvS+9Vlcq
m4muhFUGUFIaNtk/o13+eiXE0EXPwjwob/WfNWI09KAKd0VK/ryL0XH8WCMQqHv3OTMlpN2LC0Y2
wqezAdXUx1PJbqcSNZi75b13IMjECKUOfUCR916TQrjCyq9FAQLVC3Gn0Vunja4cojZGUUCAXwlZ
Ro8dDkdFumV0MOWIAyjh6o/WS2OhFhdDJ/eAj5xUG+wzT9POZ1C4eHZphdnoZsOCNkFNl7ZxMpmL
2k0mxF8dsF2wCtXsCyi5DBn3G8DOl/TZA6Oifon3x3scCKrEtZRundkAYKiAqkgi6g243W0LBrsm
LvD1Q3N7pPZbRZjQrWQqI1c1KkYzBgH/ELH4cB8M5d+ruchRm2Hl+wSUXYoZymSb3e95kZqvi92z
9K0+NsUveuNb0pc60Pbhkf/fO2mTT4nu9+EL0gAxxqVrNn2eokfHmEnhxhtsz9ju2LUFfPFVQD8Z
rUvgF3Pwyo1bFa4ipAq7ihSQSsRf8EioXpOs/7YWrnRoBXS8Eg4U2SriPL7j+Gy1FjpeGwtU2HI7
VcfU5Fx3nhNbVV6H34zKwLiJnTSvzFYoJnaPUD2MGho/Tn3cXkyuh7dkmW+k0s5Sevg02ibaEV97
mxDhyPwiKjqMppAKcf7IUvoSRxnnw+USN5SU1XcscBWHGUYm6ZqxU+xVz3VvrY4kEBemjtOyBMA+
eXS78/4Qs97NZbd55Bg3DI9YJB2AdHb9p+CkJYhhxMh0J+e4YitBIZhyuZhznXjms0k+C8Y53xmj
lR6w0PPTL1+a71BYNIoezvgDtFHEA727V4f3o10l06PdeAHihwvgAexkMviTzz8e3AfheIDja4Wm
bB3Wrjd//O1Gs97/QE8emqI1g4wK6L+YjB/EMsoLzeJomptKG2ZP2sdpz0EiXbZIL2u9JtScnERj
1V3vpjxGnZ/jTmT8z7LbymBFYNIMGk1FqqLxzxdBjoWDvmWCciBwuG/jilXkHHt+pqGKht++ONCl
JTer2TvfZ0msbvELmwkaqOVOlA4wpBptfX/DMtHzT1HQf4l9K/kmhtG3vSgukOqByFS2P3iRn/Jd
uNPaI/j31Dr7u70HcD+ZHaLIx+BRpsXjxjjgRlN7HAPyf6vvcumBcxm2tdUDM8vRONf9xGh6nWla
MOJcoSfPviV4DndBlYSCfwz/OS5CQ3ZZ8gIfXPe9ufAY41QbK6tq31kTakBHh1MmH9KYdP1yAo12
CqGgipOAf26ixRfQGUY1Ec0KFglVqCvlrQs84iKTJNpVi+Du7pGCmN5inzrmnxKIMVxqQiptXglF
K6EzeTwGNhCNsxmK9BRfB7DtX9eTamrbNQY+ASEAyuqdURLjkJGqTzAwumsBHGfkQhij71Jt8F/D
nkqme3q7KUygsTg2nYaV6b8REGbe24ioG46ydt9H+h4AnsqHLTFIhRXZzcQCKPeqnCF5Hgz5AHd7
uJ1KdIT0fExFaV5mvyYEJoGWUvDAKsmbCpK9FGxm7SrZIxgVc5xORy/a4pngHd1sEwql5oYdGxtg
2ueZyRZV9NSl9jClNCpm4itkYZ5syWbXRzLwOp4+MEsE3LovwodM6Khx324Xi63w4noYjAZl+glL
YRXA55iyFJhJCNgCpQmAGLcFyHNMprx8wpTo23vNc8rtBEi1uuaiQxAlib+PMFycvszv0oKLv8Ps
+/ZIFZ2DL2qZ1BRqSVTwJojuRAzH4EUkSma+jtRaD79jYhvIMmXKhNJ7U2dBzPF4pxidA+G8BzSf
0Vs6rFMYDdVYVY1S8eSwznzDmaaodt0vnHRnt62fc4klps2gKa9yz48ZkZDNsMciVCa63Pk3MNeI
+3ok0L3L/cjSv8wr9IYTlP87xUgJUrx6VEzWE3vJQSLPPMK5k2hS2FfHdfkeUBftDdND8mez5gIb
E6vEoTErW/iiSHBWw3EaSAq9FLagKcH80r2tuR7XuJLxG2qLMWWlKq3YN5DweDQ+XvkJG9Vd0IFT
YYIjAnVHyBMbpymIgQVkXJUMBoIQyWMsfZgr/4mtchm26fImvcq1AqT4VDRL3oB/vwZpD0K6ByS3
Vgm93CMxQ7LD3jiV5aDadnKccQHJ5b6ziy6ntQF5yJEt0ytsdKJ6sIjjVDqFFd4U46e0kNF4C/1X
s9qfp7j859C1a4EWLRfG4Xp+vHuiOUjkLcTYVXgNHG1Uf1iVjm6ZQU2vq37XUCZGSsTQt8TC+GsF
IlVXkPODD8GhToDms7pfQ/tzTBPldDLpHJySCS/UTngzhxMjNJinKuQjnYosFyTkkaL37o4fyIre
3VktQJ+wHlTV5GXVWUrNIqPl21YRYulX9beHA8b+ZCZHsDMTZosg8W1PkK40RAdfG8xthGrUkXJz
AbqhgYum+zuSZdezlJbiy9tI0qc7jbsoAU+pjurfbC1qWDwLmsQ7Cub+ohujSGdlSsHKmrC+JFxs
Mn93ycVxUOra4v2hJZ6YP4SdGZ0elX1K8sF6UBpQeu/w/7tM4s9Q7oowluzsdoYw7AWLvQqaevmL
C3+pliXWwyU5oNNWBT+RUb7uwpufxYXIAV2unQ0gEYJ18I1yOueaqrv6RMBb/79Hzsle5g05eVgD
pXxm9tnp/QSJbslW15f3YEVWDiYCmZwfCwwzN5wulDGkhKVYE5hsB5bKWkMGm81EjjQ1KI2zKQxC
LSPGK+ouCM1OnEUgdBcJ7+pnxEohWRzGmLQbqVE/3oGkIYWDBP5525ESB0TqnqLudS/BoY5RzncE
A+YgCIzZdYbBWr084qyfMzXPa0poLvIjc+XocgkV1X3Z7bzhDJqWxeisD5Lv10Zx+p+5oENDg3oF
piRdhRNI8bdNMrPi+YksXDDsS30w1r8bJ+srZUzmBuAfnN8xsIY2vWcmVygfQvEwSiLCJFBOnsBf
TQ5uz0v1WAppX4tDZXv9gosC4wADs/KV/OwY8GWeSbjT5oowbCTh1MJxPu1eLVZQ34V8NpwVg1IO
DM5tkFlCCwvgv/Z1e1KGDrobO/2m1xFUUHzXIquTGBWk6U9InG0kMVZMTyN86G7oZKYNpMbCQI62
A7dJVcEuYD638UVcXBcd3RTDgpF16ocPWOgE77Kq1ITo4MeOF/h9WlI5e7CZxvsvRu+IunLr28Uf
yO4bDj/AGOzE2tGD9ZFNpaCgtECtb2y66qHf4kyrerW5JD44TWz3e7psJ3biihKCDec4dj3pq6nO
IJoHnXliCk1/UK6Wq7QMeZaWs2Vo4DNWKuV5vL2FHLONSmEk0hoCqnT0i+h9ki1r6ZJCmk1jmpI9
kKrXE8IQ51XVUlHCvi5WAs3Qy40sfIdGAHoxGSIpViJ7npRS32H9Kx2S1o6A2VJBV8HDrZ+mkdAs
LfdVMzmoAycEyxfYy4e2BoHnTU0Zz8wKSq11w4cIbzR0vopwtSQc22EpDv5vY5Thh1YNGSkjs86y
3yYYFkQXsvBR5DcXcbOrOLh2t3F3FOeQs6N7hIGDPf/TcjIH3M803IOOoxi2nS124MYCCiArP8z9
2XlA7FvZwD2+T6YAUeu6qJJ69m6lCzjaXEXknWUQAK+GlNclQlMapzSB1/OhKbHIcU06bCfjYQMT
XqXItsP2G/DhcFNyqIqk4cz7vLuVnAG91nRzhxkx0Ta3VGU8dQqXWDGvtdu8AHG9R4GxOoL/ZVAF
yAS4PBxMJ83QLDjGYifS41yV5oZK2BOhyAQ5XCQpYusy95kIzKv9mV+piUgBmN9nlw+Bwy8qTd4B
ri0RK+4XqN7RIgqggbZPxh9E1jcgCPiCJr8vM7QDm/hcVJBitV6KvfjOruftVpKOVZ3FBdoXzcD2
4feqBC4GvtRPw0V+WT9ascAaGCnW/AvATGyrhVUAt9Ff47VtNNgOproGYq8RE1R/B3t0xR6hmyaF
e1CSvC9Prxz+LJoevdFwBGHH03ns2jLkbPv7X+0XonvuPF1On5+NLDRzVFbgKXTosLHmcwq+86x7
OPGtXAQS4N97iekLC7/+1QryljeC/k1Vf4HYNuaRdHOP4Jw5cQ2Rl8+Wk5DLV76btV7J8yeRB16v
0TTqLBzhI6seO33GuraXW4kyrrsirT1FertnZNX82XfLuhKH/dIWXEYnQVYii368FCLXyhVVtIdA
IqzPnu9MG9y36mwwAXolReFUV5I1y6D6b9TFUCzUWh/me5pTdELPEoSG4qZCZCEXmSkBCU8MZI13
TD6RtixkP+sdR2BuvmvbRupq3FX1E29HPguMTAunzU5OEFPwm9wcIi6ay6sJZUl5H7GTD4XSJOIm
eVQmXCu7boz2/3AyoTnwW2+E1iUvNVoDB+QC1RoW936+yh9g08dovPWN0BhbJav4BI5i/hQajP1F
ONpFCGwhSnu+lk2vXyWqCcufEAK+hjObZOYHvaDNgSnoq5nuBcoFUJi4SZl69HIAdpxErLZ68RVb
4TFvAmj+4MtC9+GhSulPrIp+NjeaemSyCY5dLAarQnlGCD4agrvc7frWF4LKopBWXVtk9jRsIiZ8
HecU8wWaMCHLPf3yg1MAqGCx1NMyIE8fAxuwGAe0yTYlN9mUM5jK9dFSGsFMt6PZHllVSD51Nw0H
U/dE5EDaUjbKGZ0xE2+2oqrD6d3emsctjBEz6PNz6n7sVuuWqadLlueDG0Kdu4gnFsiBgX/jLJRN
XcVRcIu+M4y1tka1CWJHPd0LsWP8s6JvB2uznp2n/OyVRQK7rCQ8jB4O10d4VxccuBdeB9Gpw2r5
q8S6v85yzt/5K4VD+sHbxvpE6u8mttFEGGR9D/wVuKUBLoJHOb1I6kGwKlFZHTim7M1byFsRg8cq
r7wKR15mbmOjfec56MkDvI2b7A7Apmf19b1riJ1ymE/BnWc3KayDjqaP0hU+Zcxm5/ah9trA8TM/
n+HCvk2kh26ox2QJqH3S1lVuvo8FVg1JFk58fLnvvEjlj1GDE93YXCvHg0qFVoyxKOGg8Na2oI7E
AtNICl2+Aa+CMuUbGV0GBxivdCEPZEnpasTGlqQfqXabiNHjpuyIImcTE00v3qVCzndqrjw3Ofay
6My1FGDTbLDwOmqfNqGpBor3+RqCkYwxToG1ZA6DUKJ54/GAvgZoMWbrD4XjG4D/g/M5AyiyIW8y
xUDyKAz6TNiFEsrC3e4ucVBbqzTZUhOR1TvRWM+65KatqJ4wYMjD591JHzn4b4Sl48nDwYFUNb30
0z84w3b5P3eoB6N6/BiyCZ2JRKUeGxUSoykZWawnlRxJ1tkQkO33l8sxuPdzs3oleTL3WO+m/TFe
ToqQcT3eCSR0fUi0iK6xOpcLIJ3zAhz/Va0LF3HnlCSZ18yCqQLQMeDooFW/jN+qj0CSa/WrOmVq
k+pk7OCBDKSpAx4WyTqmhDfnElynAKtwofTGWQyn6VcAdEJCGiCp8l4nOnOwd5FStxHJSBYKR5Eo
KbGHaYc9WaV5Q8Y4QQRMpTWrQW7WPn5lCns7isAGhMO9jpgC2ifILbGW2Kv/+VzFq6WsL9f0rVuf
+lG1O+kYu2w3dJ5G0lDXlbGWHwVDX+Th9uJXPceOFoaOfmA+xMaKwMx5IIk36f8tOKvbBUT8m0aF
DV7ZT65GRX3XTWyUROg7U/GblX+g2DQQgLXVfpIN3NJA6lbCwr8HqSsmlWhg6eYJY10+UtVH9Abu
/WW8F6ycn9BR76CEpc7b0GkFHmHB6gGVLKY/d7wm5E4kzak0eP1RTlucSGch7wTE+Ep2fDi0JP9N
SEf3vi3b/Qf6O+2uZg3rXumEEW7lQFyHOPr0uQwdfGa82icrovBArpbXUWb0NvWBiSj4iF/BORqE
+TJNuhUqpinVKVUPB+/qU0PKl1prC0M1gzH5+b+R2d66u0Nwvm8LRcLnWWtRvguL03uZUUtr/hF1
6iZJAKGjSzmkEFggpY/f/hsIXu7K0yHuKVxv5Ht5UjMktIgxwdr0wo7GCgQByfYPopgOT1heY8KV
iq4VUAudAiV3UO/KkoazNDcm95XMWFu+lEYzIvTuPsTV59cljwfjZjzU4iopVfePSQuiEy9mpLtD
NtR83Vp959FeziHZx93T/dx6yNflNmJqXabQObR30gQFKFBLUH41aYQJ0WWqj37amKQToUhP4M4m
aB8nLem4CJe3uQlMGkVIOgdzd3752CLh3DDTCG3kglSGXDR0w1RXRUwvQNGimRSsX2z87XQ/IpLu
vIKCiWhexumG+DbBgJpA7iODukvm9cl4rRYHfk19e8SCYJFWJWrqTgrSh8dVKRDtE2xLzcAOpBau
k19wJKhsmT0tNl5HfqsZfsJfYFtZih0hD92jej9uISSg94taV3myj6S5EDGkwcOZhTgrEqd9EByn
5hRoKfXPtWc9Hev1ZkWQKNvN+U4cJ4rDiGhV1uhVjRwxiyBMy/qrUmaaYr3MVohBthI7WQZ30j4e
On6tswIr70tYGnZfjp4OJi56DTpXEGLMRz4bPAv60skdmF+mj316dKGubvaj7QuKN6e3Hzlf6AXg
0mx+sNbWb3W0ftRYp4Utb0pgA1N6RbPKHsEHm9Y5iCrURXLIuZgbJwkNxlfZ1KHdyaJZkxUL/LFF
pLT6d1AYW8U7NtLqhKxAkEFN6kmb8znacDAhNwFp9F2q21JHgdFjNMo8BP7f4DrOw2LxzFuJQ2Nq
6BdVeh3qtLVnqRy/BLLxgYnuUZTw+ydA45prd3twpEycY9q3hMN+0Uz4eZ6DFaGZ6FrnznFLvV+5
w6vYnsVpEvsAm+ghKCLo5L3JEk/Ih51X1t/u/6WKCCu8juUl2ez/fowSVUHEnT0dXGG4/fQlPZ/5
BUpkgTRJqdx/Sqx3JiO69k4kVsvsriWj/2Eqhrk/SHU+dTl9iTXa6QEJy5hZLJ17J5Vnc4J+j2uM
Mfx6xdi2kG5MwmwZoIiEGBN3zJYssQkI8D+geMPR5IVN7L53FGSblCqj8scSzDUWxwn3mYQif3ZN
oROlRihRX4xWacgMY7K760dmRHMN0gOZHvU96X5fYjy8lpm4VtGn/WHBSzK9jjtnq7HRxV7yMJZF
UK6gxVwsfnWaVCDzlvVn6tQtUL9gEvX2szP4CJLuqE73DQeDARyE6/51Q1uwtjJ+Oq3c1MU1A3BU
XQ3GTsMDOBhIsjUxFOKHNQZpZMp3wa/wTBNmexVx7a5YkI/4QSD4tZdjSI2ttCiY4P3GwpbBteWv
24pnpwWn4i9WSwfeVapRDxcy2cfeR3kMQWbQh4SXoDzJ9jIHaoBdEpPU5uGU33aT1xKEI22VoCWq
K7dRd58Q83B0Zqi7WMDnzL25ya/QTWJONjLB8f7d9WrX+JHlRQttD3JpAyUpgedWYzbGpLUITjU/
Q7KA3gHblg/KtIKz3+EocC3EzGU8dy6ghvKMVIy8wt1v6oMqgVBdo4x9dd7BxykHsLgzivzY7sxR
ZC/YWw6nnO8FxBL1XTohh/WehNT3axKXT8JyjSv3XHcbyM32Aclwl+3uQUWHHtfQWsDaGRZzFi1Y
wFlLkaDmcChqDs0uRKdjEm36wp6yzMVnwRlU2hrvH8r7ZoRhWCkN24f+9JnzFuJ0ZtffGC/Cs0Sb
aavUnBplxpLAEAkOkt14MAjCNHUjVSUCd5Q2eqE2Z8muPLYVjSJf8EqQkrlADoPuPHwCCmHxbfUh
ntRymTsi7NQsN/UQ8412NcGzNPC3g5sxgEqJi29WiSQqDISptOLi1M9oFOuxUyVlbfiXETq+UgKt
V9oCa+qbCYit6WaXLqXxShXBFNJV1XdZcBa5LTDXHboJ+zYy0HqvOUkwrTjyHipgEaxm1cu+Dt6t
CiGgchCBrr3SSGS8NLTze6CsPUdLbmLEvReughXr4e0YF2fS/ZE+2TDq6Dd3NL0JVxHGotuF9C5/
v6paslTwBzAE6pdmlt0OiDb7Nr+CnR6NuprHUnPwWu/otLSX5yJtbVQXDtfccdd/KwX2M+Oy3vZz
VIJK6Fi9MyPpdcFGantLjSAIxskMcQPJbmB+Yi7Zwq8+IBQAyzdZ4A501AyDJPplv1uQb+25y0oC
W7O5QnxTUMlXZPGLn3LCs1dzzgdzYnrz0N+Rzc4hy476nIVhqbIZ/CLk/tENWM/2h0H++vxkVDpF
RNLxL1MujyiPEylePdM7z9jJc5GsVbTziXSOjK9or8st1A1NoFUHhxI2PV+fXjy11scGCh1OTpI0
5aoKZ3WOoIuWUpTu7nHaiCx06KI2iDApBXI3o3qHfbjqSyzMhjeVFTyeYtUcoYl4RTzE4X5EroXN
eAZn73eAlxCbRsQSx1X+8zCzF4oAp2ubcaFqnOdTsz/9ueatqy9iO8K06EFR5aSCtJ2u+NgBdmH8
euBt2bl+ENy60mNgPbEiN6cW779dw4lUAmnm8iMgfUCiB4/28zT/1485QcunrXma36a+0ZudmwkN
bbKkMs4OAZLoUSKHOjTdVAi2FhNHxGT8WwbJFVCCoYkmbHoLqzUJhBSVKubugRy4FzxfBfTqMvWo
SJcJVywm9UwxqgyOGlNdnhVNUyg88mTqerRese7OVda+u9/Z4qdKUutl+rCgZZ3B6p0ooiQa3b0P
KKX+zRHB84n9jXUUjjSW2wwR8Hg9TglI1XVi90E7sxxl+LfPhTi8E+7xybvgxMgMfxpByvUdzUFT
m0OsO+yJlZ5tKwwWgvjlwW/XbbdusJtlFmooR/Rqf8Z7wBUwcywEZsGTj5zhruG7bM4n5DRTFAXL
4HnlzK4EAA3EmBILn98quKfGdKvlZdocg3EcQcTOyO1c3k9vIuQ6U7uvnaiMBMNIA4dR9r7SW/5z
JKu83+dw5jcWll7eA/+BFQOAHgJXVfxWBMyYmdxOuitLGd/k5WSDuvv1ArYJUZOsv8YiolLubQ2V
m630uUI4WBbaHR6SOC//j0Uvf/NZPaYWFeOPKrFaRTjQsKvgq9fb/aKwuNnX8/HMh6FE8JtuGLZo
NJr1BC5BrQ/dBJuhlKvzIWflUZIB1N0536nycCEeGIUMJ5UGdIApmy7UO+dzO15+KeS1EZetS7pB
mVqoioo2wOCp8SL+pYq2TpddmMnQxr+I6fNs3xgzvLJL0h2gG4AOTAI1YhPX1/GqR7i8GyHkBNLm
HXe6VnIIG8fjvvGuIz/zUfRTjXHr00fnvBYhZ9v+8YfMaC66Y1hM9/lD02lpS7AKonlk9r9UFEZ1
blu/XVZwh2/wzq6uCuBHobck0Cl/OLg3unHHcSGco0S8qARJyTyr2yOr5aD+jJjuT3OrOYoewWQP
rkAAXnVqb2vAZS8wccH85MW1MZvfyzHcBlDEty71wAE0yt2FHvVP4Vs9R+bR08hQUGZKyRwN/LiV
0Fcr2XEOurcNpK1V0unRa7DdthGFLMTp8v8bP37vq7MljsJiACEjBeFSQ/WlHAXV5zaCYL9u1jPC
SdZkTeYlBv9Nu81CoLRJ/Vfsu8LZ7CdkCY8Tr4zRC5VxQZmy3XkTaIXKgwqAJjEy6QrWorimfxMM
5Z/T0yjEIxojQfwklpjl3Ach9rbnQ/q+M7Xa70dpF/hzyyUmeN7HsS9plbuxEBnP7MRaT2SjtaMc
R/XbT43JTSTGCw1BzZncLhNbfXL1duf7lMAPo6d6gincOJZiFJWwIMYaiE7iccShft3YAe85Sbgn
PIw1Me4T1vRs2cDsQkS82XvSKXPgFYiIgjYZeu0Tq54WebXXs7kd0GMOIbbfRr7kB69rm90g+F4U
woHRfeghSEb2XZAzkODzqR4Y9+Ag1VThYMLntxqknOoA+E8Wvx8uPgSOOfwq74PGYLLarkQdXYik
wnriHvi/hkH3nRqqI0ebJ6yoE/4k4tYTOtsxP8ltNZjuT38ib5gGJZEHh6PdnNB9DAb3+NJgZWW2
gEcHJlamif5o/ZKUXXvygJzVIokp6hQTjb8/Dhct/C94edhPf8YilGLSf3JYp39apXI+vpUcPs/X
3R/5fsQXFTy6hPX2tziUgMiMwTmt7cygGkcRLxxvDECQavtc571OyTKijwWGrW0EUVRKi0zieb5d
d70Ca50xSIEWk20yR89uOlPB4Q2GlZnUv4aNCP8NuLykKlo+sILYLYR6EO9pzw10+OcsJWaK8fMN
mIKXkTflJzzg4/VyBQvVKzRcWhfhIw7UkRXJ6JxVJai4DVYkplsvmhYzCk+Av+HDwIG8mlsds8wF
ytPbFMGhmK+qJITcnwPWfErbnTCmaw1udxu/1UBh8GS68V0c6G+ntDosbJSpMGuPhqD5E81IuWDl
a7aA6+aCLWXEbO/a5yAatCv9IzaHu3HugRZR84R3wFhR9U0nSQhlBPOqQNgNOno8/7bLx1uqi7v0
XFFAqdF1cOqcj7IbvIqlrjwxowBirhOfGHR9DuA4yaomHDaboJkfS6lCN8PsZKt6iMpA/wlB4Myc
2lUFyRJqAaP2RDwIuMliZ1uG6rAgFmybk+9lwqNDAzkXhn29SsbUOzzxurAXbAg775lINtohSMEr
9ffoWaXzHE4c9ljHa4TG8pK1HqEOs5MeVuSHLTYLyPxG+ZgjajoUUVno4Bqay+bdXA6LDif661Ow
c3tld65WOs+9r1RwV32ft36TO+XykmfoNMyJEAQcuWZthl6gS83kZ0KGCBuc0KgOAXtf1WMpx5M+
UqiCuYJUEzAw2Z1k5nNJ81HZLSDkNCg5LkD0qvxEmrthBZhrWZzYRAj83XGEKk4RPbZxx2qwHdW6
mfW0dBDcPhWey6XGZnPBFMcwZmyMbQuPSRUKRKX344C4odp7xX8ixVenGKHXWexBG5qMqRaloZwj
riEq/041XPA4KAFXULy3foZl7HFTYSBwgvap529Fsxpi6vng9KsJFjn5hq9SstuoVQeZ//sxKSNF
/mGC0JW82Q8KYRuhKJObQOEkpNGMIuqzIy7KN/g35F8VJ88W2i5w4DPSIM8OZXd88QG5Uts3x6FI
0DPMfmP6wl4KaocejYb2tDPtBNH9+LJ++m3UOyTMgfpHM+9fTSAOwMvU1CuPw0Q8grDlJk5qLCX3
P3cITa+Bm5lmpYePULgxgZUH/rZg8taS7vrzwlGsxZ2UrRmH7stZjzL0AcSswLCRyccyHVrMdWZA
+SprfqzBhmklbMjLqGi6AoYZdTSzcAcNOccyfmcLGhUTPPFdkdyalP9frWkNDuKoADrhG+NE7stP
K8nnwgL4ZP0L+9yXq3GLAmE08R9Godtg4kkvFNdKs8nPGm9Vh0mVpuPFOtuASD8FZcW93mB0c5Oq
OtFdCZ2S1wdKQGdqceyO4OhGrWBO0m6dtSVwQ4kZSQULWqPCmRENhezxLQW3eCOU0JVy4tzAzjQT
NBaTaYNauOdULMMzQK3UiQ/W7iUAPRVSq65z8mn5IAd/9VPL50EcPod21PHKxOiEyK2dwaFL9eA1
BZvc2A24hIUodUkTSftGE0KQ4xDZ3U1fQJZGxej7V62N9SvuKGA1G8Ow7/A5s9hcj14mY3Q0uTqE
vD1XvahlVYmyhhTKBZ77h2WFXCBGSGkfaI9vDlH7/9PJDd2sSdzf/ZLo5R65NYAJMFZLy+IB/osB
hZC0sKvaVcKmdt1+L8sQjTtqAV5iO9CWos8SGueZG5/1HxzvkgRqE5ugB5HrtIE1bqlZQOzov71+
bPxtRmvwwZcl/Q4wuiy1lAwCPbgoq0RScqaQd6Ec8qJQoOxrccm8CIkdoYhA8OIbsSqVPcOWAU4k
B00wMXcUgfuKFzaZkUEkeo7ZTiDfGtf6e9qZNLHyzdHJXbCw7EaQU2gMyorg34TEj0eYECpSF5p4
eGiLkNqJMt0rEYeK8unIPKX+b/wzxnWsBH3Dl0kn7N3bvKVYCJkbGPhMQeplPs4hfb7mXY4+U3li
lje8P+JMahfVzS4JSawlkDT91OhdKXtccPs81IKzhXf1Oqdew5Wxw2oRMkAhb+IGk+16YBU/zW8/
UQN6e51SNlxEj7xWKZvBZwfSfZl/DccRI5gyJOYKtAdnB63FeDyuIaC4uuJmh2vpzre6ybMTQb1U
yh1ExwAHphGijrN+TqEKmJyoFiJKyfvj2W6e1ejO9+SARuaGIJjZGnEDn7yCUZRNbxPYCKsPoKJl
5J+fx4DfBwvhn8aUGs9naYx/F4l6vW+qgocv3N0v//prtEL5joU56xEfROhcbbucSEgeh1PSv9q2
amjrSxTz8o7xNGc62bK7BLwjLHHfFfQOao05a/YBE5pej67chlU+7nzlUQH9Ps2QqmsAtkfEp/n/
VJpauRU2eonibv9ewYhCKaUv1wLOsfF1O+PAi7Hk+LVKPX8OlwSiQ3nEPOPPcMs99mYE3+YBXnp7
EAczHixmL0owpI0lfvrN7/PDddoyR2N3w84GSVPfYxzK1Zb6HvY9qRZEED4bQFLWXfzpfEbVf6r+
qq3Z60GDdEReKtiSy1SRC+LZ3RCtuVyZkL6QMvqtvL+wL/xinpp99DF2hw4NBH+hzzobE7Cpu4ZO
Xtr4QGT8LD38nVoxXNt/Tx0C5fAuz6KC4wEOYzK1sEtuCbL9fEm4oedxIlVHfBh5cj9d2mASmGHh
/56RoGK2HDPGojkUalqp72nRD7aMc6n8UIMSCp5MQbUbU7ms8qVdUC1D6zmDkCqiViFhovLeMXxd
67NDyN0r1GITyooJIEgnN52DughyF8WP2JDSGVFoIZatTw5L5rl8384s5rOncORUSJ2JcJ4Z9Pmr
awOKUVZQG7D0SoJGz8cJDZXxJir9noMKcjxnLonkArG6iW8PbyJPUYrVX6RGGEyb4U3cuhjKeTXG
redf60NvdyWaLWBrIm3alodNncjY5adFq10XTeads3z9fxEV4RmTGFvI1S0sDCYQTH9QDHAfNd/t
/mj95HucBLk0jzBLIZqNBvez22dNfrYu4fnmZB4vF0h+ZSjL7v4csQ056Tmyalk9aC/21yDRof2m
TysJIF7SnuCJ0hg+x9bihX2Oa+9bGdF8ipafBA4qLuQ3uijEK0nlIG1qYGOsOCy/nKX2OmZ5+GZK
ZHBvcWv4FfxswYcxrwitUjB0YxN7v+J6fewoPgeiH8HiLxVbgrXMxZxDTwpZEIDxO+McYPRIfCma
Yo8jXvgFtaguWW/i3KqJrZCan4MX+b3J+8xa50yIVelmYTit8+4Y58MUNuXRhgHMPPHTwCcu5LOF
GBM8hAaT5SE6lxJHDz2BuO6CS4nFGMczaaA8kslopcVOhyUKNvfYaOFyrTo02WhQpOUn78gucdQ4
iL3gCm4ytzjqOr+arZwJzyXqtURp1rdktylTuZumXrie1Cz0Yu3ecaMG6XL560FqFUvNmONIDwXb
dV8P/eSLpELuCfmWwfc7kijDPqpqnGkOatvcB1MNL+JaD3FHPalGZyp0zHlAY4JGykTcrFnnaz+2
S40IbDP7M7sqmKx5IiAB05PRPThnZo/phUVulSxsqU4kmmY7z3+5+L7SpP41KLlnjHIhilUKiHIs
ldygIFLCMde32dXtBnrd2PRMqG2sumuhi0Xb8gaCRtirVAFXAnkLcQHc7DXL2Ip601At3Hfk6PfG
BAdJWaszG7v0E/F7h1YeFmOot7+8YgGm7uSiLCUTSBM2UFombwP4deu94/rlq9Ywh8mkkNZQFNrc
b72VExOV/flK/vvf4HmiWXw7cNIKNjLF7NcUf+ykNuIZOIBNa9qh2u2foV1vWMR0w5ZWSMQjQguc
HESEWeZm54qCL8RnAhc1nhd5mWgmaxZCQOAVaSkWcE+tNoh+OOGSJiedEtsR+7qAR+vwFInWmHy4
1keqToJjUpuhwRLyg/FB64LC/FGRO9NDsKUKENqSSRMh6igTzxVz7G9niR8sHUH/IBywQhxKg3p2
/5AI1RVhp8AI2L6BNLb9x+hoBC8AQAAZ5TXwaVu2XD8lCJFp3enqLRvz4oj05sDtXVE40covPmRu
f5E6pVUOv2WavlkdGy+ZghQuA/l8HxAQTdfiAFIfmk7Lx01+bymKIe/M8HAuAvQVQdeh3/3ptj9e
hPSn0GNpHQx4TTWYYqxAfJtNhkRktqFfRnDshYrA1XUblgKG7BP+wmxEm+O6tkcFUZSUOwEhWyqE
YvCEG8kHPQjQTxWgVHNmPZMppWAAhNTcfjgbs51QWOAzXARSftevqY5Cg23lhPz7rqVFUR9DaQwJ
KYA6Bog6ioBwoNhipBe8+P2repL/sl5UhBZuFfg5bzeZs9RKCOExgURUr8BW6ye+6igKFArSKrT4
qCJjtVYy8okTnU+AbIDIc0GRpHBbIV0u9WEJQy3tLpJcfja20ME5uBSLdQkGPbrhkcS+5j/MXokd
iViJYmHClcvfA5BykqiADRCJIJQIMwoO8yccPY7yE8FsC8/+WzLAd86WYrj5pyvR8dGmQSztTy2E
oDSR+z5reem04pwjKmLevpUyOOf4KSOldHxIrzdDu7vHvW9pehUS4w3sYiRF8OOorXY2Dkf7IfeI
MUQ98t25o41znRb4T3hTe0Kx91VQGpxNOqbvnm5OLAjpYZJilF2AI5VYvt1wpt3w5n192X8dEIye
xq9h8xG8+q8ozc2A4Kgp0bTnlwMo+o0NAPZA6LCm7lbMf02KMDu/W+L8/f/dIwBwjW1HiKNxI5ly
HQkeUMWY41OYcldEJITskzWkH4Gcog1QvHx9nXdJmUegcBWtEBfx9UBRm8963WqGv88w18jTCaj9
tl4AkNtiSuN/06EUDNWsD9K+Pm3ybPS2/ASDCU6KGc/Vz8XovRtcki/yJxLc8PY0qiyjd7H7pBCc
ymosN6B9cMY85KCwUHFDc5zsUPPTwBtIQoBcYJOYimJbW1/+yR+jQtJBBBElKKWHzTrBXFAPJWWi
4eVlG//3j9oT1h8SVB872+Yrm0YnxQ7Z9i1yVBhkEqJ/1H79C3QeRNRFD7U9DtXZo7zUm7T1KC6L
tscvRTSm/GjihKzwabm1PQ8VZARcXRHNon2CZeZqkDwzotirRXV9/xZKFRuzPXy5iCjGv3iz8Ble
b2MwNQApX/Wohi/IA+svxs7/oYRI6mJe9iLjvh/bxIAwtY6FPBwzRJx/nUaxMCfqhfSE+NRbKns9
jp4N1wDsk+WpBtpH867ILm/gUIYS2MH9lAYik/OSAYNT0bp0DOs7D2D6AsCZaNS7K4AO/vO6Xey9
7c0NdXZaAgO8lejvp+w58Uj62d6eVe0bQm/DjHbEHtILr/xrQ/wDJxbOJiFtO7gxi/aWOXnqb0K6
8KiTL5R5ZcpVItlWJ8KSwUvc4EDsr4py9zjwYq5S3X0ZHQ2vK6W8aLG7uTk5e2ddD9inPDjzo7Ob
EfFbgbf3brV63rj7qMn4baQFVfXsL2OaTiYkGwZXwu3IgSfBeIvRTZPraweND7qbxdgCac+UEKFE
b6s7kOJB1B67N5RkMgN5W5Z34PJ2QVCsZ9f/9yT23EzvUHI5FWQCnwPsK16y8RmHve0+upE1YPsU
bjhwa/gwNNEigw45VOyr20CAP4iyCK1bIUnHazb+AFgbY8RzDmf0phKZ7R4oEpSozQ4taWEB+iVg
T7xE41+6gnqhW9f+bpTSsLFTnQM/cBrEV8nbwcxMB6wYvvSnqhxdZmpkfisYZiCZT10zCyyBecFz
aWbWUaDYWDdGJcMDqNiev88/6geu/g+iIZRhDz+fY1VCUmNQA4flrEqFjrPRhN2Xhvi5qkNgLkjq
0L7I12/DEy2UMlItptNDkXfnf9Qvb/ZRYCZwvQkRxMWh9SCQV8xOLPl57C065SSykf7slYNtnyqx
uoyMJuZTDgi2QtyRj69A0IusCwrZCAWd/rPHA+UQ7ACSjQHf67robMOvp5v11ccJPaZEuBfM/4E/
FDXlsstnijKSilyauZPOaIJywp4hKcB4hgV/FkkYd2/6s9EBVoy2bnXTuvBie2641/k5g8pkj3/W
HmRak6IZssKB31/NaCEXkFv7FeblkoVOnfXl5/0+rUd3eEtiCxdJ0EnD5/F3kRlh9lDrhIRTI0Bh
gvmTPRlKwiCoXmxxFuoSaPP/xMiSQpkucg+R4/KoUsemMQ9QYuOKMpBtVzHbKXs7/9Ij4YGOkpQ8
JWjaV9AfXN5qUTaDNDKrAnilzSZe6BaISDb1/j8F46ALfQ83umgBeUM6rW199wPOW3YFIbqlOtuL
8FkM31hgO46ARkLC3wb/R9NeLLELl6vh1b4MjUrXh+vrDYa/FWVNyrJqGmgLYEAEXaBpjGFls6zW
UHpnBwoaQUhUaJi7X8RBXH6L5bp3/zAOOYPVfIPm+EUSu50FUO4yiLTHmYcdltWntfzridBSEU1+
dUBsyBkaYUU7kpstmPLpgDHOgEsAvnOSWNsgdLJnKC5S8nOA4xmazPG+D+CgnNRAJJt8BBRo8+h3
YZWNQRw/Tmm59siai2DP0GSaHazTv6rZOXu97dRZX8RAuvyuXmm5pEdLCG9iUBJXk5ZlLdvbVynp
a4KtEReEyBw0gVz0TvcQP1qgF28zKxlxApsWSkdYR9r3CA9R+7g8DFSl1ngSSPiG7SDvb7UpBe/F
unYoo+D3mrdDdDNE7l+3jK9O3wxlH282JgKVfx+2ZE/kASVo0+E8nT/WR1/GiUY2ZwX4wgImttv5
F4/WCNJzJVCwiTLZtoD3+3A4RItoPCm/vN8T4HQ0iizG6TJB1inn7rXGw+0XuRsK92Xdoo4RQ8pn
vcCL1AS54KFdTjyAxyuUKiQGp45RWeZrmgaVC8xAbS9FsWGTKCCh+TdG8YYFnNkc6J0UTQPSmPGa
tIwjCX0y+8R56V8d1/RZ7jxvp/YSAJpR1EjcicDF29LY+NM4ksTJAZC4VKG1al+08i99fXQRTUDW
ZET/WB3YFcDDuH7agobRvqbkxjEVLxSZqM46JE2DuVAcAFkxDSMqwyuDt8yHFtAUBnl6BC1qqf09
PaexA2Xk1VnHcljBpZY3g5JBzXiqrYHWqaXEEaDwH4BABtqIhuxCPWqe8Z54kz+ALx46Xz5LnggK
YHsWXOk81iwqwH3IWV7JiYeZ3wltQMz3hjCrDr0o6f+EgAl3RhLiX7BAqPa8DRKt099ZQBbCs5K6
1pRDOOIBw+ZwiHYzYy+pAl/6PLGKcR0lhA+AwKYoEj39tqm2vHoKEAo0SheLB1nmZbPSDkyiAvUo
KmeQcp5kcoV0aVO81n33GXXYptc+brYfG6ZVeSR8ay2D4/23zCZtzZ6jZQd2qm7u3AnprL498Q1x
q95pbPnokIb/JcI/AcJKDOiptxchmFUpRyJ9Iq5rCwWkmKu+7QPOuFd1NNmRLVd7/ZU2IMMxsy3l
8dI0SMx0+RFx/3n8JaiyvXfX06246xYGXj/x9ElwG+M638fb/OpvEArqNeLi4w+6IeZtSdftoV4H
01+OyBNQtOddOyLciAHJoevkTpZF9NoRJafobCh19aEF5xsQHEOIxFq0QmTH7k8bIULYzc/3JiGf
BwSGE+9wF+MU3GWnoqds5v6P9P5Od2J7wJ629YvNJcOzHrP3T6z28NwJ+fE4XeSyAs/6PN4Sf6sB
7w3iZAadmdIFBroQKhIezak8v81TEXmWRGp7qbXyw2zlUod6H78EP9C2KzyxIie1p+3GvXoDhzTX
bGzfSlAOfS1cUiCFrt5LJ2DepBvO/1vVR0tPGnRNacktI6Q9aDVYTTZoMfMXEAc/enBmEMbeaTAv
uaRoS01fE5IZw3ZxJhGgvnblJxXtNOfhXpwxCttKm4X9vmCgZB7EqPwbbYTCqRHnC8uXHP11CaQx
NuZTEO1cjfPe+TtbEcVZWFrSb4epoxgIaNV/Uzpp+YFLLWc/R7RhXH00uzNqQ6e4SfYgA5PU8QWf
9Nd8jtjGGdqIib/LjyCpEFi0mR46+e80VFgyZY0CLnhDFtx17CWUHSH5h1jud7QgIDBe6E46Dxrl
hn9j1aPoOJ1tCJnCW9+aeynTm9nIDyufwAgspr8JovarC+zHUuLgNzojQ8/VKj/2zOwCuIY6OKUw
Xn61voynqq85g7To6RR1dviiHviHEUjh3GutnTCyVzQYGjOU8GptRP1BpSQUiXRWD/m8aRqoH0U6
JcU9//lMilwQIC4JJVqbUS/7DDxu0prildcV8unu6SO7CEK57/Eqyng94sYbzQjjT1mhMUn2HanM
zZOT3bZ9a1xJtIrDQD0z1e0hD3gwcIkMKfINW5TuANoyc0Dgc08QCx0WfbZQxUmI00qILIEaCEBP
tybj+ERvg64vbVSm2HHlij4YBhyit8BYc1nfLStFMtjD6Bhrs25yfng0wmI59l6RC5RnsihHrN5l
4jES6sE6bHzH4wUBxdsPqeivYNkP3KIHFvCm1+vSPdqUFPPkB7FXpJ4MlFWqIRQuoYEsv3Nniq9j
lZ5jcrxtlmz4awGbOPLLs/dz5xX5ZyQG3mVsViUP1K/a7moUjlgIjyHvnJ8afCqpLOw+Ur3xgk/i
UzKSYHelMO5xBa6b6PeuDUzQDib30Jzzzv1TJ7TObFEel94gJwRdaUM4JMrnbf3vUhUUbxFvsQAr
95PdtnnOdexCmCZx0V5kHCLmMMzoKBtqbrHnq+hegrZXW8ah8HfA6W8yM8x93v/O7ZC+tOonbhYs
3QkbM9vjGGCpmUlLyVqsOz5rNL9IZgJBBEVTf9WcA4tuOscSeELFLCYgaY/WqzXqc94iAqlBy25S
kWbrpYfHnJ2W7Iuekx4YEoQoM8OIPrWIZrPXfXacW6IOAv8uWwUIubtfWBE76CC2AZM39moupyG9
e/hB+FLoMANRo10LvzddknZTW3flxz/AHReAfuGsfnzWGXRl8O4Owv0etexd8t+1X4oKijJvqAlG
Ow5oANtL18kBr7IDWrGgWRVl/bsxXI+P9LAEf7w3NPRypDoI6nK9lcZ06Dd53HDdWZxq8P9Oy2Tf
KDEUyaozdd82Ap5KKSc8cQUxhA+lp3QZgGstoXYtuNkQiY9FY/bl1fsd2x2ETw4FW42gHcxkJpye
Ip2moDmsRkrsnEZ79dLsuzgqiD1oWCqn/PFI9LQl1YNfVbxqJg/Vc9HqlLeC9CfeuTHtSDkv8hH/
QKnpk+P1L08P83yEMgKimeOVRp28GV9Mz1gTP/g/6cEuYcqxNCYarfk8X/AFQkAo/fLbIxC8KIDK
jpq3ZXxaURsKEeRxxrcHLNISVy161lMzcWvSKWMAh/CswDSHcfUiEOL/4Im/MIna9aQ6edwaFeiH
hoSv6P3bkQg7oFq0xCN8rr4wEe861edkMoQPWLML6dqxl2gLpFip5hMP3si5SqIekAsS0K1hfJan
/AZInEOtxBBw4gNc9Ck6aN3krg+AsTKO+LE8EEzCAG9051c98IMOmr4DoWN5ecRh6H5b9VRfsE8C
SniRwcSJ/VB6SH79E5dGLL+5CEgOSaN4Rc0sn+FenkADI7kWQp7EOZ8S/3mckJF+Q1TrUMxnDp25
riPeLzLyEaCFdiVJoNoBykZy3mSOF3HzF1koywfspdIDA/Gz5TiFPtZme8GleHhenuFVUC2V4JWI
0YFDCc8d8+3JzwHZ/4356UZyFWpdQXn6YWSSuap8yaXCh4dvHpOvX6rVsbblT0VvJTofJXUPL8TT
v7jUPc7HD4yk/gG5AdkBmw0++BWS7Z+OFcwS13rxjYHKo9jj8XnI5RlJ63kFh3dFZpBNorJfSZ/N
Ydw4v+zvGg6AUCh3X6mtY+rLB0LfkSU6G934GKphdPskR27JqCDKf77Bk8H+1Q2h/JaCzxMITSQE
1uZc5rYRd/mpLIrcG/mVF4uJWOjFbMNrBRR21RAtzMh1j6bXuAL+VNysxTMKAtvXt1Ga9osFTzrB
ZAGV1542taREVnWQK/ZWWVm8FjOUoOIBPL+Uhpfqr1UZcKwaBrm6bUcXZSOCCqFBGmVAlgDbdMu0
RX+1qPAmXBtWkaZmFPweT6xfwIkrhIbzHoVUJr2Q+rmZSM9CiAnI2//mc+ijOzqfJs/zv41O/+7w
l1KkmWfDnXWpyKJYvxAghyZffHeFF0i/cOV7kvtj72+RbhSAQbVAegRRJosv05F2UqgKc1buWX4o
YQARfuTUZ+HBP/McMWhLWR+hillwRstF5WQD0nwqCY+c2spnW04ULPdZPVPqFMD3cuBxszv07g0A
B3P4urMrh9ahQGM1JmdLxYPWY24kp27viLmbdF8WA+fPCQeqNQ11Vn98GtVv3luV94sA3rTuNlYu
MgbiukjKLBU/xFVBUt4G+6nL5QI08gJwbbSfMoHZy4P7f5vXr4VIDU7UJpg3GluZkj9FgHyVHlgt
6Y7dAL9f6WBYB0UZGYBjQBBQpFzgix5pSo/7mQ4q4RP7yRbvaXKvoQN9oQg4mSl/+EJIq6t9f7aV
cVefHiW7sEJ05vGgHLNlkG7JSTMsPSWL6z7NYubCa0Zsa2WlDk3I7SsV5tHoht+ILLvxc8+U6ogS
KLssy/N/yANwpZHe+fIx0dPe9COcpbwqs7uzslzxOzsOit/zhL3Fz1x3wGVzGClO84ks0LN/XrVZ
SbGteGvMOFXbnSWHsn/Pw/DJOTQJAVvSCf/7BGCGhGx6WL2WAj5mhGUHrKbIlBSsOjL6LxNT1slc
J7/rx9/seX+Qak98Dv7WcyJ37m8yNR7Qp4J8wjLYD/5pKKwnRYwL7/GBHQEWj3osOIGQ+2dR5v+0
eh6FnZeIAqnEsyV0L+tPZR10fO/KpdTUi90cg4T8OdbSo9iDzQV7/Fj5ebH70ckEHCA52NtwLBSn
6QnacZrdqXuiuP9qbdyMmiqCJhCXd41114HTYdxqsJeGsShIf8GTVd6DNNP8iqvAqs8USXg1X26u
VJT1oy1WrNEYETV8FQWPNzhm7Mt4sgOlb/39gLAR70VOHzCkb545da+VoB/02m8G3bnLIOKqVylK
o8w1P9p6uuiZqXlbvK+ieFsCWY63ERxXo2rSyseEWrXF7MHKv5HQMTBNVz1wuyFr5YpdsXlhG9qq
/hrDQFVrx1qBL2YlO8d5RWYh6DxqCJkJd6YEsmsYNJjOyjc5LIs8TDB6WDv7IS/VzKlOSBB5xe3j
/9oekVtFtmUSPOt2aI/mGg7zBIXmFg9MYhwrR2T2eou3SIrH3ojl4iSURb8ugOXoD9RzD2DHnDoC
mIFOOfno5I+5fNGl4ulAFZ7f3+UBpQoa/BVgtsG0lQjj88G4kK9uDVcFQ9BH7JCNJv4M0fNNdE5Z
NValBF2i93uNFcO8Vsq60Os16sN0nDzh8GB3mg4RzHyNN+BglIW5n3XiizXavrIdMu1kA6/WLzE0
tyZV7RwMQ3oFjk/8kv3UNeMduABiNnzpblftmqXzDc2qZUjc/69ZydbjmER2lt7YTMbaqLAdybMc
gQZ1k753p1Wi+ivzJf33TeKA5TpMXptiJUuYahypRxghc5esklvGl2MV9J7YEbFRJUccJcaUuasW
x4YJ5yDb5KZ6Tv6ZWGgraLSIpGfRYnbhmkksit/6+xXxUoblSHaRICS9/G/7+0PVqMS1UMVrX46r
6gNQpUa8xhmli075HSmOVmOC5nKhyAHt1o9jve6hQS+/6lIOUj9JMoPSm6rxIU1OVgbyuDrikijZ
GDckkiXqmyiIksTw1fcbisxvorr3WGyV37yXUySwrzk1PjRj8w8bPCC33O/SvV1PZAANotGVN5Fr
Ptq6EFA0rQFgHv0R57a/DfkecKZdgSYlz0q/UYbnd0aUJdFIT7xI1Sn6ZN4cdIysQ5uuB8BJRo2/
z6mBRq29IMJe0GqG/M0e/470NIVkfKvoV3zVqkEuAlpC50rGrEq8NRRJ8DbynqA7SM/NNvHyP0ve
fgK/HgRUKPCSKfwRZAt9Dbl/SRuric+WMWfEIZOthoMH1J7dTimUtNzFFcX20tPZnk8JMZimYugw
8D9e+ZhsYdvAtT73NYl4f/rRJzmZezyyLjzy9nhwIjphfLxrhqiVIdjsFwudHP2ExQXo1RmhT2y1
r00PCnn0o3WEscjePOMo9908xou/5IayfKkfN7gP0yFlriiVe8o285GYJta3tl5hcPH/luqA7JMU
dfXC04PQMz251NOULZR7EmsVnxgSVq/pM7cnEFelPKep/Xj3tOqKuwhL2NPA63OM8yqGutOQt7LW
QkUDA49SRCUYKcLy7Rm3t39T2I8oShU+u/Gk2cTqbVmOCxwvMAodGfV4xAh7m2oYzhSX6IKpjUgB
H/fBiq4Pcbkj4N4Ra66EeAupW5ZHiAkQk8Mm5Ny3GoknlA6GXLOZnNVieW5/lhMJlh8HNMCa6Vqj
zxVa6EDa7YkQmgM1M4BSx7F4XU2ZMwWFAmR3AhevYV2hdTNf1ccbUzA6ls4dwPOpyyguqni0ohm+
6f4HpZigjho3XZUXcyLKb8Aq2kKftymVfKQz2vdYMAiMlFTGPHrWyNQTm2NnveqA3JVoG3ljA1uD
rl7TcFyFmOMfoKWrjgthGMmHNDYIy3CtSOn0SkdDeCB+IawE6ffnb8m7V0syPoMLme1O7dq3jciS
nhgWG1CxOtu9rKGIbr5Y5pp7lDm5YEKyi21gO5Mv9oU/lgiPqzh1x94MbLjrEP2G/v9gF+/8RJWx
D75IU9OELxfmkU2eAxRtrASwrXQd5S4YCTpI5HC/9rr+RsER7djg43X4rAIqBKsUu8+D+l3cyqiK
rkiZ/hsUaE7g960kQnxipo1EeT0TXF7IVDd50AZRtm4SLHaId1gB7x8NwDnj1f9tUMQDSOmMOmj1
p0jxeac32q29HrYoyMuLCy45JriEXyyXW3xDS2sZaUyliy/vkVynwv6cpVczRx5mRvCUL3R2CGr5
e1iz9M+rTV77gkxDaES4KER3FEpxKaYgYr2m7iWxGDECTKFk9QlZGw07FxcXAaZ71uDahKT2BWB9
6hKtl2taqQx8ZIMQpeuiLAosuUFYcogCqX+sU71n8x4r7NP5L9FmIganwQmq/1OL/wTfFsS9ZN3W
7759jWNQ5bVqd6sBdFX3+VucmW36C2+LWDrNeGjpk/6u1XrXHXyH3I6L5nLHn3aLv9VjbTTIutBs
gnyHTSUdDevRkGh5PAXmfx8ac1Tor0qGbl2SVG3jxQqcvk2OY/IW4qKMK+3yRFRwm6ReNh3KtnzN
YP/3K1L90wrtP0fb7ohZh3vVNUngSnyT1kUtY5aiaW4XibHW7WKICxz+78MYJjzalDuB9wsC3FD/
pMQdoAdp/q8oqNOemjfsNpCizv5StaIlzeeAAhTe4n9i+yclcZCbBPEt2IujQ8r0o9jhIFjPhnSv
cpDsXaP045BN3wP2Ds7RuSWoZZFMub0+Vy+oq/sW1bz66mvDAZ3hylsqkmoWLu1Rm7yVLEYzStzh
CP7XRX7A0x5QkSAZfEfPSy85KPuFMKMXdF2wsf2zB5rkyrSbhPWgKL7yOaP3+BKOXtVjtsaXXq2P
9gn/xF8RvtLbCn7mDD9/LHXSrSVWg34QZO8rj3iVObNL2BI08JNNYLWw6tLoJUyi8MtXB7Vjlq9l
K3QaX78wajKrTMMETmwtO8VPMX3SXjULU04KLS/WlyQ4BZoiwAxjdHNLm0qt1osQ74HZOst69Ne3
RcIXRuWfGTHnd6jxusO+p7ZizhFOIfN7itdWak0m4WhAerwhMHeSv3TL3TwODhhLIF7L8RUNp/6N
VQTXclX913Q3BVK982pq8uR86eVq6w7N7AOXibXqSOfEwkv/leRZ2KB4aM10WpYpL0NXlWJq6Fj9
9j+RZKdU/MJsG2PvIEfY5WkJtdtu2wzpIJrGu1uJcdj75cdwXDJUpHUuh77VYdhl9tZfIxc/jlUw
TJ+1s+ewueBO66X6SxfJPXYjDQUVqDAmK8LdTDrgcg983+rUNOoLVwAyThj+90sGQ5josvLy21zh
gVNNnmUIfV0iKGMY+6vg0sSMcolaAQycfFzooAeHZpl1aEiH86HyfKbNBsflJ8TU2JX0yubxIFdc
nvN5msXnlIbaqQgMJpd7SK9EkG6hUKIEG8OBH0RMwfOI9POENN5DkOj3uGxhaoE5e/E0KXqsBa8I
9eGMOEAobGUzc8E0VFiGjk+HQC8T99IfqL/LteqNtlidybKddDwLjp0T7N1tfP8ru4ngiC8Edrtn
V33fddsV+LW2mjan3+MObkk66S9vZKuFUK6aNfCa8pz+5ynHT5ir57NHhx3ZiaWz1jcJis+eYsVn
m4MfvzZ0NbY5frKnF1L1jhR6bua7IQJtwMIBGCZFQyB7Yh3ZZ3p7qcA6m8Wwt4MzB726TbruVtn2
0+7kGjJMj8TxWOg0tntAkPe1pZa5YNfspsy2QxxPs4BvGn31SY+Ad96KBCGKI4sfMftvjKjZGd+D
bGyA8Pbp9y3Wz0aDuCWMfW8Jdk5pCTEVhS9u2p5Ut8nvbI71HiLv8KdkTsiRVY1Ig6Qn2YeVHvLX
3fylpLyO/WwFDF9hmlPeAtWus7WGvDIop9N8dw2IK97JkEYNPMSeWQPWrzCP8M4QSQjRd0mi6cE0
mzkvBbNiOG5CTUzkpOPHxH7hiU+xYy8Q3jVJjLKmWomzfen61DMzJ+S7sM0rXQVK5F3KxGZ3czBt
tJKRYImcmuCqYqHoCJ4AeqLZrGPIa0wL0rKv2Wx4uGrWWK9LS4R8n6mvDvnmy1Xt1zSQbJncGRSu
yCtRgMvzUMDVXpnLOwSOIEsZKQHRqEBICeqqFN/hr0FOsgmEQhzemmT4kxkJEuJoi8vtEJMIO4F7
4iYmLBvqI66NuvhjcZUQfcM1OlkALkBfDYIXJ577OyCyTC2OKzLEuWWr+25sB240v5HtTscDHxrO
8cbn/ZYHTUNEEzujUvbA8lAFvypy/T+JEfF1Hb4EtLWh2PYijkhDFKuuWocZ83yFOR0mxKrpYFgY
uE61Sieagx5O/czYEGaUUFCle52cnr1eha/eW5JQ/7DF+9vBBzE+XaySxX7YVxa/WoSA+lwWaUNm
R6F78iNSqJuUJSZt+WH4qBd06EqmgzVA09KGCwW8mVVztJtfScPl2YJTDOX4nKiasbcWmbsVzdDy
4nlVFOtsCZ+BVXl3u8PnudrBOeYX6xB+oBtK+wDo9Zob8RsqTW6/O0CPv9NCm3euq0e52iZvQ+DG
X2t2l8MbqTXEGB2HJVF32oKkvW7BlA5EKMDl6Ejz1vyrZglX4CKT/KWARCBmvBaSAS7FwNagUwhD
Vb4v5dcHlwoPum0VHmWvX6IWBWBtrm9+bF+krpgv4MVbc3sGCu285hwugrhQgOofvUoLNev1pkdn
rzcEfZ9xfrx69qORR2JrmLs9i2oTC6DLXFV1j56AsenuipXHeWdBDgOno9ICDEmfsYr3hINKxdRm
OA2eiqhcb8bAGbsldtWVOIc+qq/DtuHq1mwWNMr56R/vwsY/JhCf2y5XAPFjOXDhs3fLmPqxedYC
BsuoB9vZHWgl3P3g6Pqyvu9vpZqvttl4qWCg+ohy6PjA4MUOgHZCPRF4CgYYuNxH7ubqT1Umwq4Z
ZR95ucEURzsCRUGi1l+gAN1o+NxpxrPGrDl9eIM+Kh74Slk6Sb8yzDFrFFzj6cn7rmJ5ZBM81uGv
VoYZg2ogFXRYE1b+ECzsy9PDad08dPT1xRSa+gYSELHC3v6fT4tyf/ZnTHlhM1LTUDP//NrQ29Mv
MlQSJzZBGNJ+jQ+MmgpR1bWKw+i7IOAFKtlY7Iqr0394f/OVr3FKmUy34xKeRPIj2P3kBhnv3BDx
DnxcZ4VSVS8LlPF6u09DorYGSdWENno83T8KsHhJmHdFB/juzbMhaz/GHNfXRViAPpoT84Cy0lTJ
JL/VrfyQF4y9lmJqRgEk9zoghMd1Xggep0o/IxgF6xueZ4otEIAtpoJHZyzjPnQpjeyF8WUfMrZB
c7BzxjpekCsNw3B21hMRrb+W+WF9vJrWhnHROsns5Ty87qhZGKwkcurR+zaG036lbkTamGpJ9GZP
hGgl9jXDNY/YC1WdeSwF+aQCtUfdfF+TFcHoxokL+ZAzNdHEHpV8y4WNGkp8eHm+7PKUMJy3/asS
BOs/IBX3xqC0fwc2pqn/bGEd+Mx7WJe6rzbiw5lC0cdqHHUl9f1ys0ng3DkYx8TOIRyiVu26ykkf
xQgcaV6uyV9/1B883jwopFVVp541iDpwyyn7vUTaoe6LeLocqP3y8KDAG1tL1QgZWLnyDTTdJMnK
m7CGCF5PFVAElWRkmLCdt+EsYxrmxuw0NKii9ST9U8JTr/tpdadzee32nFitgu2qFlSxOyR+i1Nj
0igXakNw//5rQLGjqQCstjTYifTjKB14fRV7wO6I0Z4QYbUI7OaqgBdX0oZEpmoZqH+RJPf1ZO8s
V07VgVUwAbAUhjnKIqBehxpMn7eIBh1lnGLPKIDH8nCw16610AyVgFpE9o1t3qjihYWndyYBK5Sg
0zaxsWey73kb/gVMjruS0TAbnhOHRls8uLny3/yHpyNxDACZUt3iZNXG+3bO/+0xOYwVTvs93bkj
JHXjcV4xh8uQDBA6a9XOqDljtc4E0/NJpKYAMqNz5CgSSrfX37CBKKKWGkVYCU8TnMqTUE8c+xMu
OoEd8XQcwZzou6I2lwS04Orlpl+d81EnrcTNLt48iDjzLx+wy0XwBrpmRANCY1jzroWjiv98wc+g
8HW6Mt0xATb8D/SqGOSluDIdWxAGyiJGG5Aix4HQ8/uGHNZrxaeOqz8IiMEGDmOvnaFxfJKB0Ely
93RI9kRufuDV7j5+CDW+kkxZn1JhsL+Yvab3ZkjxCdPCM0mrqsDzKt1gw2KUEv6COhbuttbW8u76
LgqjO/GQf2rnA7cbO2moWJrCnbb8f4QaXjnRb+GxxiH3nkr0HRHsox3maBhaGYCY7KStIl6Veisi
boGVUHAyNx6MITY1kGsiLcgTc8d9cFzH/m3zMFL0HyVAaj3PIt0CznB1GWfYcWThnO7+zPGWWLBj
Lc4RMbPRq6Ol2SmsV1qmhm+Bn9IFJup1zcVgQPUjdaspilkdFS7ojlwrcYD7dHfSo50wpFFljW4T
uj8UV1cmT1m/U3xShH+JLOpdMXIMKQYoy5mwReWki4MUm1uG2kWKTcldNORRbqegq5AVpGxhPc36
5RXzNaDF8VL34vVzqcZGCOEmh1zjRIBkSv4PKPjry7YrkXF215xBAzAZU71xYJBKLV5AJTl/4KVc
uq7cYKpbBWMCdb2GGmskXMSBnD5U3n48bl2JCBNxmSI92PICpPl5pWjB6tr8+9LnESNkITGNfUI1
dQIeBFZjwdhnpT/OkEM1u0y39lI+YgdGKKtMQ0my+c+GKB0MNxuKmqHqgX39w3HGbUggR305YUcR
IatlHIZcr63wG+5aur1vtV67Veqbd6ICHSDRQ2rA2w9rfc+ut6jJl95QRsPxJFB0pwzq/Mhswsst
/Rpfh8S5SLKwhVRCnHevzi4cASvyeJWq0e0yzl9d6MZQcaLMV9qGQ3K1lUi9bCaUlLMpiYACgWp5
pJ7i1dYNetnZX14wYb3gYZZoomK8nRK+vJ9vwxiePFxAwDDkm+v9bluu3vGYFNS/k9TJcYDA6c3C
m7sO4f+sPjKe/BEfR/ZzgSv5uuVrhA8/0klNPD7uRql/vUmy6d7zMYL/rOeqMvOrlX5bTnLE9VB9
jx8vSq9ox/Z2WUXG5E0Mi1hBMatvzCMSo4XMELnDEeF/A1KrW890rf+9jeDSKVtt8WJDa3TZOR0l
gaGCuVSS1KWsUSbZMgsfUDIx/sv/3Xc1W3pG1EwiICK+DfjSzDed72ow7Zx1+AzuZbVZMqvAWiVK
9VhFndMXrhXZyXYFkAbRW76sDWe++9hVRmw8L8rbb4JUpQR/2Kx9Xet1tmaravPHPMTQc8Gvy7sw
JQCx9VEdmHbsaWrgDDiVgWNtPiG95WoYORbgHI9AhvLoe8xL5OxK5L9Ox1WAkJxjsZ3ndnfVrnAI
3UifpJHu3mqpDSa8gs+UeI9kwzZ4KgvR8afk7lfJrU/X36TYF2ZI8i101Eyq8No9HIH+jrdTtwA3
/ke8ZSmiLv1Bu0jgrWxQ26S6SBBHpgYVOYT74pwUov6+jvRIF8UZvP47IZsO0J0mrVtcznjtUUVY
l03JfA8yaAbzZK/LfRWS5wvvktfU/QcttgsU4VKZos8zA0o8ysugPt+v/taWtfER9YEtB6dP1Uxp
ZGxuFOYsj8KEKWH16w3KGwEyKzYri4QWgeex+p6CQ898JSddYDsc9HAmHFuT4OL4qhQW72JMVeR/
tn3BZlhwX5ggkb0rRDDa4kLkCw2jTdLXzmoXG6VIWrrVFqhoBYQA5BpAJczROr/U7F4uTRjYO73U
9Amq1LSQYS0TnACv7FCCnAXTJgbS8BrkmQoYLAJUVt61L0sQJiN5SdGxr8mKxg9Q7z/PxFtJwYpf
ouchzZAEbIKtQdmIBsv8/IcqSse2Z6Esnq8Q3BjPmauL1uXDpQux/EETgx+bzvUakyIZRWb3QN94
JuzO9nWo9MmUnyRjqZfrLUSlzrkRXFB/TJdVVQyKRTMPa8wJ6+9hJbmiEbpYzFys6XCjelejI5gr
8mbG7DeQ4CGIVreO/Dr6MNFHVsAtZYshu0HAPW2eNAik9+Z2NcMHStnxONmHx1Zk2FcD7BOI3mdt
9INoo/BuhL7w8AklEGC9gyOLf0EfpC/oHlX1mGegbzbtUijmuukEr2zH5Cp3AyTjuUTLYySlDLIh
fL+lI29bVeIG3qAF8QhqMADSDwpT9KAgHIVa3dR0CZgRq1IZ7AIhQ9ysXm5sxZ+7Tx0aK9ywUlF6
ndRWhchMatz94CZHbyhetI/EnMCGoHYX1lAcP0S5ZaYs9zHUYzvEmu+A79dCU9q2iWB7uTNZ1cxT
yzAiAXHE1zRjb8Wq6X6j7tlc1H88JIhrCPHVc/CCMAi9zQX4CLHfQJRmxxiJwYMNB3uVS6HFBK/K
GR09y3NVqZyeu5968QeOlgWlKIQ0md7UtJbBkNnDOFtJUOvl9k7Di35idGZODoQMrW3R8mpdSXYx
3epNc73csYyFFr5w4aKUoYmjFWg2IrXhdL9Em5ppYsemR8FDwBMqWjSCgL32WTEnSRaKplN0iAp4
s4QZ0LzJrNU/mQkvQqoA/385Rv03xn8L283oIP60solDOKA1qXgO3GLnw+V5WD08UthX+9Ipd7LD
j1LtDevu1ShN+wFoBkGFzCExjKFHmQUefu1aBr8HP1rwoaleWVfJoOCfVhrs93PMW7yq2jGBFCY5
j7PmBrIvFYMk0PcgOPRwZNbw0AKrWF3a4sKH6zUZ/q5uyX8kSbD0A6gmyl78bc8nAoRjAyr2YpB2
BLem9/w1d/PcwqsPMcHaMDEob5EgFG4J5sgGhzPW6+KUx7yGNsknggl5xHEitTkYb0j+7hbWq93R
0Ya+47W8cgv5A6iVEfq+7XFd131KglPygYUwvashlgkxueQ3bdmhhNzPCbAfalHbX5VcwbfUHkOJ
8C9+chviXaL5BGaGBDWTqHYxKVj+pxC1s5EJdneQlkoAMYe3vykIdakw1ezrS0vBBKCjqbwPtyNw
ZAJBkdTbVE6CxIw0/bTNBwyApLW/M7BAZEKQqL9qdhWNyU2WlsnSkQNH1KKd40VNIg2JxOD6+WJf
CBsegr4rYB3h9TBKdacRl6T1g1SRPJscMthw3SjL8ayU3JxxajG0JmKRwC7nM3bfZnNYLcxu0u8p
UTpb44n5oafCA7+c3j3Ai9MnoDflaZjoqyffI30dU+l4YOfLWluihYgDUz4cCptzUlh271o3Xufd
luvO1xUYBo7dsvFh1utO4oIYzNmS2otpymJYZevhm8rfiQnxWzzs/TMBqa9vC2XoA6751gy8r05f
PqOgF7aBADMP3FxFQBaw2ZJpRFMwrFbKpElcY7NCZGvBPEQQ273lz611LnhwCuB87VXSrigjxWJl
pkNpk3EYkN/oh9wzpd09qvwtM+2z4bTrZ2oDkor7XoRejJuK9YXrnXxWi3f53ff8VJXMXGx4ny54
ClLjYW1scJxJmLoLnWNLzbQBRUyue+mzYLp1JkWFYD+IHUC/vm5cH0+vQrccyp55E19lhIj2sVTu
Xj2gKmrpJFXp0RNKvME/KZ9VH7sH4uZrdQIrQdOg6aO/irAYNZhNATEGqUOPZ+PcnzMtq+DFXdKW
hwkbefN8MGqnme9Ze2y2gT3PAtt0X8hDX9FojHCmokJjVihmzQ2+y4UQGV4kLvqHZ4KmDeZWOkeD
kRiunhjbUx7dSQlUlrRgfHGcqQbpbiQQq0SzUOiSto4TOaUhY+/iO34aDqJH1h3mC1xEq40Gaynb
P93IQ0DO6x+aePLv0MRnERZBKa6XLEt7aK9JCmuj0F5veK0bEKKi/clXcZQY2J4y7ToXkb7+U1qo
i6LQqEJ42GX+F/R+GF/IDf/U4hfvlSTngLAz05KJtr2uFB/6KSqAR8a33VxGo17WySYcHuKNsuOU
pah3uzb1VEiQbu9AXbIrP9dF2lE+hltI9MGVx7LalpYyYdEObCXtpzXgwraPrC+z4Tb6xw/ufttC
11uQ49/qR1ShGvED9hlFvznuuhS4UxmTKLRsLdCjH0+SdvZB/8kClekcangZ0Z9KZXZ1gUpl+Uc1
lXV97niLZZrSSCCYdDQI64mcB2D1sZWRhLXN0ukKB51f/1Ii1MCKjJnxZSqzlFBMtqSVJ9a9Kk9M
OJ7E47jxnthuwCN3vaUC2AaaCAh6vplmL1HEdfaXOKvEjAql5vQXb0QQIho9PGwB+OleIaijRS+n
KvitlC27QpJrgctd4QVw6tpljtLErbmLxorzDUURHtd75XwLSfE4WvHFj9QenQWISQxz2KfIJHY8
D6l+KubyQ51sW7Ei+gnyURSiJ5/yU7QuAVu4bF3H6ayQsZHW5+g6blD/4QkpuIIYaPCvz9h4jaZ+
IsBZ8pcvZPGjs5prItL+v4TUB3qSmgul1owSLciGwvANC3E9Vk1Aaoe7QpcRzP0ytf31V+QtRdDp
QkxB8ZMV1JAO2Ef4n6NbOqg7Wp6gTQXszrYq3dX0lcuFHbL9guXNYTQ0rlnN8vGtxY62GTAizqUT
z8yzRfzmkprR3kWeZLLSL6bJK32arm4DZz+eVP56/5lrZhFi6gX2+tmorG+eQHanzo2hXxqSg6gm
c0lsOdi/AR+YxKACsdfNZv/vcRB5Ao1jwEMU1ssjqPVPmzYg5icRDdy1v2/SJaV24RMKrTAmjdKP
ISzyv2/K4nXvso4080n68VvD41sj2XH/BfX4LvA9vWGGg/XFowNGiXb5X1mjGh41NwIWQpvoPAhJ
Y6ry57Ya+EpRWQ1QBENZ2ZowLIsNjefKxRrcmuyEC/trS6JD9jrKLyc3UHP+rT1/qqjdWzATh8XU
GyHhetz+9uvf8v72yv/27ik3m7utYt3l4C921UHh2zyaiSY4bgMHcDGiMir2yAsZPZs2623XxApz
Gkf7Ew/4P70f1B23wg9eJiuW0m+LFdp70sMNLedsC3UqiHrBRVEGTPFyUTDmTNR2KCHvDK5RWfig
O0KTu+Y2/x7wjbQCmDu10ztawQsmyGEH1F2UTAA3jcVP0ksYqJEbmYh0nsM26T94zxJ4jSokEJMS
E+1jM6BFeWsgSzD4/vkq2619KnbtXCPJkpSy2ZGNkjxaGZq8W4i7yrwAHsXvlHpZSDto4CrwnQG3
Tn12crMWunjd5cZiPaLL7vOagbQkbsO0bORLTASbxWhWvmGTZ6OQ8tQIr8oYGV6VbZy9tfns2ZEk
gqUG0eKxgNzLvNvoduq3MSjUYA8vCPMvHJqVNqKXrDfseH/rjRaSdwPjhmnP7DM2q0oWKygOFV53
ZGMR4zSqp8hit5Xui3MTvnLDtL97VKyUC/Uabyp9d8AGDhUm0fSIsiTqbwXjHtLfFPAtg/cbjjQt
1Cd9q6ssTMaNczjQE5T3eziHVpM2IDi4CEsmRRXfT96oofz3eaYkwO/F1nL25n4AzYG/JCGVTmBy
f6KbZKAVO3UI8iywOjsZ2Ij6+SElconS76aaOSJTuLHmERk18f0CjOEG0S96EwlcgJCuRtsZT1w5
lrLAxZh9J6X+EZvCvUKrgIA77+tBooHGhZtUGIqfHkkBCiJtVYGIQ/myx1faxDAtMHk7h3IMUmru
pmfsT8TG3FXrb0YMfCZgpmX78I+Sb4W2Iqcf3aw+cGMZnT+tucM9HyD+FWjAtFfJZHHR6eQKxqnc
eAFZWoEJlZGktFDt97KyjvqU+1ljLpC/vJHJhNAgADSr/W7zyHZ6RpbK4SJ6SDIkE4p1wLLjP15i
QP2YdYLKz5R5zJnWSukT1y7GvfLSBMX/ZXv0qKNnDq3UoBa4M5Rw03Q88cs8+k5XF0zxuXc7gHjl
n28hqPHmwXzPgk1o4TV99jfRqHEvn4UsyXcm4GPw4ffVG7AzrPTvXIqIiiRQY5vNOKKRl15IDNDS
FELyiubmYr4o9IN0HnRdXSGQu9Gwm7uRHjGCwoAGU3DhR4514my5d9BnBH/0KGYh0JEqDm/1zdne
ORfAZlVJ2nOy5I1lPwE83fmyLOeIx2DgZfNd9Yaz8gmu6JJBr5wULCGFqg4Dtxd2W/jfuKmhwDSS
edMJwb1gwMoKLNzuTqLmRZpCnK7ij+yBRa2tFkHsKCLyMUIv96iI479GEeLOSM/btalJT9ukdOkD
IU92qVUD4GF503gBoHZXDRtfnPJqQOxo7akU21ZA6zetXKleMhylKGHopAC4YPm3xSCL8tggOMpf
pZpsQZo3LmwK2z+7MXIPDPJUlCD0h8/b+EdZstj/FIuOQMpa9sKBKbhEGmzP0QztP0RFvv4DBLGi
mMCWidVlTwZmT+W/XuDDp0Orvvt5GM92aVtUAuG29zRyZSiXs3tHpiJKiShEeC53NJQrPLgpYgH8
GU6ZeDv92h8tLQQutTfmgF3UIa13jHMtyQXgJmkmfcz9nt3I3MI0UQ8LtpyqLFoPgxL0qEouX6+Q
5MKtmds36zsOB34hCSxYQgYDPlLg7IVZjex6REsodeyQ8OA+gI7qrkWA7xqFGGSGm4HyQkZjsNlX
tOxepnB24fLtf6tcPqI9SnEsl1xyE3DxL/DieF/jB+qXnYrSCEnhpMTiXE1SZsqHrPKUQB37sq0q
z7Za0+nmVxIrVZin4735Kkppsb94TVgcbtfsGbuqHidx3ixPydDsedaLeN85nWLR/6BJMNI+p/co
xxQsII15xsRuUME3HZmc5ZxeASNFUH0jGz+Qu3DB5x+ld14h8+dC323Z28Y+4f2frWnZbHCfbG7G
8z6PLm4o0aDI36fr+clyagh2AoU8einMARt9v4949yNIeHvdkUyYD62iNqBZkdPA/8YnVC5FBUjv
fbWssh/FKEo7Cnk64bJP69N2ON7hDSt8nbJMqWMGqoxulDdllImKLOytM+3VRREOv0BSWMdDrHUc
dD2zrDI0rAZysFJAWJVNWuyaZ9w/uGkj7UNVmBBbVlG5ZHOMOWtfztni+qgFYJl59ILLTVbcxMzN
gu5krLQhEtJC7cw7QsWPfDUXuLruLh8fEIfbk4Jan6TZzIEuAaDTSP90YOdY9CAsjd4T1ls3bxNA
Jysq1EZUCM27VDj69TxzmUyNJPconMMv0jKrLhYM5b6uIn0ecXfLMMpfiQUt+IMJI3rSRxtNgzCE
4b0+GDqJZpUgH0uopnAu8vG7UQr/9HMe1u1EDhZ2ARSHLzItYNyZaEpgMxdt1E60plEPDZkW+a1M
Rtsrs9KVWcnZQM2K9lfSniqnJzULjrOQQv93Sjw0CDEccBD09fduhrMCHWxKeDjZEhy+lW2mKyUX
eGzG8OpFnmH1lVGi7nNq3w7eymeFhGI7ZOxj+Mo4uQjbnPPdjh9tMrgnzhSA8BFP2mEpnbcWw98k
eiu0WrHuNj9l1DZ1I1WJe8fUwFcou9aFdkpT1Tvh9NPJZmvqC/EL9r/oUa/SRBh/ymw3yYzkVo/g
G9Y0Fl7btwQlxspXC8ms8Y/VUmNIrDw36k1oYYusxWy0MXZgBXOtZSh703+74fBPer1F8pzPHza4
3wM+WdiO8pYFkqVBq+/DNensX/9Ex6rPG/mqCE0jan0TCb5mYBBC3k6bf4HjmEBqngvJdvF8okRx
ccH/DvEH1ORURvhKXB5PY4xiTS9qiIcdxpbvdweG7qf57QgFP6OdGGyutoHe+aBKohfdTelySr+P
9rDe3ECGzddeo1+kCY5F0ZFQtEVrF2CPoR6f3EPUkR98KhnZv4FtPMGde2flXsCA4ffk7meZoIxJ
pCpOg41F4WJmOKa/fAXrigjqCrNkhOyB92BMVRX+sexA0hnm6O4nSHed2mM3b+RtSbnVc/tm0gr7
xTsEMs6+1obdFU42LgX4M+dI45KpcQrH7Lu6AGl2rTgFBDpZVe3SP02q+yMQkz7GOxsMZuOcrNg/
lskLudn7+68XmnvDn+doGARe5itWRAXJiAdGvElv1MNf30x75DfTsddHyOJPKQIdl6L5Fz9x3kfL
SSxFc3bfJgGhW7j71ImE2PlZmrRIP/MEjcMDWUKO+4/3OM+aYx0MRbOfhg+KlhYXHRXbtLYpBrYh
4ocM+GepxCQrd22m7Rs708bW4MaYmzFOnBIi3CGuOX0MrBh9Q8EEAHloTJj80pZbgL3K5yK0ItwF
wcIDSS8K4WA5sBHEBVLMd9x13RfBHecZhTIcbntJUJuIUm3V/7wDbX672ENHnw90CvpXkEmrOVL3
/NWBKXBoJ3EMc+zq+ie6WrPnitBQ38mFvn6smODe/81jArkKb2lGXYtu7fiCvye4nG9qLSmAzbGn
gEgXa522HgpM4o6rbxbXBNwtVmZ42HxomFrbqs/olDojZc2rmte/OwKOM1kx5yTETk3Ll4fAWrMD
B2yyJdbaesGzj2e5LH0NmvbqG0O399fsSbVuSJSFKmkwv90RnLZ+pVfUNL8dU9QfSA2bZEPaIr51
MoQA4kq5Z+2/EiiMYLndsM3TKiHoQtz05TzsObnnJ6Ww2AgVGexchAaM4kBnVK8DSPHDCJdswFKq
c6C+vLUhIME7F20AD7SXsJDA5tF29LRsWl5b+STsoi/3op/kLwsrXhFdGqV59QiMjuteEjO8lZOl
2bfZKCvP/GeBQOSCzJzdRigd1zjXM0dW0LpuCie5cj8tpXhMY3T2BK9TJI/QEOZh4CgydkI4EVeD
BZqf4KncAzR54b1BIUvjvPxE0QkFeVAaq9FrNwDsVYhASv1SA2c6KWORPp5hManJrg1jQ2Dkfcwi
zn+AGalhIF7kJziD4Dfo2f0Bomq2S00BWUpF+w/IsqBPpdbNfbLtFI2/ymgVIyLu6J4rm2KiEz67
2s4DqySCJAbOpC6helw2SQSNtQtNbiFOqWFqv0GBhcDiPHdkFcg/gC47B8kKgCb4ZemvlWdmgXxZ
LVE+2f8Eor3tzbW/hSsnxs8/9a83/n9oJC7sHdVfijA3NFgCjlbXMNJWuXQKGlOTW1LmK7A0W/2A
YjfnKsoobo/cpOse/j2v/gvGqIlXL5wdFYqyTXHIAJjw7oI0zp9vvgwbIeMzBbMgO3l5dGPpSeUY
t4S0NPeKSrnhM1N1IlHYLN3Vbti6dRmEVQFkUb4Ltm70Epr20lUqgMgf0HjuwiXvwyLpfCrTs3LA
XB1WVYsa/MlOOhPqWlRPQZNB6Ze+PUv1iqJNAyyodl2bZv3jWyT2GVsIaog4TQbrui8bJFeBlZK3
cHXOe7eVnAU9kkMLwCocNa0D7N2KC5xbLSTP4MjWOEjgFd+A/9Nh6D1zXBeA2CXhgbJAFICLgG2Q
ZkNveCG5XaY9hqUPYkRghTrnhAI9t76VUiWGIO1FbIfQV+wKDnq6RWKnF1CnoG9Bq8lTtQOKyuL5
sUH7czDNIDnaV1W06R2M/vkVvVqqxDJwp9WLGvzoKXcoD3fGrocUQyCDgu4RKcNnlxnsWQEw6OKd
MyvXEdEl4xqkicoJuAJPLEE80DZ1Ll4UiaMaz0BbM/Jvr/v6IV32scPQnqMN1854WJiqkS9v8Ca1
+6an621ZziCJifV0ZwoH7g0hdkzAxBHrlMY0q7LXe22LwDTzLCQrTR5I26e/7BUD16cv0EHG9Slk
NgPdwaV63oj96SkT2b6rLxo3feoA/YBd7dGijpgSIPa6iqGpEJyyIxTqW1CAYj3XzjDwLuTfBEgb
FNTsijdK7u25LkknZZuVrt54ozhdfILrFM9TYAkSqKOCWBIW4IflBa5+iXafjaOFJyf4+JFRLwPa
wolDUK/wtYVgEVyySmm/VvQAHSYWkiHsyePlyaEaMHhHe10ja1Fb0uVRLcISwCip7iINkgj3iTS0
c0Vd31lV0O0QbwiiUh6AKgb3yRGn9C9JBYVHvWYwwCeB6FYMRejW7l95a28XdzdzzNaTNW+2MJEc
6sUpJNWpkRJ1h1OXEeFg2cBuBq+IUN0PxWjpuDdsgbypk8htdsmSVdiPvFVSAicIecLR21PjT10s
v2qotZwi3oF6jhIVGFzwDWJOSJgD2rz0jiaMICTDqyM12EQ2cJXwlSyT11f61obbe3SDztf/OnoF
WEEYDIupB291ibs+Mog4jJx5pMw5BTrYRlt6fbWhYeaAB2iysjNys9tyRbeJ0eo36mRfp2DeJHBE
sBNERNLb0JhIkwSswrHtc1dJZMRQyOUk6I2HjBdbcpKxEd6kZW9b/IlNo77WKlPlpoxCvguO4CD1
LZBK7MZdjF+dYLGNgLhSEp7tIFDhLabspDi2urWSwj2fLLu0UoTFthlqSzbjanqZmrMQYs1gukCW
wGLoxm26MAS8wdUULcHWkJLXNYWgWZ4AnkhYVjfjSRlvNpiJCxuuKaog77CXWOQ8GRQ6y+Sa6ZRz
gBf0pQbTQ9yfnOojOorB1HZ2eD6wKR5BzzrZ6xhLJQyIvxmcbw83z0x/d/twsr3bF7HjBEKY0w50
KpELaOVeFJoyUlMfD6ebEbRpM9ZCIeFUZhuXpIHIdBqW5eopZkir23Z9l2ZcrXBS+clA6JcdZRPn
shaLgWJOcL23rVMyMV2DJkwWkQYe+KZvMgqtCQS//sJ88UpMHh+ldAEo/WoDYR7W+a7OCkmGsSiQ
l45wLquQw3IR8uKgFdIQLf8D4trj66nYscR9yhDcorTSLRy0xqv2nf0jcnxE40i8AqCLD42T+mbV
K1/d05ouhSDuaedja6g+A4eYzh/uRi7hWYEXpNvB0lPg52WPg6aZSbqEVjlHUsfgbGUnmF00sCjN
DdG5J0uJCurwnEBQcVAJbORJtT+mzrxyZQ3PpYGCIFm/zIwW6o7JgNv8jM0lybm1lmJvq4vHj0w7
9LiH1JnAv1aNuzuP5kSExDbmsUEn1WN2ib/ZW8pLNMpRcEDFvQzHe3zWqRZMuWu/RgFQfHC5UYro
+ccnp3EHYsp8O6MhjHCFINp+QFcaAgSHqd4LN/J7gV0jBl5+H/R8c77vh0khiVBOkwnC28pU+FzC
q3gFEVvOeIOjHLwqUU2ytoT3cXND1Evt0iyuvIk5JJBS8IQ3/ijJSkP3Yq692tgLv35Pv3jhyyZw
MtRk0HQ8pY1FRq0pHM0/7VsvZCg+zwQmrvYaVfmLVpF8EdlJuV3ZZGGqiPqbqwdkEu6kr3xHz5ZV
r814yQRgygElUzAEX6hS7/OY2DGbFCzyR/288o9/5nvbflCQvasakBHpnw0mLBpHg0+8ffPRef1q
79mddGTIzCOhuZeQNDAjAbTXbiYkCL9XA1azYHPSeyIln1CD85JeweTIqyIBX8I0qWja4t+sJ+t7
xof1m3wlrfooZ3qBL8lu1nHqwj3sjNQg02YOHWzq+DDjET7IMdfLnbaBRwT6kefdLw6nNUj9yxBa
IsiFxBrsjKLjSPXmKq2rW/SbIo666xIcrx+25L7SL461VHkP3bsfkxV/uHFXG86RORa4hwSxBLjL
5h0u4VHU5vKQKDOSDcI1kIXy6lWqlX6TY7W+Mr1IDeRTc3Y7wZZ+BYdBV0KGCCOKGi7tr101dljk
B8QUAeeJTXo9csF+oM/H5D8lLY2uyXVgUaCCXn2GOP/fzMg4uPS+80xCAIo7WwPQBEFlbn0s98QW
A4nm2jMdX3h2iyoYQnSKRNSaC0YYRnziBbJ8OuE4icN5XdxonqvxbS42Wf4VqDkgHRQef6HLVn2Q
lkDHx68x1wz+cLzq8WPUA+rmyyljXGqlzXpN6vicvO01vOzSD4a1KpLhLLPUhNr18HsDRdt8Tbgd
fNjKhVHEOj0dmXb6NE1SOG7BYnrpji6MWjWDwjcapOZZI3cbZbDruXcSXkXSUp/qyW3oY9vDOEBL
DAXA3er0xBcrsR1JflXT/bxcVtM0yUuXr+15Jit7IAmoHmqpr9BecI7qCUP9oifqC0ppvKTvuJhI
8+kZ6OwsIzz+peKrJPrqgt5S01BM5JRULdsdtRtE4EUBymbz55SfcIizzbPgn5+ljYtvZuOOhRw9
gA1PCIwANzjXWHD/QctFEJ51DlUBKyFk5MoAx42qLPciNS1un8/JMVPluJ86Q0B/lK6iKXqh1Ts6
QO5ZTktlCo37NkkF0plUdzvlgraFeiek8uha8tAucCiTRoBwPQDvHLB7jDDR8FJ7psvhrolzYNXF
mZ3oEijQBwzaErKqoaDSBPLiyBKfJ8Lp3QiS4Ht9kRpEi1iEOpkoRZkniTisOfixLF8lMhoxphBc
WK1KCaT0WeydAUbUQzv0bwCo0xdXGbqqmW73qrx+BR8Ys94PR++nhMxOh5zBr7mBpWmW1Bk2yg0V
9yefUOUknzps+KAWa/ypOtX/zgdhFAwWFEJcNbNRd3C+jFcxc8uVvavsc6yhNMLQfOWUJz5NfCxX
Modsz7DunMF+CT+PFcAgdlTYwKC177e+uGhdLK3nz45UfXbR+vEOMrqG6rGpBkX1Gl0M6rnLrLUL
kP1Nh9sIovdaUqBM7ZMW4tV/01y4DzZXKs/7+yvwRXaXiazZyI3srxaWEkxx+ljlAwYTA6EeEu+c
ruyD6e6Hhe6zFbo73d5Jozon0R4Rg2fa6EMXKfV0HIuEcdDui/zN8L4UkHijaghpW1+hkBs6B8j7
n0M1qex/jJ5F21fJeWJflCU/zKAnSI+FofYkieX5ccP4/BSusxvTAGpDtYhmd9d0OWQfrB06oVdp
wxb6S6+hbHwdOY5Fu+z9cfyzKVFweqPWgSpsp4EtFkpCf6WOkY0ce39KFFmNKs/Goz61t+I53co9
fpjKhPlN1CAXn+gkQLNFPNhSsCKo/z6rJfRIOXz2FomhVtO/JIrL1ISjXn0ZO2xTNbJ4824H3CFK
fHPiodMTqMMd29huqyedwItVGh60gBe50jxTKEsX9ID2q8rnH22mqkFQAOVI/1PADQMGi1icR7zm
yv3qhR/+lSx35kudWkiUHgqhcbvjgRL6A2GeQUrcpP0C9269hKt4PQCyWDiRrYNZXfM8KH0xwD3J
cFCGSH94ohoAD+hEO8HfnmlfGvw/hz2s8o9fpum2yrRZ7fjvqi6Hz+LSvySm6BOTLAU/yPEj0qLj
IlWGpKZLCis2mKgauCWb+OG84NfYwnlHt0dGtf/YYGxhRn00y1+GdyTrw20hk6lqL2Gp+EqKbT9K
gSIk1frUi59lMN7vEQNef6R1LkzB+rB0V3tr3R7J8i2DQ03lGhJhsNNZtmcvPJkDTha35ZDCHO2C
mNs8JVg1XdD/frO7mMMyP4KT+l4EZb6wOymBev2ecnu7cl5QrYiw8KVKseorpRd3NvT3TKySALVO
zAlgPYLbJiVpLk56Qmdw914T233op7PtqGrQPmVJYj5WpdEl1N2/clpRXn7ZUPeVLCauFjRzbLxg
d6or65k2bM6sJNzOcjkc4NQ6cJbkKp4937uu+ztUkyLna1WsbPCROwJvq/vRbW5KiN+8tV76Nf0g
keH1OeJocduL0kKptv3KcaBEWaHz2g73GLtdDmjLMg+7sXrFBxCxtNBzM//2+lRzMI3axohDw1E7
CAOQtP2oJ9II7XLZwLCHW4vo+56HqwQxjVpXC1utcWK94esoRGLeUcjgErFbaV/L3CWkrF5gjuv2
3f9sV5i+/n0YKj9IDr3YP3FUQiWkfjxvq85dNvEXBK6ewTbeKoWLR/E4rPOl+BGkrlj46iBOmTfz
ZVXLY1rhpZ8gECw3cKD2Wd0aijsfrNW1IFgODAfxbr1k8mBcE9iSXK3hCypIN4kluL+cfpWAjc0/
+fR9A1F8YYIhqedEk1c088cxEzFRis72qi75vb8j3i7By9BbZZzKQOuNIr1TlvcqZsztZQh6jbkE
q+BLsGJJQqzfPe24Fi0/H/V3WDS68JuSLPCXKMi8hIleVsU7bPqv4ORKk5RWow+59thhZJkiV8ow
ZFNLPWM95NjfV7cYtI+i8AbBFnw3eRBTpvc7ZeKcY9Hf/9CG9NTWWECOXr3uS791rz5EigbleVa5
I4sLwrCukZnfJZelwQhy6D80CimgZ7CwuQTDDdnzb9S0ND9tcigDXL/GnRd2lnUiRHTZ/so2hjDu
wVAs2BrKQGc9t3FLKFFYZh/UD7TgBWlIlOSDhuvs2uLXN7A5BHBZZhmsodTqNi15AstmJ455uDCy
6xj7BDEeVYsme69EjJPVx7GV+FydzE+X4aXhPP9lCsrEXt08AZs37ZUoRqM3QCkqztr0bG4hTkp7
tm2enPnnG2atS/EirqN8Qw/R27vDgu68XleE3B3Ti5HtMw5hz7zvdG0UJMw8dM4YknYktdmBAZ9j
7nseuMmU3vyRpU9W/xGvUuIZyOCJwhzPfgtpxPI54XCJjJUphSs9bW5qNh0Yn/d9wGyMQ982zJla
hqbb238gFArJa5Oh4V4WTDfeo+e5iogJdVvq5g5n0JKGyk2Z7lJday/ZoYZ+mtQW+X8seEfQAasE
iBc/wDB2cHg4nF4bQTFWbFW4MZo4kbZaN6fX5+v+s6ridGxLUR5xzgibFShHEipDrrmIJ4Ratr9F
Jj07IMpCVBM9n8c99QJBI+msHNECbnMPTfXSOphtCj4hQFtAkwsII8E/6WNFSnJQtxajssikrJNv
N7IOwyESQZpxj1INUS1eSOFKMkjTK1X1f4Eft1xhCjhno3CdK4ofbGt+lx8S4tq/soA3mibqbKJi
qNeNZ3jOrxjgoIxCzwsWyfvLI5fZhKAiJI17hRx1kaNHhuRpLTRABlp/PoyrzJAuFQtudFh5+sfJ
osPRmaMDX+nlY82w5c1F7pY67HETqQj1iSnKQQgd/bXm/17lBkDT/xzLBEH+xOIzkIhPbf31dHCq
Lldm+eyGct58VYIxsETD0EZ2zYtWXRprIcH9NYC6cD3vPzRqpOyG705M2JWi64G+lBK0K7V4XX6E
ztx6RUTNuRTG3rB+s/lw3gqLHZEkkQK4tuWVTqkd5PpoYjEPVtNSFZZzQp0sTVjzzGFO27UOPIGU
HRjOMtKhqdRQRMIY+9C7vtnn9J2hGyg57GYuABEmeZItxXgOx5BnaNLCiT6+wSqWa94vBrAfMWPL
dU8W++xab6QhBJg2kdpYkadVIepwq2m+5HpsTqDyZvj5kvtg9f0x0gL+TD/2fKtS+jlYf+MepJn7
0DXogTFwbTcs2bp5mntcR/xwS0WR13Mh9vrv9LlJi8e1sgj/uOjkvlSx6TjboydjWoEKbybyHeDj
30uu1PJ/brwAtX/N0AyBB0Iqrj6kSDxvll/Z+Xf2fC49BK9dO5A3GV6bOoYTaGbnSV19g0EnpLDF
+EMukzAUqeIZXykLCdi584wsQdtL8qbgU6/rfKhm2W6/CHT44ZaF8gCBSOZGpVfkNaXrtnAzYoqk
lOi1sQtXdCw3r4o1ehJOlnJkwlb2lDawFQoAo8eaSdZs3dasONDGzIbdGacEcjplD7gLRwYHlfls
R6H30g1AYnT4d18x0/nfUSPa3FkjnSzwqD7RSznG2P0jf7WJ4oS2/xyEzcuSwVzIP7+bGMauXE0R
6DHcJSGocRmTcpCIa2QiGxkj5mdncjvRoxbZmjIuqAHPTc0k2HjIpc7Tgw9ix2I8TY118AM/j2Mu
1VKvBdMn5zPGcOlsyYBcO9wzPsY6ikIVRpyDDuRTwt747q+a1MLHpwlWFvMQls2JTOr1sEs379uE
lsiufdSuRsLpwD73x5cBo2AY5OhOstjc/Qp8ByePK62EosHbikOS6W0YrgUVDeRmktbV8VYLC4x6
OR/4T3I0/7/V8Ql8nx+PmW3X/4sdVCe96NuRxdijiBeuyZLYn6y5iAbGNxQQE/x2wulYQG9g9Zt/
REckRc8h13Kw7WHH+ySTAcP7PyAz64Q1UsA3O4gGrcD+XXpd+UTGa4W87QibEYBeI1m42ejQxAIv
B2v+3czunzbtlCB5oBn/MGlJu1Fqxfgfi5d5qPG4GCFGKfKikc7ocLoTXplZZAR/5oM85s6tULGj
LmG3ZpTMG93PHv5yTBUF8/0z+Joqd/ewXsjxa3I8GTwyqNuBdcbfmoKIb0pJhPnhshHx+64oQvdp
pkPUeJzW0lgbEdrk9fLxDM6YJqdKqocinQcSfloxHYh2LC1dKpfpOgM20WQ1wdmRAPpJOAreFp08
euPM0g/bgA4aNVnh35qX5kiAPymDy5YOo8tSav3WsWzcLMAzq+Xxtvc0A57cQcu0HGZ+Hk9HZK6S
T36cDBFt9GKqkavsKQJjGSJgZv2bppbR0ZWrVggcZgEzzT0PREFDRro6+D+OmtIeoNVHIA1NgAg5
NH4p+A2aMCUss19gpNX+S4iBFtrDL8w5G6TlF0E9giVIlB6m2xyzX550iDaHLRJFtiv/mUZ1oU6w
vYRA41mgPOnkdKl6x/5k0+0kzY+64hUA50zfS1ylecF6YnSDMjpCnwSIq+Rc/G2ZTvz1v4ie2WQo
U/k0GaoSOAOuy2o3U4Z8dJuA9RpR51axjFrrDczOa8rRuCHCn2uijV+ecQMXjIlCoysj7JL2cdOy
J1PLvQ6tRUTJ8mJ2JJ9GILmpLpKZEGXF4/8puNHE9UtuCUIkKnwhyPvV4UmQZNsEHz1GvuY7b/ud
3JQK+E5rDOdG25O4bltNfwkHN7W2HFTC+GweOLkxwsX/NqvZoF5UcIPQ5LFHu+8USE/W6wsSnpy7
rqHxiC1pPAX4koXTlZGuL8iPy+hMCF7ymvpkA7NiC+/Z45CCU9MRgUymLEoHplQhoydg2bJ1ybqk
uUPM1M9oC0MJtBeazMFanA+r0/lJecotA5445DU3I1koqwjPsF1DQzLmMAS3IPuboISdocMWxfGX
wozbA/kO+uL3Ehj0vdpWKiPyrzH7XVO4I3ELmeOQqP/bnTKV18X97iP3po2BzgOTJtPQUaUtE5SX
YecM+6AG01Ie05RE2Dpps1QP0sbsmZglRiUuBEEiLeQtfB+xK5jXVyqBCJEw9vRhbplgvOtBPIQW
XtOHICeqxXWT9UrnYacZvjn8Nvoj6zshzR53vwDJqr+4DGSlhWnW0kKz8+3lfPKXGVE8rne1CW0Q
Texr1W2tdIcG9hnQJG7LUdPR/GLsF6s3FhGw1dMKLvjr4jlkgLQZs8eGj3O5MTtJJz2cZobsjeqf
aZNRdJf+2J/BKwuASTQ8XHPkCg+QBes4dQenMiGjAOJFqYJbYTcD3w/8lMLuVewWd6ouievxC2/N
t87PCn62IysQF15O7A+zmw0HWlqyLzqVUK4pGBurPKiLtdN6E/lxjeqMYqehgTECLS9EOX1JBXyI
M4qx1OD4tcleWfsIJYHpxW3Iqot9BS/mgEw87XvAsDnKFe0FMPdMbLkPzsien6sHp3aCvtMEj5CN
DDAE6e8z+5hwXZpWpGhPpb33YYXXZrD1giB1HGamJEsptRGwDn2yx39ikSWRH3b383k8zORA9+5M
B473Yw3KsE+/45z8rEty3JclXcwHSS2k/TSISBAQXKlIQFBZj67TZe9Z/NpigvzYy6Z1hq8J+MAP
HlCeqXQWwS5t0S3V5thTTSQ1NWLi6kTfHF2NTwWMnGv71HxuVU56wX9MVkFFHVSGsatXbECzuMjq
yAhCS6Qz/+JeIZykr+4vJZJYjxY9Cd1A+ojlFXkdYKqWZ0Uu3Iy0NAb2mLIDwVwTVVRGqx356OcE
lp2vfG/Q1o/wDSdA/w26tv9874ZjjHWTPQvagbBYgInb27dkZYykPyCpIQ4e1Eyimkjo7qDkbIvv
fLSptXa606EInRCVZ2arA6oYZvhnFOFdp+RoGAZxUZ2xvvxHcAiLgRgiBSFsaNFSa9t/ksMh8YkO
FxVMgPPVwfEPyuMvkto3AHkMDB3AwI254sodDD99/SE02NDOdBis5NvrNfTyXa+9pcFBzB9CHn/V
nCYXIepn2fOs0W+anc2wFLwgtY9yq4T+uieEPZBqpNya91euEG3LpYOPsuQa8xr80mhb/9wE3j17
yIYa/acgJRdKrasuC1jNsxnqgSzStLn2qYmYObKSpBLoI7dyqRv6XkqVMyJLtecpXagsOtM6eevu
k7GCAQjtzlPDDe/YGB1xkbwVQ6pwGp1EbLdfIuHI296rY6MZzyfi7J3w9LNdI+AV46tjrIVrmY0X
rw0wJ4N9xMSKsG3E2pjGSgd48p5UbbV1mcxbsNkcXSbRMu+7mu5HAjU7F1RS2WfflshysChVMBX+
EhNuolLf0t/P7lQUlrD8SlUyjz+DT7GJPVi2zSQKrh9WYsKH8XhRuVv02glekR7we0hTZQkpjrKg
sMnkgnQIy9iqV5YL6rF8M8nLMZJ+Hk2wbtvyAfNTcNxcB1d05wyBnTDeyaMCPFpgbYH07cXSAcL8
zA/N6ZgEyU0VxcXRbv/IgTOZ9fUgn+jGtIiileSak2V3/6z2GcwNqv+54AV6rzUFAPFgDKRCVMDK
7aIiGuzOWPMThURN4+lfoaopcT906muCsl8KgaMkHALiKi1D8YE3JLtpprk0l8+k5ArWwPZiLC6R
C2/VA+fI74I/AWvVhhPvOIHXgRjtd43pXJxPouR3Ono7d823HvGQ+IxzIXXo2/CEeVTrylEcRa9O
0SlvUR931Q49uKHgy/pxMpIF6ZVcmoQplI4DMZYDIAuAxinuBldOeJBPleJZBO2c5aobjav6LVt/
qbTSwpqyqHf90a0tnGrR98JrCtXLPLmj+skKhCC7Q3DxIP0iYrXeS9WZZoS71TD7NkVwB7UPZDn5
qvTsxElankymik0OOsSDRTVtlcbr673ZtXhXCi96PqXIP/Nngk3AAzrXSVqhqlxSU9MAxxwYyjiH
MEsyFnUgUtrd2uG9WFC1/eq/jpckyufB+6paDPHG1bpS1pTUs0OPi4mgwih+PQVOHH6toxLK35s1
U66jwaRG9pTTXpmy9Wt9kiwqeKkSFg55keVp1IUn2PVBMMa8bgseXV+dSa0gcB68AAU7+CcvzCAN
ENGy4mjAupKtneI9o4W8WuunzxcX4RpOskhubxWi9/Rdbw9pb8/d8igQn0c0cL7ZvXCKyZxnFqd9
AMv/9Q4OFS/SqQg3TbhhLBdrfjMPcmg6ZJxdX27mWExWLsLsalv/RMGisUR4xDmCH3oztmi+zeMB
PX5kTNV7Ws2Stp6z1VB0xNncNQpx4uTRZnx+YzMiFxmbmZoBYIkB6RY85Ms4EM+f5125hGL1uE2r
Ss6x21su/wrkYul5LnddvmWWQyhpRPMa9w8Fmtf6WgrjzZlTQd6Oj7t54IJvzpDxVfaPYgZle3CC
7GVPYsQROMFJnoSDpg7N8fe+i+b7YXkngw9v7DUrVVtnINvCffatlRojyLodL7AD8vAe17NOAsCs
Ws4wQaCPf0gimD1Oxqvu075LGVicMuiwC8hc/GsvZyNuV5NzEORgesBNTypdqDC+Ry+NPtwxmZ+l
6SpDFFJ8gIdRvRqROvq/2N02bIwW60OfY/7nDaaTjCyxAOU5z/Xiy/C7/vKjYu0UoUN5XLDijUlP
QZPz9/4hOmG6wdrzMZrRnunZc+iDv1m8vOHsq5Rw9aLJGZLlUkCcENZ3M8C6da5Mr9zz9oNfA05r
9hWEtp/Q1LfropOagtUz+7Iba7lERJ6r1ywuM9MkNyQSj3ybRZkzk8fHEwjQGhbNyHLkEil4Ozz5
qABJHGnfr8fgrhQ2gWz0XFrispIkuqv3tWZsGARKRxcPftwS4VAdJKLgsywog3iDW+s4LZkZaoxl
D+o6WowIMKchKdBJZMd8ru9lJAWhMTk8FE5tiRooB3ENbgo2dzibBvpioaewfJvHs8CXTMUm7bTH
cBQZOgZgFTnX8di4TkrYJ0DP/pqh+I3w/kfQk9SzVF1jXmi0rWGjVgBAd7xAs0s44yxYnvBihQlg
LayD/APjT45yw6wys8DhxhF3T9nzJHv8K8x+S4+gpbeiuXRG2cPUq5uFKFVFNsETQvC0srqcRt/b
qX30nhcZuRtcDHOo3HL88r8NQfmirLns2QJ5cg8h3/jXEFgrcdquS0S9ju+5a9rHy3p9Sx8PCPkh
UF5bTLQW0aXg/8NHeexEKUF0/dgULjnYIxXGZhTZM00LISBTWFUuh+uJCiVu7l+B+nEAR+aVmeLc
DfEvlnQVHpZ3WrcZL9jQ76YgP+OPy08+W3M4guWuUsz1RSOlt6xjfyjaMZ81zmc+pEjU5a9M6vK3
nmpuV2v2Mug30/+1IdU+2LTK9UniO4FnqDRB1ik8wR0iE2cZG9Bo/++pihDqFOTx/PJAITrSa9gq
EV9wBdkQ0xaC15k9HgItqUn5FhCBgXZITPpFwKuazYOzm7wakrNPO1YOl6f5/PbZ+LdmEz3xiK2C
h4m7WUTEzv7ia8Ha9bnUrzrDymsee7b2yVKoLLMyzF+CwTL7i/ShjOkAfb65q6iaUrJ0IOy0gu1q
72yEiRZtxOo3bJPw4tPkPLrgToR5P2SGqbdg01vfdi/fNIx3rVFo/AJy2LIc44+1PqE0BLw1sLFr
stbf/WHumrcVrjNdMtqohXMyfDYh7wVOtZyM4nOEf7TgReUUS/EZIvt/GcnNWpMjjJd42vzzEBYY
MKf0f5f+bg3ODyQcKBerURTSzw+WVHLntCmB9QnA+WxgJYMYD4zLZi9q1BfiFs2rqCeM24w8xgcO
9h7AAF61llZQ1QXJo0BNDqhsAzPe17Rs0l3VeelGg9rZsUGlHByRlLMXgtToiboxjHkmpO777S6B
wc49L5CSI+Fxnx3bv1GOdSVgWkyDvxnjzzBWWnJeE/0ZY5yMyOB0ChMZvaxb9dOxcIgGbyB1opPC
d40mH2smL0WNXOZLPDrLxBuJA9oECVdkcANXR4jA0vRRvsqQmsxJX84EYbKKSav/QFHDOq8zLKAi
yqJbXr0eC+f07COrNkgYzHetJdSJJVaW6dG0Fw0f6eSzjZ8XOYNAWn0EZNcmOt7MZXFEyiB1JopG
NrZ8+r4gYCt0N2mOZ3QWbCsHGXeVUnU6ycr0pRyVcTOXU8JMTESz+yYXn1MbO7Xf8wWHeKCJIH0M
FejyutYvk8a0hHjLNnCk3aUJGqzszPI0RGkGhcrynAVf/SYHsDLCY58fl/NiavS4ENrUnT40JcYi
wWu+OdfedFk2wnkz/4uJ0VtS7Oo6gGBx40t0qT5ATz4WE2EJS/WPPM9tpJM46vo2SWv4STfWfqFt
Q7NMJZugOL7kUz1ElQXA5W2omA0pzO5SUfChv5jKNonUSHxZsQll2wKmp03I/Tf0JUSrdRF9dyW+
s01w4zVce9IsuOZ77KeqfrvzDrgEl1q8biJgfyI/ncxLmCXlyMTyz3j5YiyKeMfOIxT9sCudKOMJ
DV09bqr6E3tKP/Gm40TBpxzKGrY94JlE76X/Abusy3qvSV7JsnJR878KHIEBrax98MbpnhRzZSHV
Q5PaPS+0P2wmgnL/IKbBupVuYd+nLq+om09ZQkpCNlEA1ys69544WvTJvtmYmqKsyjhnZ5yrcwde
NxYJt2H/UlqzXFCNvT5PtWUS94sbTCj6CIqfCDfSatS5m9UlIn2suN/rMC6oeo7opocE/kW4z9Tf
O4XyrjikekFMwOZtKAJm5Cx47VzXuH/cxSKuf5XqWxn1fQGnRs+gINsgFvDLhiBWcRvSV2hTm9Fw
rGd2PivOIuUOHLj3+FlND/Q2Xg/fsmgQ2yBVU+ip1X/4LFTPs2TG6nYz0ie1QUn9nXD4E0mOO3QO
OWQhS+o0ztNQkjYyakj+PNtpmtu5yCtxxumH3oSF7PVIVS/Pf9oVu0zsc1ky34maAEIygpJgeHcR
qviq81MJJBheLdFZv6UTyBh8R3cbS8KHsYknRphAINdyXXUubs3/OjkojYWG6veiQ9neaZIu+YqB
4d369YsbOHFrQpLulXQulFqFMExUXwJNJO/RNYwm8h1cRdqFv9mLpDGZyp+hYUHm6HYQAInUQQCE
D4iaZsSVVqUn6e/CF6dHer4LWNesvjF1N9r+wMOOy2nAPeAh9b7U2bvcwQrSK7LyUDV9mlQpnrP1
e6AqhX9u7GunolujNytZOJZoBWhHEX8CVUrBS6fhGl/JWqjQem924PDj6UB8+jZpz5RIr4XtGQjr
N0Y+5jgIffvbqlaVhR4fhcGEaut6Q9t3uWxFVOIYzoIZURSOVt0UbPGegbLJumRucajsdJEk+yzi
fMts4yNJz3uXyA0Y6e+Z0CIHrBTV0owhDSbN8H6B13cb6BrBiDDfDoOHUcknAeJ/jDfuNGxcT2He
bhdnDBRL+av7qnUuKN6tUd3AzFOTnaEuco01bMprENsGsThszp1BRxrDqYVXni+BuRMEPvO8Xl99
Maw81EIRsKNH3oa8GYuiu32Hm9jIySFxO6nP9KQiXyvuVvaXj9W0Nr1llGqolTeDmdJmt25p7wn+
jezPRj0qPse7fyLa2UmE5Vdo8JqvuKhlqQ5Cj42RCmLTCoVsMNsIbiIk0rHnyP1paY9rMOZTsW/J
0Moq3WDEjzcBzRCnLxULyR9ZWPOCPgT594JnOv2Jp9YszleI0c2B6oPbJPWFmDGP5WyH4hDWGlME
1yxjy3KWpjTm4YoTuDXzjyp3Qt4Tzh93qaN/kyrp99l21o50Yvc4ODtpkopTZSx52DD1809WXZwO
cIf7acdpzUuoQXPGczfXk84cDRC8tjkS38pR2WEb9KrRamCzOlCYuEFXxRXKlcRilCxoaDe08+bx
38FwDJ+jBXiA1eY8/Ng/SP9iWP1Va+1iFdnrE5bO/gAL1RMOYxvZOQA3OQzJz2IYU54C5XmEdtw2
cq36F2fJIc54I4vee7uq5e6d0BF0HpSWDyroSaqgaZzhvhWt5F86TE8pcCFFOQzcA7EkWnbEEERb
1DpQMfoD8K2PZK5tDzvntK3dH+bgi/qd9nopamu6R/RTKZa6+9KrIgu3yyLAepPUAE8JOOHrTAPf
J150qjX82fX5vs/CCyOmsHPcRcwoJF+jVNbHHZ+FP2I0zZg97gKGccVsG+Er/jbtv7PpSSeyambV
zvUBcHUsAJIDKDiWinpHZfMAoPcgjD7F5X0kK/qpQtE265pUdjoxP/grEoBbUViPuatH9vjITpH/
zgpoTE4PTnaZS6iJ5m6idhvSe828EBucpFxYRh9yka6hu8qWjQS8RfWKd4j9+6j5bXC+fzmeQlhl
SnNTKg4eRd9flNJnnTnLLd1xVpD1kYENlggoUb7/AMJd05geREbucMhFK4HFrWI5U4+yV18/Qau3
Qq5a/p+S2ySzHw9CqTrwRdQadDlPxwGxJjtqgX3EhsVPE2x6Gj0m2FGZXVD4Z0rMhk+uXBZBuqB0
KMae9TF4oNV+OF0+reHtuqYY/YZUZxSaJwC1lZn8o7b0UF7M5tPXr5Pn2K+0t0zZfLtrnSlN7Shg
Y+C6ob9kXXm3upOy4q12hAhLTq91lsV695LoNij920BGfNCDYtvHWUx/fs6CGcguX+GewvAGIbnP
pQR4Y2u0AlnURFBJlR6JKxXu/LEI+sraZtYfZbdw7bWNUvq8MIra1tPmeugSuDX0DtoKT3N8+UDx
29lpzb9GlJtvlYwLwxb9+elMgtG9iSBIn5y5XaRAghNfyZmBaNooCjAyIUYMJiSC/dtoiXoFVNaS
j3bs4B+lLoMGtdTRYyzHJzPLUW5aX0o4grUJWAVqXrJnNGdZfPk0YTBNYkGHtHSnVYBIWQ1fqTgW
xtB5CMn3WOBpfw6MGyuWgVrxdgoBJ5Y/8Dz4/3SxEFpB7XSXae+sWan55A32MD/X0oqBjaYLI8Yr
BG11cuj8QrKGmxkYyLp6dNMF0Yq4YZhFgIC0Bd1mU/WcQsl+J0ldjhhuGarY1udsSuhmc7htCsps
sm3SSOKgen1YMRjvyC4srR6I7HOkTgEd5ynPUCOzKUQeMV+BPO1ijvqOngXLqh9VdPBBRLRd+OPs
K4tmApqDEkw7eb4ZNu/kyf8c06cxJ+YEh2TnniV2b8HpB/cnUhzMkem/W1pxKm6qnS1HO/EIfAIz
Jb+0+PI3VyC6UTEuTbcZrRnKfy42EjXznPCWMm8DtuwtHvS8LnZV3OdMKq+iAsP4BC6Ode4AW7aZ
ZTeS7czX1i5NmneDfz0Ml2KraUnl6cEyd9yqx3P62qyaJXi1uktebaAuKJnzasDryiQxxJJWM8nF
ULrbBd64f/4L6b1MywS7n9ba6KIMPyaVPBwKX4Z7tWZXiKAj6e9gVg5DV1JmGDOAXWNVzPbmwAOn
QpIKJIknpRZVjLEVjcWQmy08eIMEKxLJVOllFmjmZsy/hBhDdwU63W1JL7TOSZ7dHT5jble9sPWy
pvoe2J+jWUoTSqqPgrVN8KXyIYDcJ2ByVrvIqYo7yiKyRh2tO1vYFZEZFWpbami/e9ppqzSbQ+YJ
nZySmd6a19jOey17LQTS+PWoVvPOYB4n6fEMeCYCacmhuH0aCg/h9PffUak9yJbE90tcVej2fEj6
+S3hvs8oE3UUh6gFWSuGaqu0QkmwWERMzGeJFaSDgc6KsDEBtKz7519M8RfQM+kG3AlPxRHEfcm3
Ocp2NafMd/JotzFuRbGEDb1M+2cRPGNSetSW7/zKTNWKRQd1q4nKQbih7XxS8W+IPi+ltNGO7KTE
KBa0eShXKtD7H05vf5dUElLgTXHsv67wmF+sOfDZucLkkFqOv437oBdB5fHp84kqAlB1f4z10cV0
YZ4wuYssAd3M2/5bVT+J7X63rNSYNBsxLnm2NiB+DoZE7cdZcPNZQwV5y759/4rD7Br2Hc5jfugi
rJHZodNzt6iHHmROOS5v+dDNfKjylFXlN9ZVllcfuzmyxhbKGcwR9hIlxVJBpYbbATFpajLNyI67
i7lBBe1HCgce8t3Py9WBIUxPcy2U8QTZKmzhHDQHAtOpW1uq3PrEEC78yVBWq4n3GfVbBF9BUfDF
Q/oS1ipWTt3zW7n4BdOZfRmO+flKvxtygqDZ39YIL5Zadl19R9s4r3jkRcAiA47fzLjfg68r2CeR
SkxsbsPag+jH/I52ri++ekrhWLbbVeaN5lgc9UdLnXw56K3HiEeelCxhVs/JhLURtfmZRzIneW5i
hbVym7fcHX/s2jBzZydyS/Zn0+06RfpkUGi33s+G2hv8y+ARB5TQP61W6mXGLvKB3k7CmriUY8Xf
a6qwQR23hZIPjaKsICK67hF2AFZgscHMPMqN58joRMsvVwDz39rqe4+JViFmAUuoZPeQ6kV62IBJ
Mx6FLhp7Sth87aL5ejAxnILimm03d4SSJfYsZJ9izNwFSZmUyQB2YfOaUQ9i4u+AHxrdpvAsnA5H
LOhlxAo8tLMB2R4V6OE95XLdA1cYXFPEKe0c3Vm4No54UflBTiiZ8wXLWM/jXwOP2fsLTxebd0g9
R4wyk5ASh2nd8gkvHD2zsWq3ZXWN9GOqdwc673/MEEmI8RfAceNky05RyIgO6Wuz7U7VRyozQtCR
hMGRItNwfPMGBq973NS/kQ7jqT2uD5HIIuZXCJh1vXOqKAuyJ6eCSmG4t7MyDbcQWz09WRUkClzl
rd6p9vP9XG6gNK4JLl16K3SuvLhDZROJi9Pqt+jLTzaBM8cE+PzTQmYVymxhKz2pP1FCG9Hfv8OE
mkMf51nB+OXqt/kuwr25AHwsZCy7A8QnF9qU9mHrrs9+FLJQVe5FUxV12JeIYp7e9uVehd+lgSja
aoEIc+V3/fULvoXHfS1fzTtD62g4wjB0qD7i5vGqYpj63/9yB8acHMh/anqXhGC7gF5iztprZ+up
tCQqbZ3UYoui9Tv3eCYOEV8vu2ruaveURvJP1QxR69ooqfkVZjEnAtqcsPhOK6s2jF8xMtY4DFDy
nJGfEC1TGIMeFsRsHGb8LxN/hOKLvBd8P1makdOlsIiyAA3TnziMT6s4sqCbAV8VHRw2WZ4G5JKq
hYpjop6VMeXG77zBTIkHB56I7OdiMBvOU7NfmiwHSh9423J9In0yXXBZ76d9ZkB0Z3/xL/2ZnFKR
/tEuLwfSoB708/BC4bGsun2iaXd579kKneWib5tvev60rPr83jDlzH/t69lDECeuRRk2piKbWRIK
Hz8W+0Irc3qcmXDMFUg4D0ZigLwDdmpZqxqp08YxAVm6Jm3Xx5fMj1PrpDNrI3IsmFFUwYlH8frm
GQwPQYzq9Jn1pVAYgUYjNyg1WntGPAdmfrd02FCski5yMzSiYcody4Y3yARSixiN9aUiQ2/SJt/3
EVgykbACqpN5g0rr67vx6rX0SSnWgzskD3oUgxaJfsmAJJQeEamzXo2PEWCZMW1VHbgxEZvsOnVd
j1CQAem9pW/ntPI+ncBtEZSD8zOCb7jywMrZRtnGCzbCIueJlUcz9ar4UoIPyykWJjn8o+65tGlk
EiGmeWpTnQkOXIHUG2vKEELFskIEXf6A/bpzCkrvisQUFVy8mpihTjqoRfuHcSqoizFBS+pBCIDQ
N10hIqLn9Wv0qcuTbH/QzS3OCH7sJZOWa5t/pQLIW0iL8NtEFwPljdCkqFZuVsgB6OgvYmbVxuJF
1TiYxYHkCuG2h55d2+k0n1b7YpqZJNJAoTdy/nXTJD36QUqTwJMJmNrfrn8ZHDWf/aJXJq6owaLg
0a2HvgO2wuxgRrWixOTMnzUh2ovgJQVPGty2BkwuYwE48PQNgjq1M38Zv0Db7F5xG34OHwHmgioE
V+L46msp5wX4hBZbXziROT7EHKk+yfJJ7W6lz2Z48ybwt/6ZXzDwUmAozjmWwj1m4RKIW6+CMAQt
g3ke1gVwGOM2QPFgG49TIs8/2pWaSEUImToqTwoRwIFZP3+eMvS9VUbQ5KOdWo9x5SoeFDki7Tnx
3yMRoo25kvlqHMPWdz0RHB+AeNoxP1QHEDmnmfQ4GvN3EqwDNZMMkfZP0LjFxtrgBw7MykbdVadC
U173ic5/pVmaNtIqtMd7YW9xI8IyopUeV1cBmjOqrfxOGmMyph1Xjryj5z3X0OlHUZiO3bNEAlJ0
XHK3lZSkXRzV0aExDFcKi93aZRp9T1/FqmYIJg9j9NVUe5WsKV7exfleIdUasC2/C+2BOn+t8qzs
8cppmqe+SXYwobOmo/n7+0DzIol0Q/IVy1duggxQbRvHBhOW/+Su5lphnGKsqlYZeQHMuTQC5ZBm
MjeIp/btjoQ50Eegcks0chtd/l7liyGsS6jP/asmC1i+ZuCLUiXUZVlfEkOldIzl5lA9D0ekY/jl
P7pw7oUPnzKasWSJNyGIL/Qqw2V7II04MCqHglks8sKfq0qQEyWj2K9A82JGunwwrB3i1CRRP9G5
zb5kYp50rvY53siXzkgPqRFcj5smBS9awwOBiXiffeDjprXNBlp60NiMHfyzDuL8GAItiQI5PLqS
B77ldcajrsAsNRTokqbqOgstrc7MTBCuL/TVQB5n7sZ4EnR9SX0Gl7tD77Za5YYAdvAKwx0EczxE
t/UFmHg76Itl8RposCHX9UW7gpgIJxCiTKms1SwC/oH2ia6R4u29OGvDp/iS1LsKAHsrm8oeAQ1s
gfUs7YHKAePl9rdIkuVB4U8PCt6vb59loHCjzQzYKXJQkFI14xiBzN7KL3+LZAIAy9pgBGO9SBjP
xSgjtOK2jCBINmOEZNEvNe2Cwe5lEoU1HkHNQvhQ38FdSeuFSjPJaGMwZH28MoiQoq0gqXC9BTZI
/lzTyEnWER1oye6OTTp+qbfr8n0xjql9b/NXDqJ3kIIfNGmULQg31KQGO2BlI+mQalr3WkXrp7QB
8bX2e3c5scVlLU0cfr5hvp9r1uVEXVLV3mw3HcZnENx76dtw6CZ27WMQxGMd6lPeubtD2UJoF6bF
F95Vaa3fC855H+VUlrTdF3tAcI9fKyALolNr0ZT5DjdivBU1IKZxbSIcYcQzzs5XTYdLCSL8lyzc
Y9j931SNNUGW/P7rOXaBXpY0NdRLXipxpctzG01uzqERlkCi+x3XgcVZl1+WzlwWVyzxHzdmu0X6
lnRDxu5DfDluOtWdwOKQS4qvSYfsUfhgn3Xn/lbObyZxAK0DZwCIo5svgtQbr2gG9owvsghvV7qc
29E9vH6zzP/B1fO9AgI2M3O64cSLNVj5bQHl99KmNQrZFlZijcMdW3qyXYfJKGPNyZ/F04X55XZB
W9YD81pvxMK/YwB30mtloJCi9nn1QI+GU+ctLjiKPYqJ9zkeYYlhzu7/5WMQuMeBENg9HaJybb9a
JprB/39K24t4d1p0R9H8jR2lKy3hViuT/Wb5GK7VqL3hBoRvQtef+mXTHNJalOhLzGXaSyOmTpr0
V5GIsIxyiLTUl91GMX5fMtrko6rSOlqyNhcEk54kaJf1NwR8pA/dsq2TV7yorHnLtGUfhNTDupQ1
rxAASsCzPsFA+KRd9Ivad7BOH/9pZRU2ycFbtKPOtuol4S+y4o/xvE8JqzwGFfmRu18xOLSPMN5l
AUx3tFtDYWRl1MCS73eEyPguMd8PI4L2cjcb6+nfnrU6hUpfyULUgDugkjcnVYlRwsKA7wH9O5cc
ira0zcnRMhwEBgozDyUGXKOLZMdN2D9M8IMRgxVHyaWKmGVCABMHblcbv1XJ43BaOp3Z4/DxyPdT
nQMnDHmmqjjkSNW8npug9Nh0mQXZtCsqqdWA2PdsySp7qv0F04ijfL5aTLR1VCgpEXpFKWMzX7Ow
a359c9fvGhBdja+XtQovC3Ui5Bz0XUyt6MwwBHCU2+7cG8lJI/wn0XzPiakl6+fnpOhBrb29WDIc
TonWhzjaLiPsQniWZ1XA3UVXtkeWn5ler5SEV8vYE9zrmRNq5boJ/D6nC5V2H1EsbK6aBQGsAOmX
uYUkOwd84hkhKY2R3YaqjowGr7XWx9/3BcLcwl1b39Q9ZaUqouuMz1Vk6ZjR37xRMZmZpw+uLa+e
9DoZ5mmzs/E60Yy9IQ7Kwvgpnnl/1S6O74lSI5dSYxQ14sAucvgW5DBkDHf/PMDwiwJ+XWfQb9/I
3ZKOejLaE+UVLtZtIJhSnCT1vVSUJJJebfTsfwBJJNIxT3j3qLIQyoGwi/clmqtjz78bi3XMdFZK
in22iGWuPr1BkWLBx48Q48rwugnP24BdfAVpaBLC+PnteAIp18w32uXNS8txtLJfZjhWBrYKzaHq
duHNoKZ9tvRbKUkwyPwuomy9tq/jdaqFl9AZ0PQkJMD9uBLyqjUVWutRFmzIpk4eEN1oxEm5CRC4
KdDdGdIs27uhVVJ2IYmSIvpiEUVtFaE1+gXDxq+Oo8YgmVCjoKB3OzxrMLckqSCeMQm4Z4HiIR2m
X+siM3evSWdPL0GISGhqSTjVRdRhotsDBFG282so89frMf++8QMpUNROvII+cYVnhaan1RV/yXJ5
5WNFb47rS741S6Get1ZBicHnHMhRW50Cjpe9cRIZWEMQmfg3x+A2l62Akdw77kxOgedKgGTXxo6j
TxMGfTfLJvNvLJwOmdHs79kReu9rjkmGFtrHehj7jcXbYFzWHtVxztAJTrfAQJIIX9cINhYFrCbI
7U10IqUslwDtC0SvlPAutR3PnZSF9Xou2x4fDjjjp+Rh25Ih3btqrgz+0Hs4yXjiCPQhjSz7Tp0h
lIMroUiGiy9dJiawYJOO99sJ8KTxrOvZeylZYcSnGSLk7N7GLw9RQLRrlbNWeBvI5+3GZG8Q7HF2
4RX7p1DoxS4THygB++OfNS+aa3tKkodh40tby6qCQr0pk4yaTn3p7t8FWn3TVUhh6OipLdJyH/ws
g1IrA+z9PmVSSqqW7FT/fQuFZojeEp+LHA8vhhrdKxpydPnYlwvjZfFUMQPpQwtCQQLSiOHe5WbP
TERR6qWV5LEKNO1hv33EaEB7+2zcVsSxU95uoKiUfSNzBhwMemFZYZ5qzlIr9YOh2mwD8jpNm24M
6IefEFdAb38TK9dsbv8/5USy91OqcUCKxAQzX/gmXBv43H/OUArYihdQvhaErvaneZSsmSmEi+zh
G0MTCsgGG6wFWA+2c3MyLoYSUjSClfTxucOKKUAoF4miQsAjLjkhlUrJunmHbz/xTQL3QgO0vtJq
uCM/y1BEFTNxG9cE5d/SmamtyB4aftenBQNS+Qq5tELFqXoMU4WPhhoCconrzRV5k1iiDDTThN7e
FoId3K7Myvct1Bzs+5YZVmFE1ZRzVASCAnFfu9xbMR/FngWKo2zJz4K1ee6sDHM1Ae4zjZtJVuBm
XWkPgaaApySMAVspRSUDAW6x9rS1jgplprtI7kMLO6PKEjI5GXSce9MnTs7i8/MCajNXaE7mlFvG
wleW3BZbRT/2oqC1MCTLJfvxRBgg7QfLvVkHOJY/fJxGUSiEfGUvYthw4OvXyjXNhplE6IVoJdlq
OfLb0eTR3H0Zx3wQd4poTMG6eMQwvEZx9uGI+qB5PWXdM78BxYPw1ezkJ6yWxCigIvi/WCrdbU3O
cylhBFRgYt3EAzjdl8k+y9GR7gRjcrEhyavwowqwF6dl2AL3F5A9I9Wovfgnp+IjCHRLf39QZibm
XQkdTz594JFnI4a/sQDXIqjWPaRzIdko7q7G9Ep7MKKWseUkYAf6YUTQBinhBb1lpUxQaLAtgQr7
u52vou1RaR5j0dktGXzLSKFvdk2TYhvWWK8ZvVkaWJ+dWogYee/3KJcYhxVEF0vL0Zk1G+KJgUn6
yF5mWU5WtR7yeFTkqCSzMUJIX0WTBMMPnbGQK2YzWsvLVq0LYAFKUUA+pRm55Yei0CzYE5BvchRX
/TlCKu+3L/iY0hd8WpZYYqLOxVNfWrkH5xUkf/3HHM96jcozUmkARsbjBGwxuuDjNvDz3toIVgS7
FwwpDpgDDd4gwLHCZxBZFIOZBgMrEfgltweuptKuOQb8k02fKAKAkEkiOchCm/ivXJ2MsxhLiYOd
AtotNdnuhV0GAtjqye7jpwBR2R0qaJuqzUWu3UPmfPenBcPvsMvBBpSrKhjLeEL8izgijQvJlJQL
1thUhIFarGS0sP+bavHKjaWPb+WnDa6M4ZXa/N/AUfKetvp0uY/SIJdbPge4O47rz8R95JB8IPh8
dUXgM7IgK8+X5K39oelkQ97qiulIMBZPLnA49SKIKKI+Y2/DPCBgZafTkjmFTuKmaCFWaUs3nCCX
v2ol0DdZaZC0Ch4pVs2FMq7MXLvz26A8JeCzZbO1WzBKQkWqLGTt0GsflgFAStmGpdXpkGwDFHqE
r4jfE/2P5HQykIac74Xq1RjBhdqdb/X1RtOcT3u1vKEZeLgnlefG+2CSjZusYdX6r/iiiA0eKHW1
EsOM8X0aTK0PE2AgqaZyIefrenQr1to3sBGt1iGcmLSMlvLRmkzuzFVmJq7csdxwWtxyBWOrH+XS
9HZPZ0in8eQXHABsFoD3CWDRP83IGo7KJE5wIoYOd+T5ggJLn/O+f8jX4TGhpKwiZd9jFSukFs8W
RmQd5dDUogT9Wh6TdeB3AY55ZxOLsOxnYKZ9rAY+Up7MkQ+jy1Q5+iiZwjw0sQZCwAz7U7tKMwGi
khA7OPD2mPWstYBxum4Jjhud22erNOIgykH7mUMJL9h+/UwCsNOsnUiZIwbqVImmdzSYbw3A4DpO
xvvUBauGqr1lj1OIyZxR9gr+CLGt9/+YTcikx1dU4iNhF3DKIeJGbxgO/sYBPyDl+Q1l7t0cyjkL
nGidgN7RScU/nAKXQNwQNH2HsW2+z6rChLbyJCveIzEKn6CppjKmcshyXi2m7kGNqad9MZm7/7Bh
VXiH6qmF3U7L3YGRa4lw4NZ7W1JcKxj5wdnDii57V5ZVtFMgEj81lg6BVRM+aRN5elik+0kH8kq5
PNKqWXRHjVT5PcD8pYh0ZKKj5X6qUywDEavQ1RDXXzfjCQi8bNADyFV/+x0Cxfhfrh2+XWlZ61iZ
SZEEn5cXUshYcNP/Hbac+wXWbnSQRAXaPTa5yzkSqAcy2zISUG3ABocubveYnWTCE/H3ZulkzdNS
298UBoltPVjd5slz7bMeL1QNDVe7HMboNmvkYU3+x6ZZhsVFCMcTgXgGI10lxhqSXbTPXm030uAM
/rCqc9Rv3s19apg+vUGOJ8eqn6PSgPHrKDJVh8ehc3+LJMqWOSWYR1rTOfJcLP9AX4aSuAqE6Hgz
aRX2H4mL1vNN2Lzi9ZSJbeVr7+pzbcOolllexScCfE9B1XkkUANLHuXUdDpD8Id1zzUXShIfLb0r
ke0yWWaTY0rIqrjC7bvC/QtFq0MMx6KEHkWC7TY9+5Ng9dgJj7xek+DDY4tkk1xftAVsZlo+kYu4
fqC2ky1ZTuRQ0PdeWnPq1pJgJ0wSfPVq8GnYGgUtDe3gb3kUlRUHIpO83oEibR4SOtuEmZzArIdn
xYNEgSP+S1/d7+zY127eoCMX+7inA0E8YHZ82Py3Gc2uGZTAo6htzjrh6933igPm7W9ShnFDif+g
husXuBb0dp2nLFsxGzQnEFoMYN8oxNeKSRvZX6eSMy7mMPyzXVYUseYP8XGC4Ptke79jlyvCCKfw
CN4Nt6toXAMzhtrIOgh4PZ7LsYb3E+LO0Nsq/V/dgv8vc9fWqcU+gbp+nbzsNYbdFrohw0QYtGSL
NBKJEkH9NH9GwLKw0vxhnLOM4JSFw0SGUgxYskATtjGMhXCEfrRi857E8gWZoyhNW8RlcFyhLXQa
Ge1jM0yBymtftSVKepcjfr3lKlq3LrJEmNGeps1ZdbnUxnImMSyyL1QYfAWrIypHNm0RzsNPIoaX
fTyzuUeX73Uyd4TEFY33Wta+fGwSPP2nML9gfPDtIiKF37WFPL0M623MiEuZONN7tEjOdPPPD+EB
aImcXxj2QnLnAwJMQHS/dHhAxzuZbik/pmXcJSl98iNZEvNUBZYd2T0pqColeQ6hHd1W9xCBkhQg
Sy7ET3S0bvKj2H1p/XksSGWBdE14m4pCpOAnPeFgU4mYYvHFN0p9n8MJgw7+Y42trND/yb9mKi5K
pij5l1d/rFZt/agbzYVM9oNy1X4vVbyIOUK1mx3Kcs80f7IMPNB/FThEQ4qiTVGpoLdklFNb+z2p
4WYvGx0klGY17749v3vRrnC//2q6Jr+4c8JdCQW6CJ8x+N7U6m1r1tUolvGCgO6ZsuWf1nQiqm1j
pwzUfjkFoKE7nRxjDRpzTqIoBKaw5oJ3Mp7aaxZXh6IkSNGmpGRyKddGkIsS0RQQVso9qUoJnvbK
1xkc1KNIIXqqVJeoHAVbwRP268+MjlX1cIMGVYPIKKepbgqrB3wtGGr0go5fB8DXVemiuGa0g3VO
BxX/LJWpyX6D5v3zLpXKWFCLjmbisFk2dWSp0XjFdHfvvzZYnzniUUmqHPe/ETWRWAEI6e9WNsTT
ZIocNyTpZPB1efDSskeyZEYWmAsyTIn5F9TMwjPPcUYGB/E36hPaoZuw1kfknZ51N9+DaPpIXCPU
eYcF0wOw0wSUNNC5U6R9pKNrhW2gg1R2geqdPzIZRN5Wd4MlxzA5KHjlwZN6X7CDrkdmpTaJlPrB
8Kf3SRnthLBTm89ThFOqWsNQhvSYvqwy9JlOINaGLQQoQRzG+u0H+CgHUYx0M5EGbxueYP2LEYwu
1kEL3zIc+6E1eTcXbBLvKCxe59U4zV4crDlCx0NpknTku3Qlz5rvFDXYjWDGJzbhg6oK5htZAsqo
mKhNi3arOgqdDJnAbp3N0ckEkw+f48lAc385gdFVfbltgKWtesmOkNyT09iFI4R8OHUUgDuVRdj8
Jmyoe+Tfgv+cRZ+uF68xxJfugZtVaKvMoRx0vIl+W/4NzlH3z/xeh/6sZbprEh5+DDAaQEGFzW97
qMS7wtNeoGEJ6LM0oG/sM6IlrNZNUHKJlhI1qyxf3qgXX9A/DMwcobiB0ffRtlAF/ud1Ha0pGel2
KAVLRcAe25W/Bt1gWJkJ89lWBe0pcN0lhxBEYbTafcNe9bB8nc17PEadlReE4AtkDK4rE4Up0QNF
wCzjvVSwpock8agyITJQOw/nYwaXxVaWaUzf28NW6D0yczl3dwXXL0aLW7WaJRTVFnXrMl6o0VcK
IZ24h2WeNeTLYQrE+B37lGQ+AEpQYXdmCPW3ixVr+6zmMGO6DtTpa3cbeUSPJosrBV5PAkLr39tv
Av/MSCyHvLNJ/Dn7mtCXE0oWGgT7eH9ckwzCOAmNXLk8nowzIqYONJDWN/InYW5hwc3cOy0ONdSH
QDrDFZ54wp5stAVtJOOVcllezH41WBConj8ZWXgIljz2VnvY7MrwwFZdTQ0bgFyOzXGLRIRu08PL
ztPzsdjJMLrXsmq8Af1NTw7UgKko3PXqFe+So3XzQCgMEQpkz18V9GUqOdpXdaPvbWQsJlyV1fi8
1ufshBrkw7PkGT/sAeuCLJ3h0CJiEsie1JfWk6OZZOXsUlT/vrMxPO/lR0Mkp/wHq2lcQsfpkUI6
7+eV/vvL7EmYBx+399Up2AyI109ZWI19t+fwTTYNHfFz6yfTvCHDMj7mslHtHDzW9xSrq5IbSdOm
pTOl+j2J4+dGYwS3MLhPXgjW/I7HbAL8O5+BwRe5L0MH7C5bKTSScAexW8shcjoDUTz9OW2I/Rq3
es1Dzrs0aoby8mo85Kyw8qNv6QJNFKCJ1n2DyNPpZ7hiF7kKW+GKZqy1USBojqU1njHuyYcUXd1Q
JMF8Vv0DrMjzCVNT3tl6pWEn5aYqti8/GgS8zpsHE7lA4JfHurSRINc+KGHdWcMGPOULjjyReNuF
Gga7z4vvacWhn1I9+XaoOeC3sHKYexjrZUdlpulhKAQ1exvMLgBFwOGi7LyQ/MWejmFHcMa9ZcUB
WQowNqMjRiMQER5H/t7BLVEnmfGIAnd/AaPkqMeUb2bIR0jUmT7N/+tqd0NdUSQGrl5ZpLKMTO3h
qSYG1Vjr046+0YiveAbRPGWeEdP3dBUq/z5GP88u2E36e4sWGRg0kIZprjKsj0uRs6+xzdXdsmui
wjgewAFEd6X+HwzHYJx8lZiY5DGQrpASSsE97jaGWEzwboJAe6mnYNJGXta5f9tx/bFRq2CEtRXn
BGcmXhp1j8uREJrxN77UaGiS1e1LyNYQprU+pHjnL5ghbIU5h36oOLcbvuAbqkBFzNVbttLZ/LAn
FRevueLzRf6VSZkjcrAn8PoMBonqekm5rocSnwYXehn6PEkgnK6XMn5d/I3NeCkkcuOpWwLG5otM
L9x2XoluyjnmWnr4fCnzkNsAR501AENvUWCK02wbePRS6MvxXD4Zxmau4QOhMSWI4P94+nx4R3CQ
QB3MRTUapvCO5BbMwIZwMmVMWL4ZFlIt+EaNENJuAsgm48HX3ia22GId50QpxFr3DzyMu+bjOtWn
fOOb9Rx5UYt/HD4PGu47av5a4CUlYG2AWFoIg9Hbj3aDVoV9Zme6/rjA9lP9VXPG4nzA1faTI5t8
QKpTD/7qrq9q/kTUXqmxl1EGax5fZMBHnWP/DcO3sHDnjW4/SQhLVjlr2XbZGcTEiLIIbiO7g17x
RdAAOH/87DIq36XpxZm7yc4/8xQgkY7EUGk1pn+yTZsETZs+leMERjKRnlB/kPb4DFibBxFCPlak
9mc2ZbNo7+p0wXDwi7fbVahj+iQUSrM7g/Zcrn3WmFvXYpEz8ca044XizxYdpUerETz1oZgAmR2d
2dieCe3nv7NVOCcZnmzYulr3L4r6ZAwFa8zDt4gL3VoozOYY56Ck8pqc4DL67TPYBv8v6loXbxa3
9FymvPQYiShTITULd0BaHfbVoLiSy6OUvxyDp4SBVVW/rXAP1s6mfu2DmLQ55SO4xc0hzQtiSc0g
NpmRkMne0NAmhD23UmVZ2Y1qllrqcA3DGf7v8ZOYKnGKs1Kuje3u1uJV66WrnFzxiLhNRQnJ69HG
5iLo+eoerTRR2vF0jytbOzIUtOl5RlNEZE6weBPIQNhQ/WnWrdtQPkLx3dU3NFs0OLz1LyLqddlJ
P93pYTpjEG/mZdbX8weCEMqWiKIG63w0O+hPoGm74R+o7AKQMCS1WUUW2exky1eg8Cv7E6xzCFBN
+usdtT7mOYgbO415zkw3QXMWehRd+x13seHjrwj7Y8kCVOBacCoZaprV5ZiSldGHTAYi+4wDDDDy
hz+n1xBD8SfNSmasRubOl1aOJu/7vS/AfXlPGNIshQpcIm47C0kLuwfqAsAeSq3F1X6P9DHUx+Bo
ScCbiAkHS6LhCA6O6thMc6+ZS3hYoko5q2dmhMl6auB/YRuG6y2f4D3FI/Z9wDMV4q74y0k9buZ5
xbWzjOQn879i3flPXwLZDJbHnimf162s5YEBQrGBF9ArDPp897SQeblvUwC1irQmrONCFVziCaHB
mIsde4DBliM3lkY4ukOlJno4H9i9qJiaTFicYXlByNG0KkmcWmTezu9v6QAssHWFBte18BvpEdSP
ahClmQ6rRiPnsXqpP2UPaTdNHUFersdoy/ZXWK4SwF+W0Hd3cXzU0kIpzZ8eJzrB1T3LVP30tqhJ
TtBRKUCRRtnG6Key2blOdkPPVV35fVl3jgVJ3+Wv/P62mgHCQqpKhdmnY/jI41nizz6txZs5Q+tm
5NvbSn0kzqp3yZn5soTzwMAxj2ZwUnEfZeBlBBYeHiqqEifKXrMIDQf3gTMaPRX9xgrly8vxL43E
wvhngCFbNEkJSgasByYaqYIwBCayWJUR2A5X6aBgW3CjuPiSUroqYf/zNM036mznYm4xAddDxnQH
hvzNIchIyS2ymQnC4ooAWyn/32217/aprhmSkYzN1BseEtiz1gyJLTWm+2V5LWY9cwyfEd1+raFC
3Wsk/r40Oi0UsPSue2ozXTWWLEpWX7HImUom89AkrWahx/rHRJooECSvvi6FnRts1RsmzQnRhv9W
9T4vZ/ja1FB4v3Cs2h7+WgTh2pCp+o29ZAkuRbqPJmCj60biaaQYzBomxDwS0nDM+QY6UrmbwdxZ
VdS0pHwbA1k+z/0BqMjS6FcFokKzuMiDy+ubqfhcnSLP+LHm8TfpsQLHTFyj2csiAs96h0iBu/VF
lL9IQuEkOMUgoHh5BBWRc7wknMUkJMuuL6P9yZRb1mRrrf7NH1XF0IiB6TV2aBLKqu+RkU/s/rFJ
hK+8fBdTeqKj4mUdVkFh6Q+FqfgP41xuO3PPQuqJ3h7hLBPdMtmuFJdnduy70BHXuWYzJuMsAbo9
EyoQSbsntD/uDAvNzqDz0+pQIPRpf04xnym+GzffviQqLJDaIrIpgpB0958GrXLzQQLIa3Zxp/V+
xg/l6zMlWctTrH8QE6kgXbheAjk0NT3SZ1G+V5ZXRAP9hqGvsOfN2lXyevoeofiL3rD1qi9QI1kA
msSpqPrtRSbh5+uSqyzBrE4syRUj9jJMtnDk5UOY4fJmjL1Vwuix5G8Rb3IcKmDuuAveUfiVQGKX
O+mRX0IAA0HED/vLyYq5t00Jgk61IID2lJ2He+toP8nJ31BgTiGsWGPhip/bFzdrH2ZgTXSbFDcl
O9kIwWlnE02c5q1f/NLelFnEEkztygL3LzlfJ3ws++zp9V2tdLGjz5uqG3tOkwMWE4M4JQ8ulsvf
zvOgGKzuz0RVGUfAMmHE3TYoivBuWBJdU6FywIgDcqik5O+AVPNUmc088aUGfSAh1NVQBtjRzC5B
qEGo1ts+U1iU99syxxVbM/5dVLmn1DkaBi/yWts4kH5IukCCxYFVf4IW4xlyFz3YnXJZZudoOsgH
+pVUW2WxPE7+gsEioOQJMzGBIylsc7aktiplpfj2JofYMYbN3wy3TWYMoplFa2MX5RFn1hoMPOQb
xV/Z3rg3w56wPDrzterEjcVGr9R4VSkHZgEIbx8tyaWa3lhLi9XxmUsRQ7T4hVtvTrg0B3fkYAs9
mt78sDbJr/iloIr7aFWo/sqzqZ5i3P4rpEkxYIczEhwBRTT6Vkjfnrp6WYsT/214r4tNwJr60epY
n7EylfAamU3y1tCRJnjTUGHvCjL53m1np4MEL4E4p8UbMPN/7FWHLS9d60g/wozFAolm49yWJx1c
me9sHzmNed31PHpXjNXkySN3kZPR22mDmvVqr2B72L8n5HBYq9motkSYIOXOX7nqRu+K94GkiYwf
D4eGpiGqTCc0scs+jlXDC+cTPdqZA8V5tydYuogg+SizN7PuIzLPwBx7gu0B4gGgEE/wMjffYNyx
S+iDBusgl/uALWucXAIK8B/wTS9A6H6SpdbmasRCNsBzU1k0C7MRLZ1VLjYMASlQV+0B5hQvZPR8
arMEcgrLkGn9gVDsr2M3yooNS6aRNvFF60mb2/F8FN8se2yytvo+bKfwvoHX2XVVDpVBhoi1lVxR
N1zOJA99+e+19v8xaocOuhNs2y8O0NlwhlXX+KU/+o2M8KLA6zjq0VSzy2MZmz4zZ6JQPFzonG8h
ok8v6CJsvK0k1L72ENebOgqut/yXEfBhixXOIgMX2rmssGUxg1uLY63RHw68SwhRYitx0vM9JSa+
ZIaGx5TYYG8nxD3Ce9YY8NUBZhBVBkOy9m7B5NQB1LGUN62cdV3b6Cs6d17Ym9WZJ0V8j4lsAwoj
n/9TmKRYBxovh+UTWdgaIbitONcr38gz/bB7Dm9BBiutNGlj5fqIjR7zyizJ4jH6uBTP4QOt+am2
jqKLxCZsCCz5ODM3nR6j6ZSU8Y8L/8iB5kJcZAswZVklZUw4JvhXUXNl0J398hoifRbPNtGeXFWp
Pi4NBXUyiRZO2Ij5+GXKFfmabgJtmpdPH+a9BeSrn6Y/D5b1d0H4cWU/wnWk2HSE7vby76+CCgvc
n9UroHHtN9Rciqi3Qg80AeEbIvwYAY7hDZ64+2Ick/1y5Lfsf9zvKZy82nXLleVwfpk4OnHFe4Ma
69pRlAabAGs/SuzFKBqU14edJcoLnIUwUQp58+988gk/5jFilc7hG98+gLJwiMTnOJJLUYDArP5b
xP34z/rM/4cU5udsutO6BqTpFvEjCzrZbHI1hasjQacedMwYoin0NakCf2JyJbsBygq7xQNQPMXQ
x7LptdTXnSUWXO8ieje2vsHwmpBkkEEmSARnfk/lWtZsnE2xFjDs0ro9TRYMbTpRx8n4ZxscDkVr
GksRJi10aT8UfE5o6oQ2hDOigyqa3HfE9fcfdRFcmmaYcknOVyThYLr5XVQx6ZPgaFnOilIuphE5
S5+2hEMNbBv5puCfomZUF7oTRVJFwunJqHWk8gCTTGCICRqWZxIlbBeoQ0/SlJcBG7vf5e1/LHCp
3JuFnGu+d6udCA6fowzLY1jCJ6Mg0+taxcDsNMy+Cm1fmSqYnqWBt9q+LN18CtV2H1ZN+NwjQJcp
wGmHGQfmTUjn41+xsP4bokzkMtF69H1lfxnW0ydglgezzkO0lyH76Yfb/ksrJwa8ZZAkDFnL7UaN
sSe2hWQpEwswuh+k63xwDB5YLUO/M75AFLmCfhJ3w2rcWqW/ip8przd1KAXuAjAd3Pecp0/TS5cJ
YSzQRXKnxn4Bu9V1BFx26aYu7Z3SwmS/paglJxRVV85PygG11q5BEys2LF2p/cm1PrIYnPBZrCns
JFIDtGmZg1XKULVx26ALliGlY5XRR5NSmanAPV8FB7359OaRCmcjF6SVJA1T1EsgxjTdBahr8mCU
sdhzSaAKNNZGLas+djO7ipjSyYli2f19lETSUflpl8bsZIIr1e+++T+m3oElANLFhbrtlb94FE+E
swjP6GOsJPkmuD57XJt/EBdTdKF2D5g9luOwB14GYW8roICTetcxPheOckl62/cn9SEghkPwzxm3
R6VRWcRRn/FOfsrgJ1/GV1i1ZUi5ILT5cw3QStCC/kq+2voBH/krxlIz1/Tk7gI8dwBqXrDGbJEA
7+4dgJHipwV4pxxxuyPt2SP2AKG8Bg6ZHsktvkWjth5Yjkd9vanh4GAFWw/RSNO1qVHETtzh/Fsf
vqRr4K7Gg2XtcT638tTGzF72aua9zmqiSo7kLwBIakdIs3etugbxg3oXxNEaDrE+RZxDb0k/Wkd3
h/x/T/9pRyasCgqzrSE5huWrTXLkLsIZF5w+6fbVhLLvLpbB8R/uM4/KysQUNTJ5sbVZrxZMyJc7
dP5oDIOoB4uWa03ZPjT14ag4t23mREPWz31MC9NxdfFacvg1PW7NDDzoALsNbw0t7z6zuVbUTeqy
u+AOZNsMkqpZY7vFWxUbNh4O3gZHXsH7W51BHjK5NVJ9YlsFbj881t/eVbta83IpyhF/V4f+PAFJ
rPMT2zKMM8d7/n8728PXgGcehrZWZNrw7neoKo+m6xbrnkAw5rW0Yvao9YqpmQrjFoRFqiMWaHBE
fBenpfYOSg5BFjtiHtCeFquhMOMpUPjKTehNbY8G+MTMCcV0hiyG8GASNstaLbjPXQaEvNGr2pWT
3B1zb63WTbOpSXU2K1geF8rZjJq88aVj9lwvxsq+FFa2Po4lOduX+juVhIDtWOCq240gEuGapaEf
/PlHHYgLuXWMqmIA/i0Xm4oAm36r2luYlfo55+z/FC/2gyoRXsv9031TMa7bGC/x5rJB3l1kntcv
oRHPydwnM4c9e0AOPtkJg/JyOaGtK/Lv+/xHPZWfzyS1p96EHhCTS+JopqYEf8m8OjpwZXjS76Jt
YvxzROqQo3KzqRPe4Y4swlwZPbAq58dcd+ALmNieJsBze/kNe6Jis2vf4n8IbG/7zuTQmw/qb7eR
BU57yihc/r1OgmJWJfAs5j8/r+hkHEzjJgQsumPB0MpImoSIvVfpILy/qBADO38NcaOrkkHFHVsc
WPRMq+mLhsyQqXzeen/fTkf3Tvbg03oKbUJ6zhtQez8zwyY8RcbCtqrTy3+JvUZ2co6TUYVHl84n
Yqu+6EQpIK44WMMbi1Tk0/N2yH1pM1nU1TsIGwpBqgnTpBidjeVrsCYe952bxZM76CW9i7eVAYzb
g3UZP/bNAPOTg5J+cbxIObfvCBv9pGncs+wTfO46eRrUvCDz1z2xb4Pbw50qV3kzcbpEMYi06WX+
QqnDcgMxKQ5bA03w89s9UvcqOOIsnnRe2wLTrHgL9q3JypXGwgz/6YoDkWFNPOhb11v93hDlaf7/
7rqCbnVTRim67W4glTv4dz9p1icyvZdIFJBYQIbiRE9YpxYMh+ApA/y2+JXnMbp9s4TAhzSJu66x
eu6WxZzbRk9UOQCBQKVxOgCodQNLQfzLsKhwigbsOhc4jUt5ipOai0uNb0MzzAS6B8EC5E+JTF6c
LzFLQbmhIhVQRdPhcGW9fV5aD3BPl9aUdx0CArS2JJ5qZM6H9885HtVCTw2tJMSKx3q3vlQy4UJi
oOossDmNOd0q6P2I2a3Gsx5iUDBxsFevz8eBg1IMAptwFNRyklqmLpuuD2a5r33YJu5LhgrIZm+H
3fMWjXJr0ayOmALUgh3SpaP/9KQR0C238jd09e55q9ZarvyLMF4/fFV/fYcn094O6BvPGAWKhc8h
lrZbZzRvuYy/0FdihRlXqdrgRVyL4LewmOcJ080cd06mqaH/h7Z0EPgXTn+Z9SuFy22e7ueo/5YZ
/CHhl6VOlR/ZM7gNYqp+cx5JZlov5kCkiZTx0ta1oqkx8ARtLMC3qmOm+TWAefdCoQKNlPEU5cmw
/s1cfciBOq/UI0zpehZvSiAdhj3N2Q8mzTS3iIYRzjZSZqC6me20YxgnEj8Rm1G+1xe5ENj4XvSn
bgc0f4/WmaEvwrFBBHD7CDvx15w0fOEy6lUlaEnZHKcJ6PezM7irhw9LSukUkVbX65W69JW2Qqh1
4oS2ykYTap6tCeel8sSeLD7HBDkAfFqwaCS8PI0RrBNP9bg7Z63lsen3R38R/+zJTzSOWAYLdcfT
iHGkrOQenKamBNJc7ZIUPOyqUM6qSFWyFSzag0CN9RgF8uBwFfK9uIyArsrJ3jKrhuVaf7060sI0
Bp0Ys5S+vxt8zk4H/2F8LVt7VGyafHTkHjxt9KBiFKLj0DvmHEXSoDG+PnJ6lqCl+WOPs3yQ8ay5
oBdRlU8G3d3u2XUtXvonnc+i4oCI/lMvNdD4fOnt8tmYPCrl4MAajgMuu1m8KGEmy562nB5fgluu
I0sH2+764Rx4p7Z5zm8WEGkut9RgNV3Hofar3Oi+xJH2GnikubmJi8L/Vht0OEZmlxBIlE8+Vud0
mpguENcBTpSo0pLv43gkz075X+QTPJkAj0l4bmkg1Ci77mlvwTZeJcAmcerXnsj0hFCrKZsGCZnR
L/f0Art+jpQBpYq+kh5DmmGZG1rlYkMEAl4dZ/uIa9B6BTRX3tBjRB5jTQ6uFHfiIkoWStyZCtI/
LrbBUm86SvBHyu3dJi4+mnCkTgImIY66uPjSFCm2zluPsgbe6lqLzd6UVMs3yKWTedb6Ui1yYUu8
CnyfbwYEi6cVJTeuHfF0lNEQ3ohMWs0IuANtCYyr9l5jXZCgU9j62Fiy73pkeAQJKS+fBUvJks0m
WwuIc22c04hXZZAePvkgAGQD6TbX+VgiM6QdF+NoADx+pXtz5/CDogY/LnxRU2RyxBma4Q188ku0
2eMEEjqWsn0d6MGzFQvHn/k4xAczUYXuFbbIWBeUbx0dOIjL/cbmTOI71M9l//LfKzcA1fMT9kan
m+MV/bYyoRtidNqWYyArAliL0JSIhMJn9JL3KuWvkLkQ5YNpNM0vLfJA3k7rDf4n7fy1nYgubTOz
kkH6dWcuiSCh3MiRFVMjuu0geggOrSW2JnBqxXhoTC6tZJ/rvqfxJbFjcdN41Is4wl+7JW309ZSY
ZY5orpG6t8I03s7h6w4LdxO+CPNvwb8ngk56XkJ0DeCLUlZiO/8vM9bjAmH/OcM5AwidF0H8zqhk
qNk79kl9/U0McpjOhoA67xjiA5E3PLCvXtbY/mw98avnY7fKaSrttIdn2jfEMpe/OrmeTHiQiB81
uXHg7xE3qjZGu7WGrzTP7x2v2bXlAqmaUFg4aHMuNyDmKqSwxwIxoKpQ/SSW8We0kR1CRv41q2Dg
0TmezDPPlXX2O3S+TcV+TcfC91M6xgUdQ0nJTv1ESXk5JdRwkzLoNPfBqAvHi4F68LqrXxUX8wQZ
y5viVWRpIevmkaZSPYcVn/d4jBkGOVuHVdhdMVL4xVltgJS9p+E5z42xYplOSb4DVah0KRSqgEiu
Ht102mAvNUM7/i06xLHBmDi+lPGUXuR6gHQy8sJIM6mtOveZ4s+oMVl5ynUPlx8uQ3ZA67+fnsx/
GoTvgdBILrVLkazakeima/hcu+wUW5onFhxKkOTM06mDnTJiVCOpEu/3RGJBmLk+rwW62wyMdB+N
NCP31rRkJUq2d5S/X/CWmfB0zae03euuAvMdCpoloDezNMugOW2xQM/UZvcx9KlfoJ1eGkzzaC/P
nYYezpxZ1OhqhVbCjfh9ntwgjAnKtziDfNiPsYw7U9eYfNeHyXOxwNaDK70tNyk8OJkJl3dkNR/l
IywxEn+PADa6d5YRFCrnPfdRMc9qF8gK7XQSviorTCW2sv2orpDuVbK0ImkjDB08n1naDnnR56j+
RqFLjADFHt8cphyC1B5gULJiewHOw6IpYKybcJ7HnidpByuWbGy/QZKXW4UKQ2ZkwVRSGxh57mj6
grpXeQ5AmPH6GDR94cDMPrXDsxevh/j4jj+ikHJ8paTq2EsFC457uLALNmNu4mJO4jYiOTCaieHR
tGgjIUQtqSsnHkLCIXCs2iTHWs3usY+yfzp1t9Sut4CkXxHj0mbmzgwPghux6VqLa7BUFG3b+ZIW
/DZHFmrZFL+NcipQgBqBZHpd67lYTFTsg/EPucognc/f1Ttnrg9CUadqhwB93VM/U5C4ro+KEoSB
AiVypS5i97eIGdfyxKAewtn9v9ZT67+T/TpkUe9DWJtzjwgCQr0qAIQhWqQFdnnDk3yDwOETI2ul
x13nAuo/hrjyc3HckGVEegxZ50+bnrg7W5IDsNMBKZF2Ue+7kD4Vlv05VmfYnLW7i+LbJCPabOvA
XYalI6BjlngxVSGfVZrIlQopwqExZUU35yK/wU7WW2eiHdbgP1pTRRfm3c4SHAcNuBvL/60h6tA+
5IoDUeE832NwGnGPgyX4XNh7bgJqu0hmpBzQ9kF0Luya/0RJSiZ83ZHnk7ir0nWkS4ucGI+e7PS3
N4A/6LhHmNkLGCSNvD0W+T2lzQXmcCMMHquZ6lMvARooe0NMcpT8ME0gWBtDKNJFU6iVGkie2Rf4
NgkYBJOBVTycFDaknBl1GCV5F+S36iiZL6/q9yHylieo4IbShPgGS48phHu+XShtUGS0ozp3ihzm
GpxKgC/Z21H1TaknsPIr3l9G3fbAw8+gDMowPEfZn34qcREdxSdtlyArQQQIo4sTy2eNsgY0UDJ8
kHu4TU+R8HrtaISU4D/WuiejCzO4CCoQ4lnCl/YFW8Wz++HRld2JlouScCLWgwQG1zwCDbKsoXCe
vDsc+AlKxEra+C8DRoSCFpkw3twaeVMJnKuEFN5/WUjBt8iMfESxL0MQ7+Tdmi803J1mQ/uuw1PJ
oMmz7xY1eEK6LuMxKFBn7WafopnvAWT3J0JGqth6evS0phJKelUmUlkheRpe4msvyy02gR7NvK0R
BsnB5mpkTe2MM6LyGWEx+qIsI7r1Lv0QUTV0ukDMi7VqGjjk2aQqdM4Soq24f2Y9IdQ8ZM22n470
5khD0tp6g1qncVVm5Y6tIicIpbBXhcYeYXAC91RdHfZ8h4XoQdg7T+huFwVmU4xA1aTRyU2pl53p
A93CFxD/UAD5HqfTtaqPxdUuruCToKlGrfZoRNDHyt3DF3B1ACtG/W+9aG56MZzdZzQTGgrIdK6A
ghpAjrC5kXblk1nLgYPmwQt+UcpcWC8xyXc3EiqD/uTa38EjEQ+awU2xkBFhZ4GlDJDA3UnDcUFx
RUXvb8F63H6LJd94orXPLA2rQaJ21eWHFn9C7c+NsZ4HdcQbePtza6ZCnmSeR5u8Ymw+knuO2OBg
VbsXZDEa66wjfVTxfpKPw72kkOBPWpK2RM6hPDtlrau17ZEahzWRuLH0TexPvshZ3Wbr+j+a2TXd
nu+phBMx2Bp63WZGZg1tHdOPjMg+Rnx/V4f9RJWL2bQ2uEzEu7bWPj00sl931u/VylVVp36r/MNP
b7br6iVDfEmm7t3fbv9gAJBgdAgWypiXJPMYi7cdApYpa+RO0Pg2VMnpIt4x2pxzsDrAckzZnmZa
0aPudslt5YP8vebMk5T+IMvVogXsOBGw3BZ9gTE1m/nxL/BiIW5gEjpg7P3z2PnovkbiOrEWJcL8
T0qFEDO46YmJiidR1FZOAajJ/BoyD9FuCkIzUoRb1+Dirf4JFqm3MrudgfbbAdQ/hIzyZN2+SwPZ
dNKuqsmMLvguSHln6++he/xoxaRoVBCDK8vbFmuSN+egheB73b5YhOdXky/xYCEKXdAZusg232vP
4Z65U2cFDu9+nw5379xf0P2kJLKYGUd+/vaiDErXdVjP/NTJq85hgeHNXDFOzHTn5xSmeEHIny+W
mevLtGPiUf+MPC0PK9XWotuTB6SSJfrmY+EQLzEdpt3ADqMGNYdtl154r3PFG/lYj3M+u7wszLd0
WvBSDncE4oisb7kV6k+H9DpgSNWOzdf8KNB7B5e3I2pqePh8qotyJ554eq0REKzbNU+3BEABzm/G
9VwFjdoNNlwUtn7RBzFTgajGVOybsuzUwr3i9agVlzvdcXcJxxp7Fr0P30pdVDcFU+I2bJM1Q1k1
/B4GrAMgkNGIL9ePXCBETBTRE3Rrv7ABFRJ7mNuCfrVwI/SZ1bZFwbsPbNGkkxOFKs0dOPDCO4Dq
T+DBELgMdE3X1DWpyPZWdrQyY56idujWaLsYooBTEJwQa58GRoS8goQY9J6TqRDxwJnj7uQStkGA
QWf2wbJIv+wlsxxn6qEHItf5kIpsrfB1rHjO/fDTL3WLul6eiig+/iVhxqximNRwy8FCbYTBsQFI
2CadS54d+HkL/6biDs8zTUl4D3xU5B83AkONpKzTqa4PrTt7qqWS/Dm7xRfsVioWsc4tHi97hVFd
OjZ7hdaLvzETaAYdljHl7PHyhA7UYUMydRrQpi9ToGGkJv5syp1LMIUJSc98FcymIuG+ATeQEGXC
5SmUNj2RlBlXeZNTsusDCHgp28qQQVjtTAHyi1+Hv9lvQwcms8pXgMHNiEFPSzUiE/KhKMG3BBfY
L5DRnNTuF/jYpaGtrTGSrHFTqGjo+emjrLvRZ+7PEHY0Vvb38HFCAcMNJ+LSK9Owl4Hq3ecNj7R2
YSG5kK1NprhNwPQ7eLH06WSO1Yuq84mq7d2x9yR2iWjAbDcR8QwfbdK3nnVc9G5XA8ufmiQl4cjS
oryg/vjjHBYpLRbxOJ7KxiJHv5TrcZqYqIruNZKaxhg+LsGLdXXSeudv2KEmtjGZQ/Ez5hL1claj
SWmnM4SVTZ9MZYtEHg6j85rK4e1tXBau90cmnafMkFp5iLlNaQkXerDhDShZ0aj7VDl3q1rlyT2u
yTr13FZ3RFSaBz7OnoEYHGSe4rlXJDhgWTH5/zLqU0DtnU3HOh20KW2fQlDm9ytmITKY9tEblgOT
yRugiMwoJ5cwRQhMEwE79uwD8fmBcaBhgtQzh2nVnXI4zdW/kQIB39zECA6Xa3jKFjLpowi54F3k
vT/e/to1+ayq5AlwvOTU2omNRLdsE7isq2zKvnhUUMPUB8yM65X7FB55kDa7a2jmeyC1Gbva7T3B
rIjp9sl5BjuXWLProL9/9ySflDQcBdMh6gDzJ3RluxbgGSFMauiFiBEimwR+jtGBm3ULU3+Sbalm
7n9Bjsub6S2v8UyE96PcQBtQX366X6X3MJMxbPs0nkrnYQ+g9gj+Nbh2CTRHvkNTRqLt4oRZ0PlX
D4+Sm/zDv2EpAr5sj17PuW2wng97sYTK0hsQLWq8VOg6y+cuUadYJrOvkgTfW2YY/qt7/EhDxPtW
ANr05kG76XKK6T7LN4w78GLs06yF55bHuxEgvyD3vHiPNFge61r1oG67T9/X5cbr43d0lRDzSnQP
HrGOZ2clVSfCe9BRc+m1H3FuVZB+R4o0kegtPwbMFoo3I6URTLPVHwNR+BbVHorkMoIPU5+/+2it
XRiLW63DGNhx65h/JPjh1ielbfEUKANdjmQb0OHrBjMYS6QlGrt9C+QDOFOzW80WFvKzjuFcqSos
R4F6w2RFnrKrRiaE7ovX1zvAgJmUsjVO4V2u8nlEHw+yHbhBPK2ElfoB6q4PyAFBCH1Ubt/NL2vy
R+QCzH9ORbIhuc93LSkFrq05irLiy044CDegrp6raj+neg9yjZYUfgajfctHk/Cxiqy6EqOZBXRa
zWQUwvNZfbzfReCJ19RyA6urMVNT+mzvGeNyH6QofUI32C3HrVU84ZyYauZGt5PNmwbsYtXMp4kd
cXjMpkTD50htphMetcplJxfcpSru6/wMegQ/Etb16BNrqVwizLPfJ+7ticYZRZ+QLj2K0tVXXoSK
xRcqSo4tNeGQ4o7BzZB6h52/jZQsYxugsOWoXopMkZ3kxR7PZPRiy79svTvMk95rYqdLdUEVjqKY
GJ7LTJbn4Sn/DWbCJN9wF+AqKSJnt2+lW1rhsKhwmPD28kd0HT4tnV3nQKf9zk8Qq2Br0AP7amD4
O2o0zoC7PUzbbj0vk1I9Tf7H9+I28A7UMlGhveKWQD/RJdasc0flCjvMYClXTwjkSQ23knaKqHXz
KEy1AMd9uXJ5CV/7Z+oUg2jzE1n4og16kHH9Jl9gE76WP7MA6MYu7E8hG4mHbaLnrlyOiYgfOJry
4UvyfdqaRSfuvWcnOrqquNf6YaUdDgOq+Sn/EdKlM+Mx6SvOOzZc363PEDedV5fsWJM4UuhkKSwa
o3nP5ZyHr/fagWRCs7sw8zKPPuihAdAb7DkQcap+hPgVjDwRO9pLhMztTA7US1MisS3EsPH5rQWo
kmn9MkE788M9pzKli9ZQL30adYao6nUY/TmZ5/hSbQXU3tIJaFxiRQPWW0agkN+o5XRsF8V2tJPx
WfyfhZa88nrT+6CcyzMrnd37TJ3ywuZki+3bfI1tNz8AJ6eEK6g0Mh3lFrcbyjf5Whx9IbEWm62B
sbEnrasbw1j7NVlYynV3SxCKURKjyjaDtuI4g1Y9nrNvng0hIj3Wz9o2FofkkAkZPoKWUyknC30D
nqwKjPlDdA3GL/dGfNR3th+nmw1RXqYB978bjgmIRV7GB/YydDpWjD07AP7E3SE/JtzGekfQDve8
66u7T1+bZX0ZPSXrNW+voMWngE+k0+kWhDu9bIMYDjS+f5kMARG2iqzRzQvpUWBg5w3MTfPjciue
5bP+S+XH8kQcqeSeHjPxjvyFrAzWe6tyqu36tbMvd4r7xL3ctcZSJ9QzfVrMQMCq83qLpxf6Ue+9
SZJXV74YVSnK9GucyYSDFJpa91ABrTq5OGBRYctwN9ydKxQ5+quymPCZKKpFY7cdIH4vov5jki9u
C0PXixJGJP2Vwz3IotOSuuEPS9+tncNkKQsEml5vWdqAfD9sTumGm2LNOXLOA/nQLBC3LBbEwYyf
4TAyiqjj6Vi09euw6PbOa2mvsVFZSnCEuXN0V8+kDRuki8s0iJt4rJp6Sb1FNwjFu0f5skkRzf7Y
d0NuX/yk8mJ+cJ9/MHAIl9k2X6GBx6ntYFho7x6e8aRJqhgKbpqmNzKLDwaVToCjJ2z81fsYOEhJ
ocAulcheuTevB4BHo8i5UFpRZF5I7H1y8ptRscdiGP0zQJMVLiftvXsVwsMV9De5G3f3+lQhgwmn
ApaygaIXQf/sQq3gmnzxMWiZXYxMgNwLDXBqg5xXqrFZAwsZ2Z4l7La3tgkg683Bv3tseGTAXigu
7sCqRXqZRWGpOGwbRj2My3C3m5FlGv5NenUrk7PcVn7mPfNnA2GTR0oSpAhbZqQcFFI+uG3peN07
QaAZHaW21klv/D6CBooIJp6zidMqPAl98f1WhR4iMKua1LhyizLj6SmYrVcW5J0L9stz6I5Hiq+Z
A6koki2gfmwm1aTVR2SAiQlg4aE3cxHEmxNcws4WRX50kCMGObMY66BSal+IzCIKGdYTry208Hbk
XccQAlMZo/qWEkVz31MuXMEw62uMgm/5JkAuVpNa0M/0OXPiCqCDDRGKGShSzxcE+f37xNj16ukE
WPw+081R3xCqTeimqyPG2L+OS53WyTJXRYftkkULa4uov7sdeDGNeodizISajBRA8KYjUwLrYR4x
xI3DwNOO9imzEQ6La5JPvoVmlM1ohkqEA1ksWCl3ovUr3FgIfcqPn38Y3FMfYKNW49TlBKevF5cN
v6ZVys8yafSfw10VovKhxyDKc4s2hWCO7AkTZ1obxVLJeU2PjrSekIVEgU6R1m5tGv2qdQvtE4IV
7bR2SfHz1wKnYIVR9yam7B2gPXy/7dah9j8Ggubxkl5qAHkmQtG5W3pC03ZF6UgLtdJ3MMU0xx08
EzRhfKEsHNh5TTdva1o5gOBu68BnhZoY8GCVGxrpHn3azj0qGy6b4jw32GutQKQ07SyN9LxR5Wls
we/J/4V4ue0trOLlwMupuEppzlSxM8tJz7mZ8nGUJO7gYnWjFNxG419RTu53vHtfDsZcNNkOrMVS
muzdZBxIHeWOp1mIpfNJl4C2YcgyrdDWHvbNuo+AFlWCXDS9+o+AP8V5RfSc5gGNA/zUGefdpVzp
0GXG2+0WnRMc/udS2Yy+4Tz2bMLrWqukYU52OkqrML3Jp+0d8cfbd165CyXltQIMp8Ht/4VBdJ+h
1HddwZJoWBCG1sMEutOHavvuz3YCm+xMeEgqCSFE5biFc0uVOVHGk9UVaoqF7QOP9KMWFBE8/4h0
La0zaY3HudkyoVPcfiyWvIx/1/sevNUqdY6602U4qfS9jmzbDhDw4C/fuHl9jSzK4MJdA3ZpQ8kX
rhcbYaSWdieWKnneHIqD9vmuY2+8jx2tAsVtFPrccizN7sprKp6jg9SpsXR3Q4EcDI0I1yzCiYOl
Uuccf4MAvt02hrFqL108heuz7bd7siSeMW1FrSigttuw1tY+dvSIIs28U+Y7qPjz4zf+dQXHnVi6
5kD3X2W1fUbXYnZ7/1FYKRhHj3T7w8/taar7sX1d4uUcETVwyR6Ek/dEkjxqOgG834qzLarrt6o5
Jrn28z+LEq0JQEAj7VH6bB9eAOCmuYPKljA3ySaZWlFa6IT1P1otnOXHUoEV0HEqlNPFof9glc+F
Ji8sqF+90nJCn/oa+kCt1BYmwRZi30L9gHlO8fbetywIzOAgKmdYW8VnPtBieeJ3TywvX7Pr8X3u
Cil7mRXw0GXBTy6nMW0csPE1/HzzRHn0lndRKl2TYnaQfM0lVturBJ5aKY0AzsYj/IyvuFmXOnpq
zGIfMakE0W4yvGkF7WvBQvwTWLPsq2Rh/haWEtQYxzwUveM7voQwY462yNXn31Lba2s5dl59txuj
MimOFKrOuyuAXXv9pl9i88oEA8l3/aOrnKhIfNIYTMOxpzjSOYfDfM/pDHTWb1S8O8RZRQ83u+nG
sGu2fN5iOI1JtFgqz1ZBPP/899UdVXO+xqWIcjDkI/bVWfQArgEP4Awp3PU36APa+Eanm4/UuI6Z
h+GqHNISNQlb/xEn9hiIkANJDeSIg4HECuL5Mcq/0YgZCUnyp9RRRrVo2v5NnoMZUwuTx0x/BtSH
mRp6/S4b1qxrA0wjQfO66EreXZhc4wu7YzT1QXbrNttkoimEM25K5F6kd6M0MGNDVOxcsdWENtX2
LUBni1tO4KL4DepuxW9Dr/MqF/JHfqhq0Zfjz6COrGSSsjeChLuXZPlaukcTa6Os5haD61ZzvjCc
pyvEsLlljniHjRNJd10n3f5PtkRaDA92ytFV7me5TYX+aj4dHCcjC9pGV9Ue4n+iqhPrXK9v0Plx
mIzThbGb/RlvC7rIkf7LlWYdbAoheQwjyXxOeljLUnE8+Lk4lU2yspp2+FCIRmXxbTo45HZ92siM
PXTh9BHobT9qWuOgiKNoZ0vOrPGDh2MkBCwr1t6EGBBnS8CLjVoHw3OEAm9zC2ApgPaLoICeh8Kl
OaHGILsyQhDDlwRZdp8Z00MIXjFPBguRRfb7AE1jTU0YPpkYjhoVx1zIdxy+eTwW6OpaTJh0Dckc
EbCkvDkXVB8WCUpJknDSD+tuCYfm3k6I0IQyEUBlzFPe47OfRPNlnt6RevIwAZEnQcjYH7yRaozU
WSm+aeyGqt6kyFgadRP7PDOd2ZzHpZFmEJI9aXAQPeY+LN3/nY48caMKP/kdVy3xS9xfkullQOOV
GoTMnuDM9O+jXsk2A/+BuLUEayHnI6bXCvjNo4PCXzRtiTv507V53g0ZbozUVVIMCs2NoiuEgrXh
ppaFcszJnZxE88Tx4Mw4C8d3v3jhWiFSWrYj5fm/KAljTuPW1QNNaMK8m7TrWP4YP2LPquhQ0jia
fuGQN3GLQPyypvUwyC1XJMIy0mboIgomLuTE75Ifkomf6/9zV85Jcf3F3fs8pVLDfgAeWUQOOi/3
4T44lVXgFdw18I3rd+qHuZDMcT8KO/gHC6EBzzPkjpG/lpkMFbNUHErMxeIOd2qNr4FzeNPBtYNX
2Ne/ttWg/2BScnhpW1T6j/ZwguQQOMfraWwHOM+uk3Vh+HL1Ht8Nsp8cVLAL7wU3i1Rx0DNZFYUy
nTzqzJ6FfNHxp6vHcuu6I8DXwaWy541L/ZcyBFvQEggNsM3RqwfpqKEhf3SHkvn+BQaQp1j+9mWI
3DRBhq2t28b0ITxwvt0Q5FqqgwImn17emw0EA1luiQE+op5ASAgHC2DEbGiAXRYCMFgD7MQKEnEW
HKuZmGStTMLm3zoftapXP/gfk7gVGM3Rr0npvyhXNP1iaPu7Qu8JTfKWgeroruglcrd3HZYzMU84
zKt7k6gGYEzLDls4XXBOHkPZzCuDE8xpe1PTv2P333ASzjeDOy6cJRYXKwjkP3LpezbNUQdPWyMo
F9VtWbV+MEUcIujEOJEBiQI+nI7EpA2Ds4t5zNlLw8gv2DsknyBQG3307o4auBTPB3hCZ7sawfYH
VmGKOo4x9mkV8OAmHE6nSV2R1pImmBcoatcusBNuEgKMYgS7Y/kf5V++i2RDhDWVYWbTYDUOIjuQ
JotJUAJkcVMRKC1h6kjruIPxvuGpy4hy8OYpMKeQMqbOUwGWfskthtcduuUStAwqngM8khsBLuwt
ajLU4a/k/mg5QZyD3X7kNED7LtsH3EZINpLbnjj/wr1C/vexyMLgR4OgA82zqtg/TQfxBxJ1WflT
4s2thQDI+51rnNi2KFe6E4xvimKdsn3nYAM7I6QAjh1WYKb+CRJjbVDNShcMhHu6PeBY8cNFsGM0
GuCkk9PsLmKfHYKvOwCoMNGhK+k6QAK3wnKhTfszkxh/2WR1oq5CehM2PiHM9N7LF0+tcZ2CLMou
EZUYb6T2SP4dsQBXiZieavYMgE97vCB7b8FCXMZ41dMEPDNJpzt4HU7cexgsdUtsrQOgGsvIwGN8
ZXg3IGJnoyBeYlD56c18kbpaT7ISHM9hfUfTGyv9Vioje/tS0+DKK9X+Rd2QqPh/AWmeERe2BnDm
K6/oZDLf/cGKfHV7+tSN8LxIgmnaQ2mCNFXRv+qhr+YcefDvDZcfzubyO6kWfNzgkSp0HBSAQTAT
r6W/DCgZvbsdKiVBRAZOkwsyGTzu7npPEly6rqj5jUQ1svt7zucbQMPlno/gHCyBgu8CpYf/70U/
/qHGrX7QtrHuIrPHVsbVMsMJbYfGWIs7PMDrK4JUeW1LkmPxoPSscGC8MDVzVD1N/GknbeOv95Xs
QGVpm9RrufIT+YmwR8+qOJcciPOlY689Kn9Tt1GpLwm64gNLBiriKV2Hx7rcRF3X/N4Fz19AngCO
C19QvJGrVyH7AMu7gGkbTXnSmNmBWOLfNFopW6maAxw4acK0N3OOnoQykbfNmr7fiZD6AyyJctZu
H75wPJLCLPUHdG9lif5PKVQTyHp6zfQrYsRwNROTxScNSstgf4M2YO0RMVRJIiiErf/D+IIF96sS
ALHnlb4s15krvLf4ad0U4xyjKrnbjzcnAhppsmKaOErRG4/bRPjxXYrkYIhVrzpWiPndN3lQnnXX
SAGmwjj79NA1WGhHX60Qvy1aezUiKk+4VEarWve4PcjxwuphwDRXDCl32vsGL1Jc6EUKh4QcJQrw
3DvsPC+eBBem71hZxKQgUlV0WJ/TbUXfN+I0M7AF5O7ChIFVWjkcSC48j71qCuo0vaCjWDouInYR
QQ6IDwX2SjyWB0Ds4aQoupSdIhIvdhMv3sfrRA2BICIBOV/kAIrgGlnsmudR8q9uYttQN0gw7Wn1
BdF57AcnA90E3Xyy1cq6m+z5nTYnWr3L/f2DODKvYg5MdAk2aObqcI1OhCV74YTZKkCPnPvpnoYM
th0V99o0Bop+H3Kd4DH4ucORSIvmC3sJbNmIJAYsOewlnTZ4CNTHwwADu76Ley5yG2sAzdQXZovJ
aFKAoqREEjwoUUs/2N6+qXIuNjQNI1tOwcOw3w1BI2x/226k5kNYO6kDSMSiuSNaVx85ky5ejA8M
5rcgSpaO8PLzlIXxCWd++B1DkJHteozYOkHitUCMTKyvWgYN79OT/44+J8u2rL4nDlaMTa4hmoV6
gTWQxNH9Mp5Od04sMYbBFqgzrH0zX3BJwy1/CsZ+UO+gCOBxs9DtkSYYH4AViZ/PjjeS3nLv8lKL
kSOqAqao/OIAwUn0mDZinoKwylveofQJrH5FT0xlISEu/y7Jmb/MZo9NCXchIc4J0Xj/fRGDai9y
HohqcjrQb4r3XO0s+rIcupBHIJu17vuxjVej08hrjSgWi6EGZorEuZxjcU8MXgDC2G+ONVpqFApC
Ah7NJCibhS+vQLWujzAdCpTcxxebzIPsfNQNw/Ug0g8YEC5n2Etg+gbyaLxcY4yx/VsV93GKIUQd
+uh69b0VDuvZJQKNuMtm+w4m/jpBLEA6aakp0Idbg6cEZwmQqnG/nJd260r9wcXz/OK7S/4MXAmb
k5CoyxXR/1AOwHpLQ0xUjf9cNYtfZp/s4CnCMNjZTgZVWpPZnKwHRBt2W0LbsyKjhSMFalFEqYSM
ld0ZkQ2qzpwbKITEKFtiwv8vcSvpXh3ZL/Rzwai+8cs0lJVVP8xksLQrHIt1zP0F3WxmjaL8p19I
wiJI+vo1/XYzJlpaacuIsgAGQ4xT0Nb3KF/ZTVY4ucIY0w/g7Ltl7gHUbsWWZr32Zibn4DmHs94P
ewPfaNCIM2//6N3Qk+8xR8sY8fvgFv4GlXza2LkQX8IVZrIlCPELUWKs2buAlTHHWpEPl5y7aQPR
PiOkn2Pjl9941kBXJqi6tPdiTlfT/bviW31DYXkpwVS6Sr4rFuUMypZJOvH9PeMUvPw+fWX9yOoa
DY6zxVQ1umV7Ka23H8krYRQpduhrkQPJqu7t7Cko1EPj2C4YUVMGYq53GP1rYKv1+7/Dy7GVRb2K
7iU3iQMUdre1DOqcRzeq9qF6yFLS1f/oht/l7267eFl3Dx7L/XDd0hIQ3kClDquT5tLHXKtMgCWA
QnItLNQBTEEC06WltOdQb/hQrQ3CVd/IRpkgovXD2Mveb572q5+wuanXm84qnFBwhoXahZxJtPfm
0EDgJmB1TaBx+ZDucP7EC0rVxbKzZL3mPsdp/Xnd0jDUosJKBH075BtQjee0oX1yIcb1gOEwSQY7
+R/5kr1rjJ/Kqfzmqip3NhJpv0esatP+tb8WVYGAzWI2o99F1fqYse8RhyxH/x80Kv2X9KO/loaB
4eTx1sD3uXR/kWAgUoVDVvInnBe6cfYCF9DqHa7tKj+ZItsQIbFfweGSi5j37pAFCuChyb2exyL1
46v6x71VXVS64gATmQSSSXzPoJJ1xDmLHeAvDB+s23KVpK05a5+6Z4rA6GvFVQznijKx/V00YpZd
XBQXnGTFErZGXRkEYgP3DL41Sm6H0XNF9hVVGJBZbkKCVxCQXx2MLnkT7Fsuguiim2bIe/UAiC71
kZl34gse4jipdHiZQ82v7VP41vgdDdzjMvITpZLr9LSzineEIXYlwEbkZtrlyTxDFP1DpLeZG9Qb
yUQ9clhE5b0yjoL9K2ypdb2KmqgG48jz+lvECCBeuBh77b0MqgszMiLy30aSxcijmpvR7qcr7DBG
oFvUXeAEaZu7fz+jAFWlwGpY5G91CgMb5JtqR280iUddK/T25h77/QJj1Je92xBOAnWLdZwzC5zT
JZCjHM+sDjsScpcYdoqeXbZ88Gq1D+jKL4+4TAFkN+sgJxI+tW6KqGTlAZ91isqxKRarL2BCY5VJ
vNuWJi1qCN3yvDlBC5Lv6ab5R+C8Ty9HAtQBb82WJQmbbulGa0VNUycd6rtXK6V4PtKzzlWsQf62
FVEhynUhqUCddvxJaoztgfYFe1b6KevDvyl5HynJIwm4BB+5e9zJH7i1jvM5FQS2ZDfLVp2q19Bz
cT0bZ9XeDRVOD+SCGqnh+98WKCCW9M6vHtK5egHrhNfgKpKCueNvdjhRyvytAVvrNTpymvQSn4PI
4k3NoFRdSYvRGgQEmUgLqSwqto8vp1fdCuep7dfPF3tQk6hzjw8oIyzMa7FGhOiVpNsZUEABmxCA
bLpfzZNqsZQaBlYIxQ9mrX8ahQ6kNYwVSLuT0CD/VVeXhKmRPApkW1ZKL0RIwqOZ8ukFTapBEdRB
QRlVH/l3/W/X4BfBkyROrRjHN5sacIA1QHe03kclVa1/PqahsoDUstyIPQgkxJ25pa9i8di6kR3r
s5O5N7IVmuaiViv6G71ZCXiZnPk6K6ymzx3F3kB3e31mHnINixlfDuMR2zBQ3PQzwG1LjRhNtfGS
Ije3YDONBh+Rn9e6nEfk+yaIFUCS9h7c3I6F4y/P5nA9oGat2Gyb7Ltg/x7NEo24db5E0iNC3Q19
VYYmseRWOATXe4qSvaBs+GCOmhF/osVwf5Kgzit8F6e5M02qj2KbIOPvaZEYNXKX46HcE/zRAdvp
my30rzsbVhdVaqrv9wq8g9cPRAwmxtXykuDWG2YAj4YedAh1wcdt4HrxodWwtZLuiSw0IBDKxxJE
9FpKhUJlad9TI4yo40HDyxzFaSmvw+2Wz+6ulovkBLtjREvIhR1zA7jcMMQusXQrYvkUfeJVp8m4
eIQUUM4Ci7kgfVPnuzhaWZCCbv8rieEQK/KD5Lq0+CiLUP3v98T5vTl1MVj/v5Vu5hqBjr8xHq3A
P0pcGHEPtiyVNO8sqU0SVvh36U5L3LzDiw8SKLUzfJtNBjPmF8nInuBbz7c6T7gBtT5G1VGCiEpJ
dJkVE1hygq2Kl4R5QkbsJaE8NH1wBHgAKzkI33mBJ0117hmdex/nGXvqMoJuKMlUHx8/eeOrlFIZ
iA0IEEBd4lRqSwhN+nHIbXwVvQJH+hVBuOADs9UpeHx17TVYYN1ySDjwfgBxOjTCOpbkm1F2k1d+
y2fKMtXjlmG5aaIanxo+sz8pn6j5po8Didco/PMik8u6bUj55lJc8JwbwQY3GvZoLXDjeBlfktv0
RPJX0NoWTydRYQEGQM6TYq+4NwLBGLSVcNdC5C4Io76L3d9mbyMmrTKHyA3yKAdov6maTzeZDV05
KzQTVMt9ac25LU0uLe4zbVK6N7M2zbgdKrn3CYeE0zSEVqva3ITV9Pr+aKAmDi9FACf5t7VRUg3V
opAS2YOOeFmrT86SL94HHCqnEYex9GNgEzrCKp6pdSGb28SSSHjHu0TXF0bMF4LoHwfdik1wRPUz
Ek4VjG+tL/7KdpfopMC3eZX5zz9ZjJ6Ji6Zm7f6wf/iu2eTo77qVg13LWEz4CGKAMSrUk5VVQGXu
05Dh7wrVjt9VM5oybkJ5N1pnuALZG28EnbUNIOMLNo/96cQ8e5zswA/VH0L20Dq2YHlDmCx9lKje
wPSIiLeGhuOsGOa1sIWgtJhtiDXjoId7l5Abksi9LSZR8ljGZoHwz97U8dWIaBnEIEEK7wO8qzti
SKQUpfcHetwHmXk38kjSPPYrkwCvy9lWYU/LsfjdmaGr3P/vubJanKL4fQQ9SjRiSzjRZ66TenG1
AY9fhjjpM5tTlAP11pwNbLrVJNg5CE9GSc0icxh2E6SGS9w1psrS85y43HZ+Eo4ipUdpQGl4ZydW
+2F4lLbhx9T/PxPjoCysqhXG+K8SGRELNmYsTcOGPQofEoQ80sWhSfBZDYGFc6ZeaZrUVPyXf7eI
4EwnE55ycQP1YGYJ65qSvkL9UKzN9wLCoNpf242K6yWvRZTWp/wCSRozVHxyPcLDF3UFuHMioyRA
TTpyyQ2AKliiOkkxdfwgoo0y9ta6jY36ShLA+Ti0r1+uF5hZ9jLw0MvouqvtNvdajoGGoLmbEsJg
MpP9QTr4rOYtY9ac2J5M6+s0RNuTODhLI6GWllGYMfYRfkAtZiE0CLz2j375OFf9c5mqRrGoGK1R
fARnNSKHxvudWU8aD/zPZTfr8kYX3w5LHQmLc6rvklA/8KSeFzM4OSOFh3RLHkbA+tex97vgsCKU
fihln9DxtBqTx2051NJOAsUEvA2FteQj4yq/E6apteJJTr3SnStaCKKV1QczJ6v2hjUVDhydSEtB
uNNJUzN7QIVlVfGqW8JxhBV1yfXOrAV/OMUrmD5uw+h5XAtPb/5ZJTwIWqjI1YtTLKIdxV103v3Z
xd0XmhR3KKfbE8jnzJKrspgkEOh/hXqyrvWPMljqqe6cPSgiLY13ZnxlepW4Axy796vCL3FBtwA5
46kNOSoBOnKeeWYhm+Fg2CwXxBu3sfLLG1buyG5OFrs73s6P5if1swc5S17G/popbsup1Olr7y3x
axUDsf6gaW55Cg6DMY5ffKjf5cp2kAWEebLpyFMvso01HdQWJSg5hcDkcD8G8tcH447nv3JRRXn2
VtEetHBaEUk0teoNnXKgRTHOScWN2xehu2fP6W7GbA72+cDMyEWjYz72mxm/XHl/cq6ENS5PPvLw
1rJoeUhMD3OZ2VLKErrhm0EwGeVO5gD38UbUbljAyYqR992OJN15XsWeo3CCoJyEiTvR+pnLa5jk
DD1h4yH3Oxab4Hz864836xflQCok9nFKO3jwcSgokWWhFHnibG8PytPLDRMcgrFl++Voa3vtPpv5
ob3Nwuzf8tRIFOVrSyli1SNaijczUSENVw6JlwgYAlRzlRTHwWL5UFu4DDSviudPPMngfiPFnYl0
X3rkp76TwUXf4YzlNkNytA4vaAlIHBVsueq4hzyONwbA9y9OCMdJgR/HpZbZ9NUhZPwECksMkFm1
OqcZoSN9X64uU2Tgu+TV517nIxcWN7l6UJgHwIW1TavtWQCN9FaxUK00rREuj74ozK3PPskCjSgK
rY4VXQVc3xJNzrMmUVEciP8E1ceUlugwB/EFuzMcuL1OpJ7Js0R2nJ5iMZiDQ0M/adzNnXHRYaOq
rt8+Ad4K9Doz2JQYFf5qKxCGJubm/T9qF9+fREsHJ2pWxMrF5nY7yliU/uqZ9ZZFBCBI4DMmRfRc
uzCsPKO9uUKhsJ6ZPUEhhPpJSqVPwOEGcObFBkPzDeVjfDBJu7Pr8wygLJIzwYdEljX/xks8Cjl+
/wjS3LyWWGTMFqEwLKX1mPxYtfWpxmsVdjP+lIOhGE5q0pp2MekKlK1JW0XMrmHVs8tj52UFKOe1
j8HitVjZgCGcxyFn2TMJ1ppGIFZSQn+7zQenXqzj2A7FF46+VpBFoJ8ib4ADpZ2QzM84P3VjbYMw
m3pFeb6zuDyPbb+V6yXCAIdSfXZn87ebT07fJeLdBTlTsCLRKlIiYb0fcKGBBREn3ik44yJbKuRu
Be0O1JnVGIeLzTJQnW/YJHl9POYVPxuAz/1KF+4lbOgBJie3zw7L/nCLVzr/sIdTMNHuaUEPxhfN
uGgmayslZuKe5rm/LsyLtXl2p1g9MC3T4WtsD/QP1jzbuR2dfTv1zr9ETUHvmM3JlrmP4fSelLya
6fmmWLyky2vCijIfWkTG7tVTOBJVQaFJaSrSwmy9jg8p991p3e/bUTv2oPWu7Gm1Ej2ICNSqhkJG
bAcdD3C+hBQFnVoTGEq3aP8Id/b82krhXNi8jeOeG97fQFPyDEDv0BEwwcj2eeGP4kIAbj3h1afQ
oty/n6RY1/vzIDhgUo8K8WASrQT4xYFPmKxyc4gyDJ04PDKo3iU8PLmMv2HijaL2VjdYJ6dU1ued
c/xDW+jDFEpIA4MnPMdPWnGY+DcBmRir3zesiU95wSSbD3rmUTkSfQwYNqxpetfxoBcdtdByhI7g
n2hGeodASPvI+MIoaU4sV1AMxJUVCY/yA6xcOkeGIFkSijJW2DQaBtSgo50LMqnwNQktV2Icnvzo
ZqsURC2hDf07djtbsvZpcDPd/a60feu9hTgRR33iedfZQA8lCPXpgZsLMcc350xRvyTeuIspybE8
gvjcFaGKU/jh41dVIvcCniqpK27yApIxRIXbAnSI/mhPMacWmce4S8f8xxH3PeHg0HzS/4mz6N6P
RCwNLVIc+08lhn0JtKHIfQjpXmkOfG5mXVWYbvW06jUX4RZgxX6g+qZ1ALlejLgA4P/uyoejTTWb
ZDhy++gtxvqJpT6x8J98hecgpw0Xzz7ZegZc3sUxs7ailozFURjOxeGZeFqzajB/SHf/8Y5miHYa
6KWuKvXLs36S2xeq1q9E6TTewmLa1HQpGR/p5mJcezzti/lkugp7WQG31L7EM/kf1IkU0OIaichx
+SQGnglXzjfu57mN+WyubHQhLTlaMi5TAR/bvwN9Lh06XUzQkPZIjwpTkZAuyywU6J762dh5jMnU
4d5qXOulU21NGtRyOV0w4sNxjKLKlLu61IpcoZ+Sya2AtC+DRdjlhNnmQWjqnDQxEpwCzelY+1RQ
PFex1icNCsymMSK+Iq7PsogF/TPsDW/nhmlFR4xmHZTwOOJtJHSAyfe+H1/oMYkZDLS54JSMYnfg
HOQIwJvOfkrYG6xsODAy+1oQkk+O9x7q5LH3lJ+3DNjALP3Ee/wjnrzA0ZoRd+4Xqjckiy0w50nZ
1XFX4PZurskVYyLJNaqC6JZgRfSddXZ7wjTQbbJN8+mSitpqKKSob5GAma2KdmjVzyD+mcp9yuoT
kcB5WEXeDvQ19OJGoTqNtyvr38RXKFiBCubmrgnrUzz2MTCLNKA6uDgS+FQN/7xo6JcbkPbzDe3p
0C3oF7eMCzrw9tHRm7a2t1Pw5URZ+Lmj5N10AdvERzRrjo1wMsKtjmYPL0yWCP5NvKO0HASRM/cT
Bpv6k10kmDq51vqzMiELIXdLacLQt0+2Jnaz+5TKVkBo8QWZryiupjjN24ZO7SP4TmQlsYeXSHP7
otAsAIWERwJ3d4X+VSNahj7KNQ9MsXE79/udOq9xV3HuXpxOMOZZ/m+YbCFOXElXuqrltqly1N/M
RpLj1nYm71qqmgMKMYxbM95M0pUPr03HY3dwfEhJzzu1Q1sNuzHqPK9ATyZKBsvMnVt4/Rfl/RkR
1/h6O4lPWpX3jd/Ux1VPGlVBf8QZ3s0IP5S7RSVyFmNyrNLMPv6jgqopAwv27ciWX3uyekr85MQB
Kua+DA2N0IJK37XwB9Y/RYABUvQbakImbFhZNhJroBwUG8hQ82h6/vqa6W/+g1Pu+C3vfVup7U4m
HMcJrCj/Iv0JtPkhg797747hM45qZMuv6dHoTjfb88WrQLoWKlpe3g557M4CHIWA/+klIfDPsiT6
ECtvxcTDn0+pWepznW8IZXowr/WVZAJtQd3NDxrG9H2Z8I/+0UvqrDw4xWpOrT/XyzL7CKYMlY82
vjECuRtx+Jmv0pypwqOzZIlr8z+1SWCktsD03GFxDzCjfRJKxW70//WwbCtbkrkIkkUDfe/lNHUg
P4jCLNEp2otP7/rRU7NTST912zi0jaMTI8r9DTIQ72TurSN4TAEYHy0FPcKPUvn3P102wiexKUoD
O5l+HDipuUv5gvmw7SqYlbMfZt8TSnT12stzhZAnR/kPzH2ndeex3iFKRqzchCGta8PQciJCW8vQ
8AdmvPJZF7+8jSjxodMgwwYuccolWjcmv7aJh/zbLxz8EAp0Wc6SW3YsnQ0SALxlpmKHdLZSVMVV
764l9qCtDfm2TeN3FUFw+9gz8ofRwSbYqX2VgFvgggVUhJYar9g1ziXy9mRe6I6yLuYYrZ4ZGhEq
Z0l2ynhP5a3EHqOWalR+j2vcgXET2SMB/l2KzPUqsV4iWZX3Pb5uBb6kL9sZzUD0GBtw7ABW7YC4
mVo3ligTlbuzTCpAILqQ10kMKv1fvcFtw2qYvM5EYOTquIizWSfq9addT5ukiM1JfFJvVIEvr1+/
XNZTmTjuLISOB01Cc0jsywphoD2LCvZz97Rjf755MJtxDx9ueCMTFw18gBlOnpFVy6GEMlpmXsJn
MD1F6g+tyicEPJjUdzlmLK6pwf8ASYv6f2MFFKE6Wg/HLBbUD/J59b4MA9ERlbwkb1bb5OrErORD
SXlICgdaRZt9ozqyDnz6Hma7AqA9TEzsEdCh9BdRpTT92bxYXsOYzui72R8h3+QfolWZCBTKCib2
lUeGFM2M8W/C1AHX8EUMjm1Id86605+bQu2ORGm8N9NtI0fZNXb17TKh9RVCvnjQOETYeyyEYuyQ
r51SwQJzbhRQrq3eZKhfHCDIPN3Z2IlLxs2Idwp4gtjR05+9tFWaPjV6nVtmqq9cV6PJVGO1j8gE
77cXCKxVGXHwi9J/aum10adEccdvc7W0NNHCM1/AgDMZNyLSy35PL15dRyFBbHAI97/iIJHMtgJ9
/dNFUKh+b+29AddtqtSjv9cjm3i1lh9i1Xy1PE21DXoorg2zFWsszco7IR4lM9fzlC93zyALbsap
EBNzh6flUKOhdmhlhC0snslShXcQ2XRWMsHgZQ2CiK0Yyc8UQ+LM3TGlvwF5+9RePvdsFsyeMc1f
cDfqWhWHpe2ic5GXlkP9gcoutuYCWjElmG+zhPh8W9e3MiSRkj75EBX5QJ10cd1mBFhHuEmcUCvd
x1eykSpjlp4NxI+4HeGZ6ZoztYwNas2PqFGCmcW3H9BMKA87mZFKBrFc2K3fAa5UZNxD/hByQQBu
026jmFcWd7A5Fj+TnIwA0uVUxlWo+cFN0qeV0kJ1KtfYEUTy5+s7qDz+8GGNDKFc9OZD1qp/vqmg
sUj68mCwJYQ+vajemnBKSKmZ/BHhwgamTZOzhTp0H35khazvJvnD5b4rgzNWOfE/HEYLwvDqCEQo
M5ByqbiBJIT2XcIY4dW+u3UoT2NcI2Dyp+FZdV1aK7Oxm/TgD+dvD3vi5lv2zatVLp7SSor11dA3
bmiX79yP9/Sx/RsUZU4Avlb3VMcB2sxjgq04arRlxxOPzQvaBPMEYA+8U2il+Y3Gfcqz51YrsPKT
SH8rKuQKdxZtW7fLgc3RzXQCC0H89EMB+PPEa7aToVEAWv6m34Cc+xMIRK7faQ+cXur+3B0xkc0l
y2dKSGh2z8gwd7BDEKwP3GHIlMsQeVbF5mqAb9fYK0gG3UiAC2//Rwfb0agjT9AoAkq5O67U0f5h
hA+e1WqS7IGdmx7cqyBDwjg1zJMtTvXFFzM+PYIhBcVUIJULzG/ZqDJjJ6k/RbBPYNYatx93ZDZa
rBOwlp5zw2hJChjcRDDPqC22JMyzbCuu2tZXGKSsgB/aftH5oK1D3h2QxKyZofqVPy+fX+6+YMXm
hrI/yiPn43wEVNVKaIsenDrkxR07pvWOshcdcDhwO3IGr38j1aFCDIe1svr0W2OYi6pv2OO978GB
Np7a1dTeRXiUwOWLwJTY7PHU013IsBuLAkCy42IzBF22IqnxCklzkjRgqLlRMBvhWWCKu3KNtQjz
Yngb3yOLKQmJVKCvCgabsaVmW4Kh+FW8E7D4tKS8+Ox44nmBNBUHyBp2bvHnu21GgCCzk9s/rNNM
Mszbgn55RlHsXBZgrYhYLLNDCA4MTvMKU6eWWWzGhH8LXRsncHq1n8WSjT1xnr8/Rtp8cFGaYk1f
NqB6neEoAIT5OMN0oy7C1/4kLKS4egLTendlo9JdUorQOu6v7Je8w2ElD9a11u8T91o1iEJbaPh0
/+cmAG9YsjTdUoirYIkNev0gZ60GzokyUQhdB2wHxBHjTay/+eDzyJ4Kc+C7D5m9/etakO0StKRs
h3OQGdz+yQodRhPpCIhW1/si43XgA2LKCu37TavCWy4OkpIpzKIMt/SN9bV/gOAZ/pcdVXvIq6GV
OI5umzUj28/PUEa9zlQ2uuP+JheiM6JdUNEK0jc0tHzHayZ5Nq8VpBjh0bLtoVt6Z5z+PCgscxUt
YwfzZOD8B59dE2thCSsVH07x4dZjhR+G1yBTugLFLtTXTpBlg/QukvxDr80RtbhdFc2E+ry7/ZTo
TsvOTNuZ4L2UicAA6Lb49XSCHLCj3EyAHNgWeD2Ytbye8adU5U/8IXGUPr39OGzhAF6ksWbQps3e
+kwTBtJSGyYVXXqD96exnGYP//8xRdwcjrWxXJQSibLX5Z/3baUT19BQYV9O9PCq31b7gV+7dS7V
fU1h7a0eog5pGo7PCwIhIMDQdW5H7e3JSRns/vUKyJfyipdl4/VhTthbNcqs7PrmBgipVBTDoT92
naTKRBXvbjj08uAEMu+cuSEA3rbs3OFQi1rkzM6cj7ci1Jp+GSUUphqm3NtcXwzrDozM6Z/Ubrqk
IR4KCpVteabWENNNujTEHti3f46DkuptGp75+6TTL0lvWVNwuglok5ixO8uNOc/daxx0hap8lGhb
bbZZIqR12GWnBoBXDsogQK7tTkWxTv90cY2hr6whl6WWKvYsOOcGPZPw66lSaMWsUVMWuooNS41l
MRQCnNQEEvL7dFnsEJ6DzVMxoctVJ/5T8TCPGljZ/9qluNDBPZM/uKhzQQBJvyolkPBF9kB2UZTr
/G+hNlpJqw6oaJ6gB/DL0C3kYUsdbDrPNXmmyx5s0jcBxBNvAvY2YWJKfMSTPb/E4tl4wpPj85pO
NcLUqRNXJQ7qEqm32U63DRKz9YCwrki0wCm4BOn8gx0bfjeKlAEjenXKq55Vw4dVt0oU8IJy8W/T
fzw83ssUyM0CW88KdwmredQxEOFhmh+IgbN76a3TK5JhQuY3mWleQnRcSnQodQN0eVkJAnTLTBmO
j8w15ZVIoU9mcvY613cWoMGaywckndtkkFYWnETOFbOyONk25xpoudNjcum6EjUrfmCcdhlUTI0K
kUCXCgqM8UZNHZxV6qTl9uQTdQARPEzPtqZ4qKc4zpICw+CgFQcIG9OcU0yANZVye5v3dqTINhnL
bGwuaPQASMPjFEszBJYcB0li0guCu7aowG0USrcKxVOw2/J7DwLq0guE6Ua68gxpynVYLV27LYo7
Q0WXiLwc6DVNCATovMswbuAq0XnVeeQl2+bA4UbU2krIJYJG/+DZ98Tz9ILB4vmyCT1nNxcQHLXN
1QHMmqTJP4z7OQ+IjgEe5FOu+a0/gGr4BYWQT76lN6ZMe8W+sfqkje0jh782lc2Ps754Q+R5kzsl
AWZOXqBghWeXgYTWwTAVaCBkwcKvlEuGEvS2sMh+OOC28bexbteQ41tq+mDe71bLYwFiykdvZxDQ
gfoXAozA2cWSSZmxaUygQxEAfbnrjf/AMZ4DhFCkOCgg/p1oHwFTloA6dpDq2FT35xrlwYx/lbjL
vQ82MkygUP1r/MjpMVI7FCK5v0yQpmFLr3mL0bakfRkYHsDu7KKN9nPHdo2Mz/i/VUddm+/q0frM
4HHqeazW8L/J0dRq5LMFfmHi5hGZ+2U328jJx6x1sdPAPSyEXLCUj90W/4xoqHccmcEyfHG5sfJu
lGGw8Wr5fyuB+SmAbcH/+AkxRdJ1BPN8OvrgbFjOYmRNI3/o/j2U4GBLAxvroo08M+GmuuVVUsLW
DMFNuUrInp7XlTvBvbmD55Wi6REW2uc8XtfFHTlNSiOangs5zrL80a/Sfm0WIMJbKSq6UykAau3W
T0vcKz9ee67dw20fNOOCIezhwpkR0xzlXpIRD4eAgw7mih2TWP1iVATlMi+/1lTJ/NEgbLxjQez1
iqH5DWqbU3QahNGVevCfLmhMPIdHXGexVMYxikQYx96gCLtGk/0jHI5vVi1CmPXJnLs1tfNHNyUm
yJAAeCqKQQgRiPQAk1GELcY/22p7xQ1gS6z/SHHszgjQYwVLf8IiQL/cFKWt7lsGUkawESi/3YQr
Z09UVB8FcETbhYTB6zNl7XXdmlLxlqJO1VM3TaJYY1ySyzYVdqxxrNueyWyyi7LTRuF83aTiw3qA
7eRRD8LA6R90kdVN/XSHKz2cGSbdO6ekVaM9SiisaOd8JndJI9FV7B2853t3x9yN4uCni2hQ+G0z
XJOyXflPkNGD+fKp2X9Eeh0UAbroXTR89Cd4fZszkjya9fd8Td5qTBt0zSTLr07cgb5i6PmkRcNh
qlmBTcuz6KlyJXs/hnB9MTsE0pHoenfsrWXDA2/SlDaxjB1tT2P85G7m958lSTEB7sxt21wTg4nA
6zRPbGpTI2S93HW6u4HziIZxzNem9R84uT8VjlBLRp9/9hQlMTQhYpFElSpLebpqBm0z2kAUdvWP
pVDI8j9d/gKQiebQsWcz21BTTlR8HGmd+PdVOkPDr66RuA2gohSFbH94PNy+NpmgseZXwImXufVL
M2nZ4AfVFvyRbP6M2R/Rxz0cTOrmSgxaSLghmO0SquJTdigQisNWA+/EgJ3Tn/T+p7HiRsjDhlG4
vm5Qz/VlPbQ2VMVzcmqroVIH9WpCWsGOAfkW1lfn7g1TLOmoeiDjCInRAfb2dBzaDMhhucUnG+v5
i83y6o5kIXvobtiqKowaVsgWTJhOBrKWJaRhOVD8edUq4tox2W6qXZiyrcaNtom8uMo4HO3cJSWT
zqY7mFM5DFNfQsXO5J03lRVR7W/egPHmQYKRkC0dndaewd+dm0xA3DQ4Q7A0MFWW1TBc6TOevnyu
KmJZo+eOSwgWK1KPjKS8DxBhBGY6A0z3Xsx139PpE8el7eLguzw7V196S2X+yRMpCvRgf5CnxalR
7IS3V4EENWcCD5gUwhQwozbYzccuNK63zwLhhngXx/5QuVd+liEkQI1eSZvhpSnFiRrRSD4DStqo
YCkUrL8Unguh6Tz4VNqw9VEhYUcg9oe59mTzuRk7DTHKkP9kFomeUQQhXIxro9wT6qyFjS2eBXTv
YYX7Y9Qsy2ZktHplm3kVfyDhu9d/7KC67F6pfwQisAFmOYldRozSza4nXnx+t5rtO8FGItQEDV33
KBIxxNQ5Oxq46CDk+zDp7nfxhGsO2VU/6OZ12iCHVwiLzng/AlYzX5YFwE12PtK7P4g70zQuMPOY
deLMFHu818EkCffTBfZRUzGNXDWuqR2daUm70PVfFp7R0DBNP9GgI0e0fxVGkK/o6fUHzngtDEAg
aLu3HkXbg4vcZraKj743QMh7tK0x6yJVFq0EnWqTDFYi9OimLbA3gZUj/YQh5PdFu+cjuorb7DSK
Nxau1iV76x0ufw0XWwS9nvl8kz7NScp/vNfdn0pbW7WvRQ2JNmrVGJdTBPBvI96FwfAwHu9mrnVp
9do12ta1jiVe0cjByxd850sEx9tc6h/0EjR2TKmZeZ7sGKOzlbBw7+qCoRqRI45VQsYBcuVHkXj0
OpRDHqQuaHvAjnJhOlmKYz+BTgREpAhMERvby68sc/8smtWGpWuRGglt+2howbGH+AR4ZAT5Jcbg
FG0qmWVJzmcW6iDVqKCPKmXXrgOq5wenUm/yhgK9buKOT3zSLgqtfxPc9ejsHaGFP7QQvPGxRaPG
mmgt5jOUgUNwXXMW56tQb9r1cT6ny/uCtqvvFt2oF3j+zPsrtRbeSDnUfoKJI/MfgZmGizFINP1z
sJApXGEhljCAbhrlLu5TiNfRCXAKL3Jw5dQ7ddtepQewC+lm73AFUkDMbouB+S5ao+fBWBXx/r4D
XrE4tWsIIkeOzFq1PcCKWOJ58pOcFZaLF4sDRsZqDd6zCTELKKn6j0H1J7ptlXViIBTbB2kjLZox
eWu+IcImh3I6K55LwU4pCb+AnYJ7u0JFGVWQVkgL0YOdySw7t0BoF6zgWNWGkSiekeNMscX8Vbw1
zOeCNYFvqQfOUaEoWAq83d9UKdShZaAhCHF189RDO41ZwaEAzfTjOpgrwUTYLUvFD1lCP6ibl5YY
Yf10ojyy/NaHzmhIXhw4uhI6fsEPquM/hRfaZhPKuxB3Ak/MOHpDvpkOirj5Si/Wb7hPZfhDo1hf
4iq1DVqEKy4PPitg3znvVZ8rhdntG+KpZWk/GZ2HR8w5PhJwy8n7f/BNyswV6G/whDR98ryEv+Kn
GFuXDiFrXOejzxS5YvGC8f/UHiB++6DCv8y3z0K7OJyl9AkGTf8EfkHRXdoSfKEckx6Px1xnPf47
gGRjmbxUpZkMnMVkG9e3QvcZk6QR90Ye51/wxKSG0SpN566JcGovLphup0d+G86NpCGen9Fd/9Fg
iwvDQWvktpicjGWc4/jd2a7R87BhpWrL/B/J0gs8xxGy+ihIsxehSxtLsdlSqlHMXCDoN6UDVWbt
aLZYbKOuoKe1r3hRSNVsot4ZV1liHE2Ctq4ddkQDFYq3FrdvEjOtOuYp+YCJVYVdvC4oNsK99KXf
vLU4YOjivawyA4YEizjlG5a5wvnIpKqQCc7nDmK7PeXiL7h9vqD0j8h9+UJaYI9p3IAG4OqjePVF
H6r2XZ/RBJbXNr1TrvuJZ6IIm45u88SdzvP26TVOKzQHD5HL68jxJ7JveQEE2TPcx9/grF/r2y+T
fv4ZAwnLDx3FeCCicCgDtKWzAGq3fKlgCWkZJV5acWn7hiCOLHJh/TEpBEo2RM2EuyloSI6e7Q4T
svxGsf2Pd0FIWv46FFpOw1uErYkxiwTJd/N9UVDr4JcKz3Y6sKKxCXrqwJbZO7ptKqCGVdgsHkMB
vND5IrJ/IoJIqArAHramcbGWLqgXTnekq8mAGbvdfSJMg8Bf755Z8HBPkxgw6vESENXlqkFEB75O
F7KeqU2tTiz5g1Qz3tMbtGegONlA16tU1+8TBz2llyTE060lWFLU5nH3CAq3A0KzTS1b0Pv8UWzO
VQ3SM/hD8rYaW1dcXhkz9ID3sjXL5tVuQVYIJa2IPvJ0UibecHIsArah1BV0fsaU6XjxzZWxS4BD
voIkNlQK7nCbTf2VngrNoiqGuOAFgif3Nv01uqXjK0W4lO2yqc5BikEwRQ7OzLL79pHmz1I9C9bz
WuSQLTnJ08Oi7ZDDYG0HzANbP3nTVrAPb/0UNc0TkkxzBCKn/agcFA6D8Hn5Ot0I64emuBaRI6iS
orXmY09Db+da68aabnYdqTQJ7VD9dAUVPU3YXnQQVzlwmIYflKfc5FpiYwT70v67i4XSl2knZYya
MoHiuUt5bC+CCnpnHiAFiEQqcbJZReexl3WIDPbfzbfuPf7YAvThRIVFErSkcxQDfh2+CxH0/lT4
p9cycrLTrIALktPMO7sF4OGX2Cf1vmROMQZvNeAMN8GSh9ZyaHNJQZo1KGWpKoDzeycF4jrnJMhr
AF186ygjOQpMP37DWbevNenM/Oc4RUU7KY8zT/i7YEzG8T2lofHSqCGri6Gq+oSjr1Xykbfmv1qZ
t35+kFw8ya7YyU3hQ647PQ7d5AR0JIXFsEvkxHjeGC6cVyfhn350FXECqClETNmNL6+kUUo8yWcO
OMOQo9JmFc8R2UU+brdZonp1GH1f3JXcv4Ot3aiIgWmYTQPCki+aX3Q/EM4/4jxYZk21BbnmjwXQ
bUjrCvuljvInPayw6F3B3W8J0tU8rN6hOwxXPkRh95ofukaNLzTT9hA6LQaNp7P3jEe8N/Tez+Sj
hWHu0DbGjb3KCxNFEoceKHRuwgKyPofyG3z/rs4Qtf+c1AnPZxznB/AGEbGPHFPqB2rMp/MjKCSy
udJJNu7yv+aYqyhWzjqKEepud1hIDMBLOZbkwROJQgdYvdHrpw7h2GPBOz8kMfTgdSHyq6dz8wkL
HsSJaU7zxv3pTrIXe7uL+OMuxHm2v6b7YhOCTgbUPpzNidOJfCTnMpQt5Rp25rILy8MGgfbKliVK
PZsMus99KSOrw3EpGn3zZGiAeoAlWE7TZbHpIF4rfkdSm15uR7ewBIhG5eGCx33V7ZRL9IbxsQdp
oYlhbXVpLW5bAv0Lb3cH0v0nKJd6/o31J+PRnL2g5aM6UxZh5poK15Gh2XQsrHswVuYGG8YcsTNv
NRjbm41g8HcInKnoVs+Ye5XzO7aCfU7rYK0XP/S99YF8lSJWyneFam4jhogtYwb8EUdhEDR3V4RQ
Z5BNUJfawDrDLLZTZpax7eIMjui9QOmlztAkb3hnqfhEG0POz6UhsX9yg/7HTa32MxE0tMOye+ro
GtW6NGa1ttpy92LWbgrjWNJRLICvskbxcGqv5CyoQ+yRR128grx4IWin5P7x/P1AmxIdhxbHQh51
0jhroKa8DFf5/UNNwJQ4z2gO2i3FfRXITg09bU0dJebvwPkwdKWoixfKB5T5BNdzcNx6aAsTSk48
Bbmx6Q5CdpaZzxYaXAkoJsgA5LdtzXjgDCR88aMNEXj4Xijp5+0bognuV6zMEjUfuXnAqppKxWJh
w4dEb3cpBKkVYpLmyaEe7hmG4bpTrQVodcW45CccMTVmHlQvBmKBGP63mAAaO3p57XL8sp32kbJQ
/+C5n6CfY/k8nCy3iVqNWKCMY00ulooEGKkG/4rCF7FqA21wpRikrh/GzE8kma7AOx+/RFrIu1hF
d0WI3e6WxY6J2CbxRiS1Ctj3QZihL693p6HXVRBIm3BaAZOWshf0M/XJCtqd9l8k0i0tZluSrrBz
scFKMdLreBYe5aiYZXIJc52TBa3VgdVXqZYtBMq3hJViJznPVM+mnDDWUWr7r44YQC6wkF9ziKhO
yoggHjiN56IilwSuM5XOGkohs+FtFzZ6eky2snZbtI2ruj6CO0II6V/FM30a8Xe3JEHTmxE3Vl4X
JEwKlsF7RMUFJONUPvtTQznxr4w/3l5KYp02iFWtF89iWRpv7/vTN32ubjWDJNKEHXKGysN0HUzY
5X8Pz/KCipqMUmEyS1G3rDL49EtO9lPNOS6mwz+tzHGuH7C53h8heVBLwmGGZcwGLDXvsdEvU2dr
cRTxfekBpmhxRLbR3hGIwlKUxy0ZJKU5H5suVV0kFYX1JUTG3xgo0eO8H1Lp18AC/ecIzfdTK81v
410jv647I8vLja66dDZ9sS/6xtmp3DDcjKlwNOqe7kKUwcfndYKj5XCiqA0hdqe9u12TYjlrtg5v
QiKgtG0aCTFw1oGyoOJQ3Dg2EHCiUSEqyHyjr8dCsHujjbmjrUAvsYI/P6ganUxhe4qbUtTQk2EB
9zAZV++eh2tRYcfVYlB3qEsGyEh2g1j9BYYLRrrRgOgMJZXCkLpPC/bxKR756zP+IocF6ANPY7Z5
onPXLGWieYawvtHXyHFVh7tUvi+8R8Bzn3oyGOkvYGQMv3OEnmyLZh3MYO+jOz+SS+hOvnRACsSZ
5a+t+2czXZJzJFFy9dn6Ua3B5RzZDE/XZvy6aY0QCfYhg1vqMAqmnfCOQ5SUoUEfRL8sGkZerfQM
uwSUwQb6Bfd/MIqLET2zx9d1/iFZ8KwjPQps7AR3n55VyhhXlnW5aWWbFWBc6YdjWldF3RUFR/4u
IhLel33qZho4JIMvbBwFmSGYk4okRhz4hgW/cYJ4KXvUTzHb2Ghc2qS7qMUzJqMJqhOlB2BFD94n
b09ph8mp2OXi0pMQ0+alPlPDbSwjtKXFELuIm97p6fPL/xIdeDuHL+255eKRNk3PijatB2zDCR7/
SiefUfwHEjh1p0X9XSpbL5yyyZFg2UuAFFdBBFYcHztuZaLmjMF+CWTqmd73YRy9dpxB5s0gLd0e
5jtXDVGE/isu3ynljbLkv4xC79HE0rw1huR9J3BHzEQmDVt+rDjefsljTPorVDyyCxti5Y76z5kc
C2LmXA9iJWsvdbYRVqxFK15Pv6FJQK4stXU5HT5wIwAKrObAZAT1xXj54GvQgCiXGGAWlRLHQ6+4
58hDTPPSJu8hIsPjGzk3tNUVYEArVRUDjTflcP3biDtoaVxnGtQEbgYhPwHWuW/oqx7bZdZeYEHD
VMIyyh7wRKCTcSCijYUxyv6Hz/KOT0O0iuAnfjmynqk3DigIo93+l6e/ONewyaGG9DIg0rxN4JUt
DsINps3uHt+JJEkCCpVahvBdw4ky1/zU8PGcCF94v5piTBLUr7YWgii17NqltTCfyIU9tHCMMpRx
sK068SVhUchakoXNAleHQhhqGwGIKF7bz/xd6bG12gBreYwA9qqKrkjSnDlNm7/MyhqDViOSijpA
yQxQRhaZ34cNpbQ5vrXYaABJz5s9dvaNiAVHC6yunEFxeKtUUXOZWWlpyHUg9YTWIYKsiYMhiJNq
HDXoHyVcfYv6UXv/zuPEka7mXgkWRPYZvSDOJsS3N36+VRufDQ1G/9c4/+R5/v1aCXPdzzOFlsL5
VryEPAvVxINir089I85wMtkjVGRtalLODj8vAFni8rfjeu0frU1hxxqy4tVdjLoENTMH5usoLm1o
PJQN1TRQFMfabhF21LmqrNqlhE9Jxonyu8sDiJ9d/eweDAper3KTytHDXrVlG3AfxAC+qkS2yJLD
kq0Q+g0M7na+zkKJRxf+YCN3WqmfRx5m0uthTzc0e2VZPyIF6+IKJnxM9zOP+M02iBddClqEnH4C
aG3/jzf6mGylRSaLliGXa58SBtIb+IVvCRegbMLgn6k5v7AVmz8B80Fcc7k1SxohgnUM5bS/0FbH
LTR8Bcjh7+sfarjVR/7/XZWko5sDW7UM/dp3HmlI9TRiLWhMv4cw3+SBSDBc6wlQ6rsu/+h8qnco
p2e+IXafydzDdmADoMuwLCwNz4cLpGuACxn7uUwNgE4GsVz5Xm4uzz1ik6LTdCaU0MsJEuQwS7ga
JHvuDq7HXPXqLaR4NFfxZUFnm3QtPO1ObDnwFIi4JpsHTJVmmf2UV59/xUmvKn1J6MhvECxHzA4y
ENzZmxZ4/WNaZFM9gqLgfkse3dCL+wOOOznCFzWo9LzNnBEsKmQhB/4sIkW2g4O7LZVeE4FLPAiU
Q5omAtuiTuCybu0xB3B+sTvIjwS7f4/0f7FharOAWSOiuOvJzlfq1iq8Z31NIkMY1KgM8iSRBm86
SHenD3GmtHgGZBQirHkAru0NO0Kb7PDgyq1hsrTnkNLJYA7Tz/J2AHO2nh3DSTtJ4vyldQqgvtKW
WBZI2fWaLG3Q2cw9xb6weC/mnqGU7vqbTb5SPTIltT5Fe+gXd0NYyb4JP/xz+YTmMyTfjDpB9wR8
dZbMQ8DsPL5YtQSqTtqOeqeLJ6ybOz3KOpEvlgQKvJwQTeRcQ7hazeAN2jGTGKs1n/9F8i57JcMs
afhLXMJEcmoK7baGpW1nlrpdrqhzbQZ5HFgLfYDfAMAajrfQ/Fj2wfV4WNjuoiaahuWfz81/FnaZ
qHVE7COkCKyYa51ERhReDuZpw5/SJeNPwMccLa9jnr2/phkXo2CrGqYZQcVT5T5wTdNZK5fuz2Fd
hV1rEhWotsaBODsAxhJaotY8tHYjDTeE9NT1dNYPho68ZfgadFRs94tSVahpa6yAbdUEjTdEu6Eb
Pn1leDw1fdCBZB6rv+N2ik2P5jD8aMc/fLpq1wJnzN4/92OhRMRdIX107fee6Nv0L5tpt2qBlGFt
d84bSegWnKmerwpfoNc/IBI+SJEfsteytPG9XLLHwBKrS3eJ5Ptq4BiyFbj+QRU8vUuR/rdfCLap
7i8Orxxmifs+a2LKDjK4NVX9thsVU80mggXPTtwGtEuF0fNtEyTn1fSFpkwTTr5ge/52PiahVsvC
TC4VpxD9zNUJkw1g8hin38f8AuUSfBO3WMKNXcS6qaSQ4eYg9PrSLxFXvdwuscIFy9k3Aovb6zaG
SAyHLApv12k7fSxw78AunWT2LwHFEInu0SG+vz6XUTLhbfhjd0CG2YWFxjAbyJMf9OJvqCdmEfQv
2Tm3FSEFw7VwBNcd3DGyRPxG5Jv2tb/lqpjzDDUsG7ItTOuod/yCVZXcAqsR5n+Y9BJj9s5EILW1
m2JgqR3P4Ae9PrZR3szOMB0+R8giyuint23F+liKbTOERt9QIFbyeVTv3Uza6+CPzEpRDVU5/PmC
NO2V/T9lweLGmCZKO5ZsLZQKFenlzhXEeI+M8bW8Cpjg824qfsiklx76k+Ai0zNd/c1osQXSonLl
4VDPWcZ88heIelVlhHVvM7gn9u2LGUCNLmOMfjyO66db9CqqtnIpyBkkqHFaZX1NwFKyZbpUeR56
tqynDrCgDrPt+U5wDk91jDFVMR9n4zHP9CuZ1clHzC4PI5WvbIcWGvkMeH4dme+UOq47Er3oP7th
NnTkFnYAt0BMotvtq/xjE0sc2HMgo9ruVPyGwDR2o8m95h9Wm04XKBLuzb/I7XEoDPjZhZkn5UK7
LSs/PPZifYTfQ0mPlVIgq8Jb6XSnigpWCGEvCboqqes2r3GogYgL0NHefIJugl/9+g/I4tQtiDd+
ZiPFy4igIBIh2X6xIMeI4umfrnj2J3E1GJS6B5VqPXtNwT7Crl9YKQa1cjMiiVUZIJQK5/cp9AfS
L+uLRJCt60LeoIvNgIkHFQNEVTGSQ3Syouhioz4pPQBca5McBJqcRETbKXHO/rA+8u2aIYzBX7r8
jweu5RGEAF4s/4ErYmtdF42BL248/X5Jl/QLt+NSYUGrMwde7ZP4BOozTd04h9UGr3HmbyPbNdZA
w311b/VcSP9tJRF8CoUda/fGtZyKtpUptjuZDrTlV3O9T5KijTA79iuK8L1LLCoXauQsBNl6cnuA
echww2ShanYa4Gu0VGULCBrK69NF7tbTO+GFdlljXNtT7oixDIvxj0K1R+2cSN9Mmw0BZRlql2li
9kRh+Qvvfh44KPNlZNg8Y7F7+WVBcZyVw4NL9Py4PRfIniOaHrzyJHKQPoY2PtyJd3GqEUhKxvUk
ttSTDEpmwVepEVBoi8eS+SflJrJ26dbcByZOd1Qg3yb04IcazxvTlJ+rVW39I0DFKStlm2lVErF8
aOhRMYnta6yT0wkF4jm2/9YUPrGBI8ZYMpre0hv+Edisdx5NhcGe+1tCB4qCI6rbnVWvC28W7xE1
YV7q290GH7bJA9UsmQuGNy3ogE+/olfoPylKll4W1G27C4/coRH9HZ73b+C613gETKQ5eqXmpx9y
TPKQCA7Kaozb+FHzV9jG4qv+EXaFoNRlZgafFvhW6kz7XwJAreKYnn75r75EaMpT7y2DnP5Bw4hv
DQnKcv5f/teRdv7TMTg+Q0RR9pgLqB7yJWJanS/pC2AhJLHLU5w2TIAhyUCOFbmqDCPEa/VKIDdS
s5O8vbxLdolEYY9DaulPt3Q5yIzxfHtP/uweaELPwgsrHC/8ut1EnYN3M/PX9DA2h1Uhpugx6SU3
9LCKSO8E43il7Z9/Xm7+xNex99q7enik5tjFB7WLWyDy9WToVmpyt2nQKpMHmw2D9YOf9DG8mh02
5aBxLb/PK7BVIZHrgbPXb/mmjoiaH11eH5N26zjyarYPKf+dmnXL3vymQy5/P2rZ1wQw63I2KNxH
G5eXdKKFQoV51poGQXZNbRaGKCZUBuMsMlkYdp0JkWHZlnJPySjc1VVBi+EXQP9YhekrEs8I4e/p
ihbJBBSA7DnJI8IqCHyIfKbQynVzapBxwox59KExmw42qN8VTWB+Set8YucQj/Q/WZZOvQny5cj6
XSpaeKH/Jjc5vCh9ne9I53QK1z3emrosDIaV3P5Fy7EGXsEhHB2NprZonwpP9KBCUpOncrRJlvDH
kUv2vQw+0YPUcEd6wcEasW4WGZfN+VUPwIa75acEGTQuRDcFthdp+WYGdpbepLQ7AXQ9QQ0S5/Py
wOs34y89UAbfY8Eq4fRPirDk4Wd5CHYQYrIlGk4k2AFMiMAM8Y02kDSfUTfQAKeLj31XwvtoXQN/
xlgjwXTpfdzjMnxX9b2fSSbynJh/Z8llbshUIo/xuThR/XnETqRmqqGj3cfOVef8F3GbSQG4sf6m
1XYM3iX3aLNm+73UpsGZkRN+JKeM+xYh2yxKMAb0pUiz9L/Ss1YOICaGcySqI96z7fxJJ1nPLtKs
ocLLHnPtaKfbTyNoFoMFIu2Lf/oJ6JZA4hNkP9bBmHomlaReVuKKktkmpwgFxa1qAcDNjpTBqgZ8
gdCHpQP3ihTeO7pTZtXtSFjzep5+W5jdURLmdbDBWfeAt7uk00KnFio8pfwbOZ9Rv+WdybdHoaGf
RXTiGSTtBJJuWuJYuYgTwFxhpAjvfq48Q/t/VjDJ8k31k/LHA1EuJiPjQeqLdFJt15jotDWPZpGP
aZ/F4VfGZ+0ZKQCm9vta48kSVzIruXK2gzSWd54AI4S0266IunjqwjAXZZMwdJm7vo4rrrFTC/KZ
vjAt2Jju/Aozco4/yMUgOqh1pKa+KmwMB9SweIrLROVCPrlmG5tPCuFvZpxa108julrtrFAjxpey
SkCePf1gsMkvxIUVz0zJiIPmleNxYpSPwbeEAFsYzETUQpFPJMlfGmhwxRIHwOkb+itapKIk4KS9
azH+S9jQOHEhkO9UUDbn7OjRVXJFbJZj5HkXasqItwaFTC1Mj6xfMRUdQNNJ66uK6274yq2DPtkF
gfAU24ZgZR65cS37kncSYO+rm1Qb9TNKDE0Ax1ugNRPt/QLXN/3iiUUaoT42KwZ5/G0PQdnvXBbq
CiDsqhzUw4v4b2+DlWsNiyr1cH5ii7ggM+GSebse3AzK521tX1MACZf11hZsWmeLjflPPrI9ceLW
whMZJX4fbjtZ6Xzxb4NEZDRrEn4kuz4rM5RChXrlsyDW/M49cUFxLATGNV6DpVtdYCxK1x2O7raG
W2h6mCzLsqC2G+3tKdh2QB5qLzKemg+2dseD/CbvOvXo8LsI3CoWUpeXOVD3UV0gpcylv5eZDUNk
9aSq0aDfPvfkidOw4V8jKy1z4BU5OU/IQBx8U5v9ZmCVKgQZ/xFD+d+x6QSwrD2eYVlxRcgwzySd
63hrGonBiDpLVTcm9ZJwciNYG9dzXO2Lw20eILzFBACL6fopRO15KuGQjr1rF4BeonIs0aV/w8uT
xpwNhZMJ6s8gpMVHmiFMk1VN8EJ0zQ4D2fSGntLyHjOB05FaKyoqVXYMa5G11IFXacSZdwejMsii
6inaEL2JGWuH3IQ0C4ZsMZ5hyYlSdW30nmFBBgv2kOMNVco5w+7WbHcmn/hPQgk1KYExpRec2sF4
kisgzMSNiP4HjL5nNKAp7zWulZUpuEO05cUY8vRU3xc8CwgkN/kAPPXbnYobsvONAMgK/C8wD5zK
luPjT2vPksZNgbt9NQv5GNTXkZ6qdrD1WqjOj0SkymFdyOfe9FPsYvGrZJ33h/o31NNrl0XUaUZ4
Y39Oyj6lPNy+rZWnEwFMCO7UF46OIK46mWXF4vAyU65x9Ck+cZmaoCtlJMstXOTN1kxbr8zb5Dg8
wYTr6bNkRmeTalmw4n9+blFzQneWGxybw4jFV9GqMFjlj6z0SAnpGQlRpzrwkJUdZpJNwHzyFsbU
GF1tt4Bdj9Yaxd+cm512hlZnG0qYk1pEMGSONbV6HOLNOqy3pM8kiHzckXc5xNWM4HK+DYwe0+uR
WNTWv9GA7cmLvF1H8vV2jMxOL3lOrBQY7O82/MUemkOnmMV1U6HiwJm5d0TaRRIK5+24PjXu02Hz
ll88P60FoFGjIFIe4fMm60bgwSfr7CuXFZMPDPnaweFhnugvunT0If1Fb2sEd+jKFT2d271J471/
/xk4U9fKXsbjXB3lin1nkPRgXoSvl2CGl03Psqet+2GzlnuKFF3tSIE8MIXkeiCKTbucht/r4TKg
pRcUG7TxcOKMmvMup48jzZvEHZ0ZN+hMxDBh/vlWeLYWbcXdRfZFlVmC6p6e8bUeyjyOO6ZWgLiZ
j3lDLpft6v7eZYOPqKqdbv7WFWgOVIfvIsheB4EySb8AtZ3MnPhVT/SFKDmzips8dNgC5Fs6Uioa
s6dAlIXYeT5k+aKQca7bIHEFB4f79QAX89Ve+AjvT/WeWXq4QgxRNm3Yo+tOSQCZ2RtfpmxUnXST
caBYMOVSGUndP/ubQ3lWbQ2F0IkKStIaPQDqHEHCEe/Kr0RYxE+bGgvEHlnc6/F2wM1zwy2RmPFZ
L6GPqWjZfvYrbC/pHZLS/UqaXfRdMkWLJ+z05YkQ+ji0yx2yWMbJnGzb2TKMqgSEqO4ZQcmN3T1K
HoJQJxJldbD4QxbZLQnJ1plfy6BkDdXHyht6N+mUiHwOeyCvr85JX7SiSCenIMGXLBTR7o/AnaNa
UlZ7lq43m/fIYxJLKo/6gM/ifFUdDfFsufjMGR8Pr0dqduaxWalHTYlg7mWnVXjjNyl0Tc8DsWv/
cMbnjRXHUWXxVATOlVPB3M89EfJOogsRdtUVNdE7sFVj1XLC8Ku+9XVP1fc3sHsLWJEVJxq4eIz2
iIK6fHKBAND4+C6sA7uEP9DkCl5keiW8HxPqAay0Jp63eIU3hBH8/210mUjmFCMASS5zsEnJixew
Q3lQuZhs9Dqb0TlxG4D2nbZyTJLJ7fLKPXKotkPRTQx3MoWizrvh3YEtvR7fkyBQKFVY8fd0szfT
S3VnDjuszGX5reSeAtemyG6oiR560T3RdJdUCU0Zm6y02QkXJPLg/u6+gcwQCpHD5Ssa1Ljj6DlJ
B2Eshuk7TCP74y3miKIU3pUPVYlO/T7V/sreqMMjSBVRrtXPLwQ9RUdVxYDA4qVHsq6An0DVUtFy
HI7QtQURnO7NbJxYFy7R+ZIcez7AzOJC/mxn+W/Vpjg+/JJcvyVcwTcbdIqlMN8eCOAQUVORfvh8
wZZZiF9/oJ1XBlPAdsGC9m3D4Tq8SGDWa/gCCqTehJVtoGWqS3mHLQbY9mQI2Jww3pZcxaQ61++O
ZSiEkesf/iEhKZbBc0p4YEajq3M5otpqj7UF0tlIB46XSsLQkvl9MH0oV/RgNhPTG1X8q/a76lMY
19dO1bp+ZgslQMxvrcVNB+sD+rrerC84LNcFkPUiZ17KqTxgz8dbjcWfr0/ZePM5FefXKkuMMw1o
dYl9/1ggNF3yl5mdg0emGX3HA4UmN7Ox3tMcw7Nw1iid+4sVmeoSesyKrPFb3QA0pgBz3e7hWnDA
3U7okhO40Qdf2f62/AtFLcwbUZgz+fYmh2h8I6rul++EGGTyqAlbFMPx9YXYqY61jZg3uttnJNDe
5FtolyVN9hRfN3YEQddpDJEf49PU3w2zTQUXDc4a33hhRkdELRKB6NOdz8k9Yt4vGYWVCHewmAq8
sRZOSGJSI3ZW6gzB8MLrxJpbzVSSLbzZLUc7+49SXpmQWdy94It3JXRQcCSmoPHGwAip8E0jEZCJ
IXO6IX7e0p8LrgMSgZeyX0u7OjC431H18vyF6yjSAdD1zSGonsIRzUpA5xaTXwH1qzgP6Sxrnvfr
KzNVY7UHKk/z6mIMTlvbiKVrGIAM+ZuaMXFqKSkL6muiws4IUW7ebi6AjNDBYY/vNsu+yYGXFvhj
TCbYFWzs6z3YRsxaZMejAPNcHfT+JVH3WhCPsKKlXUjzm2rFIYQwOKrZSMPuVyBCogtOTAyNnv53
JOK0lCNeEUEUP1T96aXeQS2d0+xoh29sL/KVkvz+C4DTRKMdmEm9rya1Ig7CbBmNn9HEbq9hN6hK
hgBRgus+qVzFSbRvrDT6Ksv6JHwJm7r9U5MKk7of2l/Nw9p7N9L3sB2ZuUlJKBRgCb72ecmdRRuv
6aDNPiBB6T6AgHHSxx3pl1nvOUNeUsbRZoI4StQR+S2X5Folq0at2u52XiyUoYPxB+WkmwqvEWuJ
wmppvEMIz/n2dTI6TgxilHf3H40mqKQuLw/ANWCmTbdmtPIgc7BtPijU48hZTEFgZlc9QP44Pkfp
pAuLSlduJ6WMPsiJkSRJlfzpCd7kWr4/S6kD5ST+PI8/h11LrXHCZmX/QD15MwE1MDvZ/g/fOXJA
vL3PVqeHMTHcGtEEQjnbupiTqNWlrhHle0VtRqKOqAEcmgvvWOrwMSOnMI+OHnlTortHtsbxEqN1
jvPVvyeatG2FRJoDWyTxOdZQJkAxR7VxOeHNIXMxR00AJTmgYLuKTlXAZE0GmoChMsya59sOPCdl
I6XmqrAUpQzgzkstEiamlqWqXaEfdMQixbbiX6eyJaN5aZ4vKa0PndLq59bkqRlH7lZ8+1ZUszxW
/qbRtOrsOvGNtI4DdzaKohK85/lx/PcM7z97takxP2dhItFU743CRr3isro4H5FuA2yWXqvFMcPU
mgPRAKzz7nzI0Ry9qerPPfedslgTjMMpjt/Vx5b7rhXPft7u67w2S9yMyg5dRE1ki9BTt4vGoipQ
CgPdZBaLGkLKiGh+CnWXzzYBQ1fupbUGI3LY3m2zr8a8r935v6N5g1g+h4y7of+SZZw2WSjWaXf0
jMJWwbkcK5r8qNORLZhTvZcowCM5rEt8Ns2XmxtPT9h4GuX33MlwzfFsVuPtA/nm3eDBdp847q//
yUysICRuxTTxagIuL1D8fcGnmHIeaA30uEzFFytAnKjLz6wkScjL/tECmzKsEHlVsygh0TLw0clz
UIdvO5K3O+B0WiVhFqlqeBf0SN/rFGPJa/lawkvFxiAXdt6EXs3SEJqx1jk29crdBAZc9EXYB8ix
xzqZqwfy00rUK33+ktgRwwAKHBkpbThCFp/uoOo8gi0mrEffz6hUFAv4v3HXISb316L46T6Ha9hT
QVu5L7JrVfHQNZWXNFuJI2P8STvykTxVIV01upZpkZ4+JThNpFhTpiAxwjFRY90uXt5/0T+cHsec
M/HTiSpUQg9kPtT8eWX/RW+VnJewYfN3d+mlj7GzlY27lhcieiXxfY7sMas/KxkT4u3ZZdH0QrUp
38AjS6Jvr7OBekAk1RZxtKIjfup6a9RFuRRVJWKJ175TVlBIfn3M4EJ+2cjoUTuBPvqx0vYGfZma
0li3FIU7YGSeI+QLsQVzD8GR+bqpEwCbnnyWz2Znh4hOksd+bkZ2DcI2H/SsnOOVisPt29HG+ML7
toH8fN3GmPm/X4cSQatdxBlTYarYvj9L1pANIyxAJk20nBQXeuBky367oMmNzIUkUw2gLn3V+SzY
S5Ajqyq/hWqTMGS/oPR3na5vpMrMpSDdop/gHi3Y5pUCtxj5lSdO5nhs6shn2wpF2xBch2DUnZEv
tFUH5Y5Ldcc6J4GAj/rLuGlnMPSUhIKw++cWHVuwlM8Zco+rRRK8CWP9LGTHJNNalfDWwiY1QZUY
raIJVvEuf08t97LxjK9FV4I3tLozNRzJ4JVbI7zqerdMLH1iPWZtWZNtGuV0sN0xFFrakgKjxSkp
5Z57u/Ryqw9aNwdNgdIpfMR9kVvLNcdXsZhv9Q+iE+C+YZzy/+CIjGTnvQNLyrM3d5qGOnF4l2WZ
+eeOtOVNxrRbPKwaVdSf8urpFqsmE5zfz8jMJKDa+FvJ1BEIsWpL/E/4LdsaxGAyGzDgOnVpoqWs
TPZM5dRpzemutg6GBBwrLN62N62Ye6te0+mGCcx67+/kRzG2gyAyqLNlZuPKKSGlLvlKdwFyyLmm
4Oh76KUXw7AH5JTQ4YIf+3eCPGvH3i0Sj/T0a7maoQbnN2MEGdc3Slc92UsZAxfqli+UOZNyJIaK
HNnXEYB/vVGtVKCRYRGN8k+OERZXx3g+dXw+vCTlSVgN/rdLuop1ZWocYTzJNEUkmSPsQIh5ICQ2
K33O/wHgwLdeeyDYLoVsvbRcs7m2UITfVRK/YJdKh2LjanFUXR4zhRydem16nhvIFPPCskd8mK7Q
4/q7Qa32fe4+Yu5BVmIUZ2AbZ4coMoERmNa3heiyHEkHwY6mgpknmBSBRv4Pk7Khdfm9CIzYK+Le
z5DjMTEnmq8Grjp0/4CT3fbzvHyKbDppU6+59wFR3+kexhDIGFHxF31dtevG0z59JEggMdOdzp2o
1qOFNK0d99dKJcYKqooeeEDDN9mjBb/Xczo9dqFQS7H40hJkD09NgEy9cmSe7lHOv0H8Q0cSj90z
smtOY9oocRm0p3YanuPtkpCNTnBVxdfwTjgI1U/eTB3MOLocJmDalnp/oKBa7sF7OQkPsyPKXBn2
Lj3QtvHGVOTmy7cdNiCnoWl44G2IWEXay/Stxkd8xQZ513YMfhQjF6HKKgcNWFjCc93ZM0ZLk5xd
69PZZ94/tYWZ/t6Tzl71LL64xZAEk9BqHpgUoU861AnhDZwCtUHcRCFzI/vOXbMl0gOsplrsE2u1
4lqjhktRT7wi2vuYBFyi3gpiyCRlclnU7T9ojNCEEy9OuYqU9t4beZRmk1L9O6NEuPp++kZFjncz
0bUn1sQCKB8aJ9uCbw4NCn5N9J39EJyDxsfB2i00SRmgucziBjYC/zNLCm3GUxaiKVP01iC1m8sE
juSb3PNzJaCMyT9VCh0laBLIYNBDLCnVAsbjvcNvFtqWIksyy4ocZLQrioQGbi1JrueoqzFWQa8K
8qHuW7Z1wvgy02PYszwtD2ohPN4hc+0V6hfAJrYw+FFAkd2t5F2+BOu3NmCqo7h3rFAJs81GMgw0
ilXUcuLLWxVtrt1hP48gJZOszikk8QpfPhWHczs0FAABcbeRqREkjM8OqyixmdEo+9ZjrbJPAUnx
Y/BrIq2dqe8fBm3mxjHwascvDzMNVOom6+NRfNjWWA3GNF07rK1kxRgqtIBGCc5VQJ055uPgYqDI
YLz/By2ni0bBy7GQET8jZ/ozx4VEOKjPhbexUzcj96rugYnKBXKGCqEJNimL6O0slrsywi1lWaTU
8D8/lQQJOdPCtuEOhVtzcM3qXRrcsl5m0Q1DOVVQVXCeDKBfemR+4MBb9TYVfQSxcwAcD6cNbQQZ
6xe3wzE40Ta5ZTChq9KT7BtvmRlQdKjXmSSQefdvDPprfZEFlljD05q20+q5qXjfZjXny83TEyKm
rxG3NE0xsAydU12gDYkfwc0GLfSJiRWlfw/FcWo2pwhKx6tJn8Bo3DZNW8oDbVFYtoLxU94wh/6l
XtUy26P2b3ystaPBBL46O2HlezCULCFBvmY0B6QagxCtcYbtXj7wH/fQBjtb2zDKss/38vnKQCbE
e0MjxXNpYbfauAgZ7dM06vcN3ESJ6rgw2wA2q+qNitdZ9hxjcg3JvN7aeIcPPJAcBvnKVjY4wpEZ
CoilCceylmCVeKe4jHQqf33Otm7mlWnmLCZ21Bsyvybqk6GQQ/8iuk1v2jHW+QFcEF24OjZhVpIP
i3wrZudaRfrWSbQ0sWxnMRuwod1xFe2CC4kME6oQUZQBlYa52r8vukYyBN7vMgu7ZfEw1D0vF0gX
Y895P1H/0Mz5oKIJGL+PDEQrRTNvwmqUT+t9CLs5KKUqI0rOWkjPkfLgAa3PZLWbEnlCCpQVeCgA
C5Go++bxXtPeX1KinyttvAOcfkVuIXO2Dtla0iB72Mu4s+NC31aHMXhTDkIFP/2zz0aiTd4By2F9
ckIro4hTOgBic42ed9ywtd1psVgr22rQF5dnPnhb9JuDF4c72n3iIuIHg56FiUlgNGrKpgpQy2/f
2lNgdGnhqZPklWNWKZ5jN3EduvN8fEEp+WF1MNkVEnTwy13e3a0aiuMJXni+TFiZ9X+fyReWVx9w
GA9KXVHbYIsqFyTaCrQM0MNdX99fySPA7GT3HoX4pY1bVCxk+t9LbZZeJTZeN3I6YlW7nQANkhbN
CQfwLAUvvyV4KrgRUmMz3QgP90IVXQpj4ICnsb2EmDv/FO/NAZWLYF51bux4/xpSkV4uNJUK+JgS
ATnjWIdI+GJ1vyMjZ9qavOeWI/4I3SkrZxyoz9srgamTN9V6UahtULx87+OvIYsBUzjDaoWP6QtW
gXqN6hG4vR/5fZV05PyMnP8xfSHEmSF5Rx4XYnOq/mAyjEnS+4Y7qnN2G0TVqYB6+1utr21aImUb
jZdRx2wV/QcubUx8yQvSiKa6abA40U0wrQAKI/R7zxcUT8vUyuRIUJku1Auu/ZO+pfyksIVk1eXN
nYh9FpBOxDi2Sug6SuHR7xXkz1WaXRQB3NXp+Xf4gAMwhc3V9Pt1H2P74urj9kpuJqet5R6Xhz4B
NimeqXMl2EAjZRm2Mrd/bki2loUzj1jEM4o2Qvu5a6VE0qdZECe6PhoPBMzvvxkfoenkd4MxzoDA
o/0G/JeYlxAXmQfujNgb2qz6JoyYBukeVucsR0/qxkwnAZQ/CQLx4UcS6gWJkO83e1VFZ8rkeV40
Z04Xx3ajr0MixCx8caQ4SYL3+qzCEi9LFJZGCxf88zcasoDpFTvSoE+ZLWeR5y8s5bWRPpbw2ytN
UM0ZWWrIB/xegXg6JOqAsZmAlMJw9o66I9PM8y+aFrqDckYeuzVKvrar2bVLSjUdzv2g3IgHSKVZ
aSX9dX5Sn005f9B7sMzPgcVBBUubdRhpBLR9lQr6z1qs0l/18qMJdb4v0n5OvszwVGuo7eCi4I7B
1b69asxt6UjiNsootPQ/Wc3h3DNmqU0uJhh4CwKb/1rysllSamKONeyO33F5HKn3F3y+hBAulsTj
G7gfbX/csI+QIrTQOLVzbkrKd7nFT0KT2XNLZbAaLI5R2qz84qDYWK3elTajie0WktfHocS0bOo2
vFUk53uUiVGnnwctCfpe5C6HxpnkH8ViXm4PNvoZTX00bu8C5V8glEVfHCZrJiYydDCUNAoPNRbD
Q3ttOPe/GiH/dU0NtwWvI9f+C79Lllt+WHUTKBStyBb3XIVnDleDjBJ4z6jXL+pHoYnW4lISSwTv
vNM16fDzKSyQaJt6P8rQvLONbdrbPKeG2Ec0Mpa+Tlq7bBWq5jxdnvPa1ux7zZUKsFYiy9b7PXPr
Igx+li2+lZ349aOcRtMMI9rKoVStKl8I2kPtZlvC+4d5Q+/P1OClSdKLTT5vycOGS5UxVfT2JLM9
MaxeVrBR4DBu5cDP6ixsOISfe/Yw9ZleD422AO1/RXnUeJrc5NUWum1EQkkdRX1kvyW6OXxLyfbz
wCGkKkt7tW7Styu/xLp9Tn/4MI3Ow4ubr2n3SJizR/XzK7HkaoZ0Y4u8wNZZhvgzpcKC+aFxJACp
+GcH4Cu4vtEp/12myl2ADLbyurdkb9F4EC5n5Ymx6Pq1Tb/dGFurE5zffNAWksgenzKz419hNWYV
++pAl9Li9MoYZzS0eVUTeuT04LZ+yHlrDiV1lu4fuMzMG2pQCcP7TyNzk9nFHTVrHM8xb0mgIHrL
I632nlsr7R9wIxZXo45PQ7GLfV+Hf4n0c9EyRZYI6PNmKX8ysmbYMzCjX9GK56RKtiaobX3yLOj1
ujPhP3e5GofmvzTEtztXWxZ65EOEBU5KVtqpIHBtRrcE7Z74QM3zkU1cogq3gAZnW7bEyvA/lqz7
Ga6Y4aj84tyKTw5c8jNJzqFAkpw+vn1CcldH0HY1/iEfqYavaExL+B4OAJXyO6ohCj2sYiaDvBM+
aaROTg4cXCOrIo9DnT7CjNQtVWN7fW9KkDD+NWsh+iZbsWwZ4+lPMhBwjK9bA1W3qSgDIP8XMfTF
sfwh6nNiF3WKYmuEUi4Vlyyybe5Q+GBDjcAz7hzf+CiM07furR5i0mcLV/X4cVhs5Tzr4myIPP9w
j+WRmTJY9wXMoGagWNhtvh3uKB34w5JcJlZeXbDQ35vY5gKfUhewvfZaCqdgCKyNapUgYZe0DAg6
3kasEiKzO4yL8M3+pqJrjRWOcBNVXPvt0x0tRpXLPQZlVZkzpSQCsPDIiQKX4RzDdQZB5f6+ngQE
hDZsuguIlk0hzj8NiQooGzQcI5IluWVoYtlVkbNsdGkuG6i1CkyCIROXFtfAiGpWLkg4/MrGFS0o
2pjHODgB4+DcMwab5WBu0UI0YpdtnsZmijECGrjRuM54iJzvY8/nPaPCSrqQ2SBb2ih/cDyH2u1x
CtaBJrj713EWpaE3t9XKJGxk1Pc/agb9gMjCy8wTw0xphehsD1juoRjv+xolVkQ2+TmJ7cZ76shW
Wk8UbX17nTVSgf+pYgY/jq+eyAiKiPdsOnrTBbkXNZCulGLfJb00i6fiP0q2x2RMbpfo1+fzlURC
IsnzkRbShTz2EArtqBnKTocvmX3oYGSFtv1R0+PI91Ur9EDB9ReJ+xTO7h4atH4fh4Awcj/80+ZT
GhgUdNVzoyAhMfCfppWolcu7vNhceBobPYZko2GfLhiBU/LoiNX5ibCcQEVMLR2ZYugjE4az6bJ4
F/o7qioBIL7yl0PQp2W3RGWkFRuR+5pBaci7Fk1eLBUKUtFu2rNZiqjBp9mGsiwl7e0FgzQwvvdf
9+nMTjRECvdu3Y3+Gd2rAyu9jE4rHmzhXCCRgfI2Eltm+MtY15DqEJ91QPXc9AuJgJW9dTMZ1oS2
e8OnbKidJYuuvlaTO8YEg1yEA+cA8e0wft1UYU8KZRae5x/qJZQnOOUOLiwE/7TugVQFHZtIihzC
qhZu2h6fBDW46UUmk615SrXHjEr+36stCnITjvbhPiXQiAJOWLfOXWGxpvNEpL/0s6yc40Bo4Vl0
tAdNv/wPs0FDFCp3s6v3dbSNlYVWdpgGxrsmU5Tak4dRifCZB82VVS4bsfJlI0LpsP7jCHtlEQAo
m/Dow5cT7MlOYy/LGb+THeX3vyqSmBDPH5bCa7Q+kXdEF/Y/gRSGpz+O7LUt2+pY/QO4svggSUz8
tg40oI0XYKgMtesSUyN1ABnVv3sk4fyhOGopSha26yq0D77gA+Pe0ppbrPZr30LdO+zoruJhWxNZ
DMfZbs2wg0Uzh/V+kfsU1/NkXZn4TevF3vRp8Dy3bURYiHPFKBXbdEk/KdLDInmB1XHu5FWk89Ly
q0HtNGgpnuth0P1ShhaG8Jz3xrWsGtZUUyYoqetyG+GCpmcEV7jFRymE+rE0L6rddvoQgsf0VDDN
oFDJ7jmnewn7RTM/N2D/k/p5DoDM7AfQH6k/650TUXn8CUT2CuRohyhEVAiNWrVjxZ3EhTsdRxeI
QKHcPpQCMyYc1OJsBrtRUl+vQEfkdB4z4hhzCC6jbKVG4czgiiHnV56HFYXwzZkiXvWbXP3i2+ki
hwREU1b01r3x/Ek+78g9Divvv2w0fscSoGL6LLXy9phbh5K+iI4KOKJEYj9BieizJn520S995I3H
y7b58rScBE7riulWSdjyt5d4+gS/3Q6yxDkElSjFWJDHUtgwsFnxukSQNwFYJcayQb5OaZ3TGcbN
a9293BmPGcGNPVLpV24EoAvR8EGp3A4EWAYkQGDgzuKviguLCZuhwYL7QSgd6c78Oav3U9nvizct
uIEDJ+kYJ2wXY8/vPtvunFaqiEaadCKWxo+8NAFHkiOZLJ06w7gaG56tSSSDTF4nGD4tD6OW06Y/
Gvga54/NiTZcbiZWwUvdSMixyobSUyMVeLB2L6D4Gxugf1WqJPzLnEsOVFL8hgXLjXG8QyTREQ1L
5wVZ8A3vU7aoBkv4SQ2zRO3kbSyd6b0v6X0jwb1D86zziYcgar6i07reXUC4eGAwIciuHdttxPUZ
rsLcPxQBWMLlJPvyZa5tEkRYQK8wUtKLYlM/Y+M86wHLrJcJjL1RihpQMxOeBExCzkCzMeMHwNJg
k9VKw9xLCbV7o9Ly8u4qGT7QeCCcj8Mf5HGMUrQRSyA4K3uxwj4oa1OYo+rn9dsuqDUFTrmYRDuN
vYEQIT0W3CU/k4RSwUsxc4YfURacGNcWk3SSpjTjW2s0BMBxv+QwRe84iUQzdqqIe0BysR/WPiRR
Dk15+fnFHXuSl1t9GjfO1oMdkB4lNIi7Zx6RjuUtD9PxajABdvtinDDv88jFKB8A3Vc6mN/6UIM0
PiLU2kZLc8IVZ+XJ0+k9vHXrHzbXiIOCq8feOkXclrT7mg4R7KoCf/lgxG/l0rZm7ONHb7kAeyhG
KxN3n4PdFPn/k6astPq8x3KzHvy5K7Wro4xoCSBkwiswQRwaee55RsQSa/BNss29D9Eshx6PDuKR
bqOUgC3L+1BU5qSbW9DKXRQqkPrbZCr7rxEbnPIkbgKrPo1laYPEl/EPBkSdI0Gn4+TncDIrtkXW
wLzuyLd/tCrd/GCS+w34BbgqxstlpdcqdxntDJVcbSmHrOu2jTOCIFNKx+nxKJ5ymNTnhzbJQ7sR
IRLV6HXtOUBv8XF8rrTgjv0dpzpHRZJmYdraVgS5lRBpWmwnY0zqdhmn99BEDG7dNvXQVpfbvJCu
KVGl0TVTJsRubRnvosagkm/BqXXbSdVqV14N8ooImzcG938C8Em7avON2yxbgC8CT4ExTl3ZALi7
NWCKDEKI45R1iZ07RM2FmImG30ToadBOO2YrX3f6cQD1g3WTp0/5KlpxomFmK8ak9ij8B/M+Mv+f
lkp8ly3FCXyTQB2l1e/D/1IbMly/OVLfLCSG4gUWZpKC2lVa+U/G/8uuxZFOUNpn9pQSBKHq5/RF
fO2/U10sA0cc9qhfHWuklEC/JhRP4DVNl2kARAFoGtT5XYLbaUXliup5cVGKpY29tDGd8Jq3oixh
9yKd7S+BlzqVoD0c8KRUTFIHsLddxNZYT62Ob/3SUSG+hjbCVLQPS2a7eFto79EGL1sblxfdPtYM
/BXR+/AsarVfD2gHHu0PnZj4eon2bpNFgAw0xUMv4d/VV+Ar5kPwjAlh6Nr73CqBhAoRVyVpXL5u
N5ZMEVEusd8mNDd6DFiGKMXFdCmhSwkarIVZfZbHoXxfayOYaURUa4KJ5BwHTy42TUjSF9fn+8vl
yHRgsq4rZk7ViIop8IJUCR44nkjByGvkt7k5Bcd4JCMqkGdJuEduUBtmlTyAGxj/1tm04eHhpica
vnfXfPWWTTwsl8YxFbbxOnJeEp3P+GBaD5pa8PmmwRbAcNqo41kGmYySGn/t/R4dkFaSWngxqQMn
hBdzKHUV8lg9SKpoZXP6Gs2l3a1SfpxJJQ8U7VgPOPvPSGoUm3sQyNigfOvfOA4nxntUOPgOVERo
d1vFXVFF75S+xQYJCAMu/SDuql2sFW1CtX9yh2jPCXMG0XGZoPNU5zM0JhAcf+6cMxX8YFwZ/ljP
nVI5g5jFtSEoKaZwzNnq7T/bzXvHgc8H4ESPIvWhZ1ObECDU+Cj8WPtqwop4hCwlTqS6mcTGvkdH
EFY+jf3DckMoHxh7ijnG9vQRgFJ26tupDgt3GVeF3eTDwXY9n9s/3tCHzoJdmFXeC9fUvVozeLpq
rocG+6wCAMQ1PzDjJRIQwA4VGpmCqY6NSgXmcMiQ6O8roUj5RCJWXb+svpETs4oVw1oGGheCkoV9
AXY8ZiVIyCVutUG/2vwd5RZAwR4bBor6MNd/9D8oIDgpzU89yPyK7jp7xBomiwlIgrqYjl0RfJrc
CZG//Rr/tqDT/zPLeRDsZn3DP55E309X9qANVjjw/ULSNgakV5v8Jdehi8yJ1xX4PNJrThCR7q24
nAEg+r1uh6KqKfqVD57WFvl0tPpwxbkJVnQpP2nNys8Fjp05cZha0I+MVuSf1dhhlkboYWiSXlA3
QQ66kMlp7ySgLBpHTPWyADZQlY2t8GsRV4ME2spWa106ktVmNecuB4D3DSfEDnZQWn7IK5GxZ4o4
LJa4sA2Jxgs1aH9AZbKu2wDOruh4zgmD3uZ7d9bjLasNKCdOZR4XcbUaftnPoAth7z9xWcOBzvEZ
6MAkrCjBOlG4StZNIahqH9cKqjTABFIMu+EhzkdHl30xwvdk0IrU9Ohv0+oAQ2jr9zVLfvBRNHof
Kx0sr7A6pux2tOMAJP2hStAc+CuKdjJhJuG2gohcGhAhB8We6TSyXk70GGq6A+8Qc2ILhnjpO838
ooQ6li6l8GBPZewTZ87UH+Q57tKxYBR89fFpTi0cnSkTcgISGpVXDXXkw+RunZP8xTlLs9dc1BW9
K5wkC3TP5dQ9NggeStYu6VzHk3k2rPRUJyfGMLVfrr/dyFTcIgjeY7TSRDqO4oBz3plLmC380sqN
wWbLC/gO8iWWsXfeY+W0h3GlcX+B7tIBYfadn4ymSjxwa81neLv5J1Z8j0heqW1Vp8B92rVSlLUd
/tjWQO2FANjjd+QfnQVy3f1PYsPl4+FD8VGh9mpiiMD6HLiPp+HH8kP2w+17JAPdEv6H7OytJ8BG
HdKuEbK+uI0OQLqCaCKgALS9L/Ye/Fn30mFVhtwcXYujCrqwiftij1X3tql/9vu+Pgd9PKJWud1s
tPV+p+Mk9m9E4+ORnoPexdgLA0fDJSgrErw9kGx1OXLa8TAaY3xNpB5V/t+cFNEu7DfBDsoAkUll
IS9x9x0S/3V1gQZTGJfA0irXE7f5rKcPHBM7SXSn6DCJq6URf6Fk7BqOjgdCl3q9WWyBCSRKBs7t
nTNO81bDxMbALIbcuihQpNwu9dnTQe7DYbBsPQYSTI4dau+wBFZWq9WL5DJCCG3gWxJ6i1J5Td/t
WvzPOu6ZMU2pEM6JT+q6ZqqNASbMYJxldTUfnNrOolTkauNYbvYzJ+B6E9k250K3SwqO55GCQYlb
Udavp/5Pest8hlz+LpCWQGkUK0ALXw5aUcfsrQn3zo9TV/SjSJSw3o4dP1ZbF0u2D6dSYDhIotBs
S5u1AD6/dZQN2SjmsW+JCCu9R+FkLHTmWb/zfp+4QHu3918Dn0WKaVrTqEBhdXbdwpwgHpJfQMGs
t52C2OLyE7oOK+BhahfKWix0I1pKmKudHcQMBASzIYIoowwxUgpFBAW1ovVNSurN7OnkZcnTr9Gn
FiyD6HM1bKWJpg7mSKe51nVR8i629U4W5D7jjX9lpHh1BiGQTg3QsWqAurUDGOD70NojhJ35772z
pPZxCHYH7OlJWVQs+sEj3m52U8GOlzLb88vnTFd9w5L0HlNM1g4uTilfO3PLl/vYAxN4JsVbFjny
/+Pn3itkfSElMjZQkbPggJrR+STvIVf7HRf2v2vk5aj/zB1/Bj/jf009IrKiN5bg4xzndmSfZVqJ
RHnrzJTnNUYeS5CjIsKDGqEMeGsOzaGJZLe+/dk5tQOJcwxrntDgP2ZgY4xG/UqL0ajTTT1mLaOJ
IRIORRBmrH4mhDb78SrPhDDJEceRat08pnJoU6q6DkpOTf4Cr8gmsGbiAjrUkez4pfJbuvCYbsRi
rpY3Na1mrPa+JaqjNN/OMi3AbNn3pYQgjpXdqY5E+TKFyefanfuu1OrUyPHaLhvuhqaGCUG26X41
QFOpwNGbGGf4cu26jJ28CJvS7MZ6MmMyPTS3el+8Lxx2UFLTVuu8TqrZaZ4MO62lIsMPWbjWl/1R
GHo7r5Inh8LYbvQK2eC0BAjAt8CH48QC8H2ETcghudZE7VDLm/s8PsAc+2H6WAec3CH1Jul4Zg8/
5ZFsDpiCtxMdnqcgYUdDfFtEU0/qeiv3qNaxMRH1UfUGZTuhgAnKk4tsjv3MtHrijEmuSs2khDUb
9IAGX6DVELmIyVtYfX20CLJMkpc6VGbicUyRRHYAZHhsNRQEBIxJsiQZ53Vs4lS/wg0zIarnRuvG
U0qes2YB5NU7oty74IVU1VC2p/QrNGYg1v2e38QqXQkjBa0V3Yh8HzoltQA/nZinEUeGnboU9UJD
x4qrf76qAfqH3bjg2a6LsQQSSJaD9XOa4rKaM38TZp3r7CLvYLBHQ/8oeNO24wZc8hQLYeZa4QNO
s8cT+8VsnQdI22HSP71PCWaS/KysmqvOA/5jeIfyQD++yHv4Oop45cDR33l6u86Pg+ny/TONhg0m
YxFs0LTo97JYVvT+UDlNe1PmAvIBT1f12KTJIFqgl+8zBjNADoQvlQlX7eJn8LQTQVB36MdWbUO2
pt2PLEsmtzxr888Gfk41Zk2Ix7JAdkiw0MOr8Oovfxpzwlo6mizd/4hqg/II5TjfMf314TwuKiUs
Sz8pKY4Ldv9vcMt1GElTLGNHiKE9+vWOwl35A75v/KlDSmdm8+g+zEhHCprhv/np2cyIj/ogviD+
wdttwR5MSP7K+gV+4fmfQTpFGRgF+PYiG+5NYKFfG7bFWrmzYH6908JWgtQR/ThkpuXTEUyyp6YK
flhDSrg+a+BSKqOrspCPPkDuzCZJ9k5nld7Kpt0qv9SU/En+cB8KONQYLJUXZVLpV3XnMgSwjWHu
Zu2GADJIIP7dwdbygS3lyG5qi0vIMShvoWzXGppU2mPSjP0R7SYy+80iKtFxkPzzdeTwfgvmT0EA
bmJ5Jve7ORt5sbuOxhp4CCyqZuABa6gJ1Q+ruWDXbWSjjP+RL/8AmES228Gv7f4l2s4APz+hrODj
h1bdy3YEDDJcs/E7oW1WVWooDsjp5Toa3tHb5or2vo8A6SEPMeFkt0FWPIjzHcghxXIeCQ0KqQyZ
SM1jH2LE1zN7S0ne8bWB80VBlTyfuSjDS7l0Yzj6lxdwvuRZle46Bqw5guyVtgsiMM56vu1jU+bE
yccSNPPIV0ewcg9VJ/TYvUZ3dy/CmnDY5ttXODFh0RDZVmCzd2a0N0yq5uiPVZZUwGQz7Bwuum/R
nz8UKoMZ5xW2o842K9P/YgPXNPfgqm3lFIuBejo1iYOymbhzXjqSBzJFoewsJA+1lEmCV+nTQWuX
o0g6c7lnyxRz4+iWnpxLMZLUkeHQYy/HoUXhZCm/5nsO7l0kCBXfVBEvDHxNVjn+x9uP4lAeafOy
3IeiJ38TowzeblWns8o+At6weH5KYLegxTvwpPOcs/bPqdLmOVkLbSKz8LAprYYtsV0mHCNDcyCr
+Y++e9VvfE2gvUe51puVlJGxCpraZCfKFVDHOt8rb9srctzDe7i62KrIiC5e9I552/mkvykeeHx+
RbYc666TPTA6ZHpSIgPLBaJhEQH/7vsJb+dwGDv2Td1mnHIWf2nDkxdZ+Jds5HKUKKrLIFIIcS2V
IpZqYJVY0DskzpXzpB1PRINBhGCwN5efx9bcNa96pTWZph/rbZXmo76bFuRHCroC2q1ngrVVhOFM
M+gRc1XIRey4cdZNdi9aeuCK1U2uFxBQt8jiDBIveKThDYppKATirljmmzAZG9raApdObwkFf8XA
vgBwd2f0Cz9DlMsypG/1LBFt4CWcaLK2KUoiyixOlD6S9h/utx/WDlu7HYembsXqRFdWpPscZUOu
BGqMIOXRuXcHbFJ1R0yT8dQbJGiGYsNo5QF5JTnxUm/9155832yhP/Ugqnhi9oPDhrg9BG4CLXJw
wyVUpmYj7aK5qwB28iPLMryfTNkeixUCM1Zu/CgO5uCvU78GU4SWQAbDCycsJzJoPgAiTbKTkpc+
eo/Y+phE2/EAIYR2xcevOegYghc5ZCN9ZVSNC0hmpQEuwEnuhmMcYHC9VUGWE3rSBoF+ipE8ypd8
GasT+BWq5uRDXPXQ4eDRQvF+Al3LDnVOWBZeUkQlzXI/XG53hlW2ckFjLGywOdd7yMZOUtdX2CJF
QUHRYfNztE8n2LUFtTakPerkkqQ9RAJtPwd/QHwE0Tszbh16bLaGyxd5v4t7BLzKpChZ3HMf+T0g
86iPrxK87E5T2Lt07ACYB/EPVd2s/P8dWe1nP7P+DOIZYamo3gR97g3wsklje5Cz3IHCnfJxrvUY
tnF/RKdPZRYKNZGF5n9Jw/AxQuh0FT+FZ89Abx8x9Cl7QbbVzu1SFOYp+pXbJFUeoG6JQFN0F52f
7I43WF8kzGLmJBOVY8QQRSEiayMs/khZ/ZvGHHTYygRB8UsGj0AAq7D7AMc7jO4czjLhUfD+I8xG
o3PsnjygD8BozbYlJpNFWFdau+ttHLLvPxzypWOcCCWjEgRLnZMYH+Eh7AyVVKqIsmeFxfaIxDvI
ocJixX7y1591Eq2HSvFL+f3Js4yjyErpEwyDiK7rf/MZ/WxeI18SuVoqdlWy6mkFgciEB9d5MEvy
C/VSk59ynFEMj+LGBGz4P5xo5EKS7l/YKfaYhDhWGXiPzXtBNfpjhNe5rIPkjVL6EVgK2i8cekxA
+oAV1vXabIMNPJFj783fa4QUf4m1eX0UJBo+wq8NN0OMlg600f+tHojR666bbHbJVLA588hKyY3v
J0XMerbz12JLfChO9EE+NKtQXb5hBSgkDgCjPXqiFeHQP6OWxi1W1GcplRDd5PztZoJpRhdsuyJ1
XpmVljmHHR6I/P35suAhDIy8zc5yyHkoOzk7L05e39DsaQUG1REiQWyhFDM/drtkgPssJBwOFgrP
NC5ODbEX5rV90t5yXHALmtB7ZWQBlsaIMexPEFoz0I6VHjXJp37sEOchyCukNDRvRm3WeSIG+lFe
JQFFdhtzrOkOf81QAtA4Kz/p+gDVqfJJIrpHiXeF9EIXnr0sL0Jpjon/xOXZqZMJ1WmeDdgZlOKI
gyJOIBsB+bw4/jEQ78Svsd7D/o13Je8eCZCI2qmwWPTIEC9abaUmc6gyPb4Lq6CZ7NE3JeUrDNA5
YMNG+crq5PwpJLSombh71vAw94xXSqEb2JnnTB2xBkSfDH3XayyhC9pGlzH4VOshn+JPYjZFdgpH
Gs44eDyzHMZTzJCJbsauJraFoIkW9/9nDQT8Y9tlO84XQ7bF0+ooZsUGwVlEqITAtn0opXOr88EM
kcS+y8hq08bt2lpiCJgsev9hi/6AcFa3gaZkJz7Fw8hQFiVVJ0l6Tbz3PZ3r4OmCYz3sOJRX88YI
rz3nFHQoYtvCmnBEGwV0T3I8dU2ZQ+U1tWPw6UamyBO+qrW9gCVqaSQAnCQfa3YGAIJQSgH6qxR3
ZGNdD0Kjx9RrRJVF636TjMhQ4Hu5tA0u1SZXvU5Bgw4FgsOus4+58/xo3FeyAUsXbkL8xL1ItuUF
suLpMXho8hRl0URKFyNFlmFdWrM+aiw8NPVzRYTMLjRbJsnVRaqXe+EIc9pBFUSUj/SifCBA78s2
vQffDEqQkEI6pWonBo2fu9nVmvJrqjLI/oSlRCF0AI34ndNSjBmH4p/cTZ55r+ugyEoFKPd+qrdG
jtDggg9dBa3augtIPtPRa+5p1ODRXo0s+AxKtgA7Fz9nj8h4iuRsaBHeZ6I6nuDL1iuMeKS3qt8j
qH7NYeYFqbVQFFj+j1Zk/CvhrX0WzM1Drjesapva/UIPhCl7CRdWr5zoX2lVZkxxbS+o2iINnV/9
Pny+LB5ZaSEa18SEAxjL4bGYAEbOO0w5xDlB4Q4ABvkXj1SuQdFRV17L3ZVyeg6R5Xuh0eeTWerV
twsMavppxbSCXlnjIXLdKPJ9rnr1Sa59O6G8sxDaDhbCOWU86MdbbMTaldJ5Bc4nSl70jWrf4+aB
JFOlcnrNNAl/LYm3KX66Ku3GwHrXXNFZlaJrKPHRohb4LVJEy0B1/VegK08N15dlGII9o7nPOv4y
pvsVt1278ToAxzWam5fKDHNF2xCoPKMBgNIYTjfFoKeX/NGlK3wKrdUMH66INSewD/Zy/yqIsDN+
Hxk+fskQ1NT6TzSLQEo6Ls5o5kUShXV7grqEIN6sb/V3CMMfCQO/EkOCn2QWC3TqAz0B6067TDXP
di3ys7iZqxx8TubD+HCZ8yO2SFr4p0Ra6joph2HHj1hSbyLwLchMhkC2ImdWSTZwlpzBydZ4pcJl
a+nCB6tTCkNrA0YK2Rv3jY0SbyVjwvphECubVFf3fmh8HZbnQ/J9hpd4MsCCbEWf2a5FnSwyz/Ji
hXqgjIUrfjDgeG3skN/FAMpSoEObSyf94f1JiByvRZ5c2GZamgwyzss/lZveNBwVz6h68qzUj3+I
hMewJ7304OQe8jsgFUIN7x2mgwhGa11xam5KlPoBAFo6NZifRwa4A37CGVe1ChN7S269g6IcC8Zi
/dHYQCQdDKLAqMILubM5M7ZeoVdZk3eDpH9ITp0WJaScvLaWDwuk/4EuxKWFOmyQ7NtKiK2CvwrT
RWEhU3WYQKejfpWoCcI3T9K2+CJuGcZ6op+zcV8NqznXHy5n8gz1Pa4x6zRzwvLIuPbtYiLmSGSk
cPoa6cIjOSzXTMfd3M+DR51gYnkO1yIB6Rs+/W9Dn68cMiGyU8sDx51ZuvDb/pj4NNPmJvCvLUNy
cems4QicxOCu+GhfJCgFpEgG9wNeAubo4k6wQMAXvfr2gCGwMNtnc8MylVRQzqpNo7KdLE+Rj7ry
RvEl0j+vCPPwvzJIWNbvIo2J8mHobs+x2c7BSAvoKpS4j4R1dTmMVGU88LOnuDpsIvNos2GeGNj0
7mTNEEM7V4scDEIffFXcyha7q9y82I64Q3ouawEwxDpbAwZR5xykAnP6J8/U7eKypHZeWrYtzMx8
/EZBUA9giDf1PZqCBk2F+2psWTmC4+WY7oFZrVFnRexMigjV1qNmsgdrZdM4DaswbeKXDF9SUm1u
YcOPmjJi/ep4qtxr8OdBAkukuyzG8CSH27yIEG7rmQ+eMn69zpVlkMsz3uJQ+YUXj+nfl75EYnje
O0fksurGktDjHtY/nD3B3h77cKHE8FCCm/ogM3EMvagC8ilpM/iGjMabioqaID2NQVUOwB6uph6p
+2TV1pPsg8DuGbajT4pi0gPNnbUEX5JJozkwxesQntbwNydbeve9qnlO9SqSxlo2/lPtNd9JcvUF
oNsetjWIWqj37y7pA4ykJDG//X9aX/6QAnjyl8U+Z8e6GEoqryMhaqxXKiQRJkLP2UUA/OveKEUR
z6OHJ4JOz2jCO3tkRiiMtplXcZAG/dmKnuremv24fmEoV7j8B1+IWGIIFFI3f2wE+px0zcFkTTZ6
xHnLdp8kQKj1mTyTGM4ZBd/EWH0vt7zCyCAOutOrijQQnbS+Jc7z0OnPEo3ouXNG1S1YrxouLaDW
W4mZ4SLDseVun41Yd1P/CSY+i/J7vtKyQ2bDCXB2oBfRNK+nKWrWmmHvULPnqxxLML+2HOGb74DT
ZT3+KnddObG/Ue2qQn6XSphb+p/Wi8uDxl+4DTUseJCKFpg1oDzyFhvNtcNiDrKdrL71uYffEHmt
JdK2lQaoHErEntrHk6KlOq+kANGRcFhmZaiQm3DB7rcgIYCskyzwSlxcR3JB/knCBnDRQA3uBX6g
g8JHf7trwlBD2kwjpqe17HNbQvz62t4hcpF1MKlSJxHC5CT5TJ+mp5PMpFRtuOOWd3EtBylD5PuE
50ALZBxJpG2tbZol6pfwv2NUJcArsJ4SJXuj3iS5aj/kbBqyYDfYI8FIAulqUDXNQLYGwNkQDHSZ
XE4aXW8P/Y/pRml7GR1uMiRlYoDCIsSd8p0x9ALsgpz2pPkHW6a744qzn3Q3ac5d9mf2su6EZChw
pa5l6zCHk6FRljBO6Yk0MacecW7U8XtR71yG6uEAvWzTY/p9VqbuYbJ+5B52CM1Qvgtiu1Y3I1gH
1AnP/EkK6Z1n7XIS0t3Mz+6w5ztXLy9W8KFfmpdQG3c1vfeJLt+tuAmvnGDLTGhyMRai6GZi/B9M
9lVhEnRDVLnlrz6DEfwl0SslTXGSIrRaezv60MJJbsu8cH8AK8isk1hEeXMxkW45lsoOenWP+EZa
tnckpZ+4Fr5YSTE1JnMzSkbSQE5732nDRjkgJOc3uS87A4jXiAa3hFcSPbrrEmoxPnH8mDEKszjb
qclKbcin/6oXTLCT00Y8cwgOCYbUgbksgLa007RoqjfniTMo+oh76x3GC/7V7xFJxcV63K4RPZmk
CeoQhD0PDgx4Vu13/pvgGbkIxzN1vfYh+nDz0ZCxIRuFSNkOr+vnoPO1eXgT7Ap0NnoOYw/XUVQD
JbVTnV7WUftqjs6zkvqs8Tb5IUCkBNbDU3MkwWEkdPeZNKBtNlr741hG521BjOaf4DGGFrX77rgZ
FGZmoE22TIk9ytBYpwxAlLFdKew1STrhn1hm5brDyrowwdFAi6E7q6wsb6Qz0s93QlhdII5fzMul
wrcChFhM/lE65a0ZRGZ5Uc2dL+P55GHVCmVfaNRYGOQkhohLBxn3z7HWdUDfLZ6W+HBB+mW1SOMM
5VBzLTduh84r/NamSBnUJM4UN71o/4iVynYtJ18RozN1lUWmeJUa3Pw5hJDQPsuzXJMUZTxs5JOB
5dnqlu/8O68FNCSgpoaPv9UtCGJMNJ/etoHYENEbTyv0bYmzBXNc5Cn3kdMu5ocx9YWEhrGTN1qI
5hyNwlY9Cf4EhMUxxTxFyVLmL0FeCg865JfXV9i7kJj2+0oqG6lS2TdZUYePZHRg+wH2DqKCcVYa
NsH4219EZWlBhjwzm0oCppQ3tqndf/Q1zb3qqxPb4ivAlVQt/3akERbYb6R3y7dPTdCRnRueJBo/
j1ELDEUcwaY2B10hQDxdDgyk0FbQVrSS1RH+GhVVGljB2BWojfaWaqfv8fABLXkCGuWIqux33yE/
nVS2mw/lIyitR1CL6lKethGRlBKj72WrwfP5mNc015GEJFNOUYgFKAMp6s6u3/4Kmz+tLe1FOy18
azhRfn9e1zRCOE0S/tRuNr133j0tnhYy9ytMMzxnR+YixwUo1GT7oh3Jd3xHrIIjf0nDVet0KH7F
T0wb0WquSjEg+NmoHvbJfZZRWO6MhQRYA+CBmHuACTq71KutbXoTV7zQkqX+g57dwXrjLmwMoMlW
SxY3U+3yBTsIXL+cFG8pp6gOfQ4DPjUK66NaFxacc0K9ywlwjkdOCT5my0VOWQ5co7NgoIoT4IUP
r7vKXAn2/RVe6I7uWIvS5yMUChYV1rDzdOrAwv50/EOdMtGcgwln+BAwE8p+wI2gWwHGulxjHz7k
EpA+IR/jVYIfC5cBOOfl/0r2wKrW/gWpv2TIRTMhCgrf8bVYk4XXY7h9rM5tDYY4gF6DF2fbYBh2
7KA/X6FjPH72Ubusnz6FhV4Ztf3AdlJTG7JneGzPNXu5aRjNGbAVFOb/E/iqnzNXiSyT8W+KAxIr
IuwS2vh/Egh07/YiWkvVebLTGNWEUNjnDHcjTEHApSXeRzH9+T78EqkJTgEoCUfH271NMEXhQiwf
3BxGHr1cwJoqm3/zuKDnWo1zMBNIOZ7x9/XDhFP9k/JCu49/ymP4Pykt9mo4sOs/Dv5TdBnGqVZ6
lG4Tk5h75QOm1u5j7kj/zJiSsqJGLEsDJr+OmSCIK7mtEq9/fKoriBHjbLk7OTPXfSmFLmWxMOcl
IVK1UoZO1xj1K8plRR8aFI/iz1bhqxStDQjYZb0HNZqxg7VhwHfB5KfWE5BmuHJbxTHVbh5dORJV
ZRHA4r1Zi+RqdnShNhG3CisV+fcZDDrQmcwUAYiyo3CegjCIkHEpiVJ8Mhl72KWsNqsMELA7KzBL
VHFyOcLRDlH7+59bvYdPfHC926liNy0SOjOCpSV/c8f6DL7/wv4REJmR7flw7KzBGieQqDLQt/Uw
znaKByxEJz90ALGmuCssiUEvU43fevzfnKcdxP+kL17nlmAeom4DSQ89JThU9kTlHrxPPIeNQ5hT
gH8Rapj08R3V4oDcvxce1msnaFEmtRYf30WOQi37n+NyYzDOSCQ+v+V4nFqAGHd4tJVsfkUVmPIb
ynAmjlO9zRHvDMX2c9+trhZa4PTfU18u9dU8XQYnJ4+S/DztUD+nuNGezGpVRXeiGAqDJ11+sh9D
hERHe2X9cJxXSZk6Rl8xywW3F+uwX0ryb4pmkH8st+ObP65GivdIw1u/b6Sh8yKSmuPWM//mCjnS
hvceF0Z2spzPdpB+BHBj1bjSoxldtds9nSQGcpDhXeBiMiY2ot7OOAk1XwzRphqHBo+JT2l8pQ7Z
JUGXeJDlY96E2Q9AQDOGDh2eDqlvfeGN4sbsaUHUoUXDMKy6JKpEHUjq0N9ziH8KRfJppfLxzyUm
tVgFb3Gn55vnn2JsQNgNSZh2KoQHVoIflu+bS0GjJRpDV5XoJ0Op7ZdYxPmU36CaHgNNvJLx3hs6
TfgcAVMmXhVuJITw5oPfE+HMLP3ngj6vgwEWLvPDyne9x7rVZEX8YLTYyzwXYbN+uAA5XIAm7bvf
Sv91SXk4Rn7z/ZUp3upkx9h3uk4ZJdkHpfnod77hnyOq4TAu29yOpc4UVcZLZ4/65VkVFfIQHUB3
nnjsunqHjLBiK0666f5of/UQdB/41uynX737svNagFUrM085q3BUYsEvto/g5Akwd6ZLpX0jabnh
yuVLV6iVBsO3WK9h+9ZCPE6hiXFcdy/GDuxa2lhRuZv+DCuc/AmVtYyelVnxscypwwT9JaNr9Ox9
7OtMqhQ38hk66JwEJq4Cg0U03Y78JCBGWyGM6NTDWtHx1L+pQI4GeeaWo3ads9IFELTXtqO3hWAv
BVWyO111z2aSLM/edbhC44CkWBiUv2OZfW9w6K5HfNqIQn6x8wU7YkZ5PFJAX2SNsVk9Ui9wEeRF
sEsJ7d32TmRtpOo7ibBeutn422gxz8TRj/we4lLjX0bhaEu5KxdymhVrjYlcbnSBGVHKmxxdQ2FL
eGT0qFinJhSXGeGGztVMJ5JkJQEXoWfvEObfFyA9f9dNbLorcLIgwbJmqvWT55uLhyXo0uQBbTxQ
g8mWaaAeeWhLyfnH4LOEnabm9f4oMjRzdBsiyO1zZbY1da0vFxeVeV2zME7pydx9Ou2TSQks+B1V
0h6et+NIVTDdNKwJFo9ySixt9hmy4szpE6OeegcdgagG3la1qndzjN2/ElpQfzCsYbKilLtDS6wA
H6hdpp03LkZMzJ28EzwXWZ7WLy4C69LrcNGtJaE/o6HzrKsQtCa3IMtktvV67cKHVMw1vFxa9dxN
Iy6+dI51EZ+bDfrj2HWunAQWGHU4xjiX/ldtZxUbryjhzuixQ8pg9ip3qKf9KJXCRPwee3ndCvF8
MaA1GNeNhmVBnqJfxeqypM5NrYjzvdoZb3K08CGQvG0f6A5VDpFYEabxzJJDu13fqau8O6KSWYPK
lp32geQ/WmTHv1Sx4yAqLdSCJwttfagdP1QXbuUGGcfGHlLlYH7//JvStUW/O0oWa41/Ae2FSQgy
AS52rVoPgZVQ3oqmtuXvKeKwoGNg9k3IhhFmcGtJ+Jgx9RlmTkcLr2YLpc47RcDEY2BNDTaE9bGD
BHuaorpQTKcjAEnHCtmPO5FhaMSwciz9o81YCPcJD+c32Uybb8i+8ZoxNDHaqEO9Y7iSqEcMAb66
a+VuxUFxKiCzk9mEgdAolEe22x4MV+61Oa4i5dn1SBCnIFP1rO4C4p8eR7yTaVNu7s0WV9fLSMAb
GFJn7f/6P62EqHDkmuuLMITx+1CkKiph1WuhlgD525Yh1IRwbCHhEKLt9ULdHKW13LL9aD08NGlf
5GNMb72A6XCOW/bsm65GuIGAfxfi43FRbcxkE7P57Rjl20eiiBqUzTARx9ggP3fcqBrf2Ux2wIIn
5CU4cIvhcqsRA+HI/pu98Jok5+FSdoK2SxXXMBFlrSD6K8UjbdGha9QeCOLhJNoqozAeS/Qc3nJa
KOzoeUvPycDLZfPxe+VDilxX4dkX90ifOh8X5kZ7ExT0jsPg8kpQ05NOO7cD3Tqb5+IW9MHEMWr4
yL4OY9/U1W3R1+QD5d6kntVI9jY5ZinVC/WYTThH35hl/21ghdzqruAefdsPkr6L/7XnHY5MSWP6
K50b6mJJ5/t7j0Po5UP+5RTwQBUUxy5vgeIRgQe1vp444GFIRREzxMh3id5vxntzAFOFBPRaHvgg
oS38AKOU3a3Rvenb+17se1zgft0X4MDNMi3bLljEIrBqQEu1zebmu7FF8X0SNvUJmcf69FQaLPVG
/ruAKWhMdrLiQmB2FA+6BMUY5GTE69mJ0196CGwcXUzzf2CgNbPDGI6i9J4V3+MH5+17Y8KiDHRe
sNPApd7D4uF4zv1RGbpqk3fkDY6k8li6ZZcHh8Z1GLqYBQn67LkESsVFxYVqF0FhjBDsTjxFPVH9
n1A9W1CJI6nBrEqR39cAiBnlc8GDOMJMJgvNnTQYRzOrjyc6JI/28FXXcogF4VaZJlZU19kKjoYF
kphl06P/caUaClr8fyPqk34zCni/smpmKx2rPp9HvVgOclWfbEnnNj2flB/xS5a+KjTSb5aS+jfo
yEZWv8F2mBoN9A8hVHxVUieXOp5Rk7AZzqvB2WvaykG1z4OFXduyVXZCsfRwRIqgeZlpizjB2Cn4
pbIYLLxfFaDnKe2GZT/FiV4LeYRQZ5wupHgfIIMBGkWq1NaxhsdbO2XmMxaQJcR+o17bqy/ktvVa
wy2w92fURRNqApNs0WgBNc2lrhTa2LF+/Cdxe2FInzPhYZYq1Rpb2OUxVTUv7jGF6mTvLBZjDD7j
ZNdb7zoWcBMYcBHOqY+QpvM8kZXglITKjV4q7pm5dKi+y8eH+3XaN8k7faDfrGKCRORSO3XcfFf/
mTpZFok07AIW5BA1ze+WKVqo6r91gJiVFbaD/Uw8bLfPO096KFvHSIQh36/qf/qQ6xVuEqHCueOV
5kgx9XNxZ51pthXK0nYw9N7rSB87UxSxVM1c45Z6yXyDYki9VV+H6SzCH1AAtUxAAOnIfpWg8SYg
0piR1r/ccwM9Nfrytn6zo5KoE3/FxlIGn6k8zluAfr5XJsdszXqH1WA8Z+xI5gZnRl8olHLgXjgI
BeaGWUayD6j9ZxCtrEgVVCCylLfrqGY5tI8V6aobr9VDiLdPFpdfnNCI+SiLOCi1LdTNy30j71zj
OJiqgRUoYZDbnP0z/1T6Lf5XpfbSNtd8L3Paz4h0lhy6pZGebcTL4Bh+Y+XvDLLi1lvfozuuTV+J
/zqVaf/um3WhfzAxwKZEAIrtclIiZdo5MoYxZSlI2cfBpwv/SdRf712FOsi2v3Rr5n9gtt/bJyZU
99XTSX8ZMmYopRBvmGBqJseggbrAj0VMI38Gr3RF04xR/wE9RKVaSeUal8reB+ViS/gsHxjbhp3q
93j9Gd8gbx15aQpX/ML0HJoTIKmll0ZkZ9OOinyXT2+nnHnle3GDs7oGotDJFJQrYZ9jUyK2D51R
qK1xb1EzJoDgqO5I5U17nsTrN7Xnty0VBTHWhvxO8ahn5hKKWFKYkx13TvGkWxeR93xQ9T1vmBby
mQh+hbEdkmKqqO/m/2YpZwR1tjyFieSlvYZTltAtQGXuWQv4xwSwXfVRH2xcts/qsQzTJ+5LQxgv
mHQQUkvXrlm7M9IVQLHBT3DiOCfVZX1rI+6qdKtXc4JcDJzqdXl9ClZNcvn32cTvAX+UtgsjPs+c
EYIvvA4RKHsGOstLfzM2bmWvN9N5DpsVCFRQ/WxOwUF1yFlguUTi91C4SWwLUj1VGQTD3tivzrHd
tOUiwtjYEM+MpAG05+YvaZcZ2cjGUF/GY0o54tsvDd5NjtJRK0t8HAcKIqSdpF3E7xb+CICxPwSI
VaAwhoiY1Hv759hQZZYxs0vLb0ON2TSMk+Hik8TOr01T+brx1c7BdmhduV9dkki/X0A+77clYd4z
PTXheuOgOFXwBycWiVDLZ26OLhuHJcFhDGjP4aHEcv5KAcquCXmEkrP9NsaahRgxjRCaT8wAj53b
/xic0u86ej0BdiMJr4I56a1AYc34zWPOs2GReCV5wS6VJcuRvmHV8CfNvJK7yKStPX+TFxkDJk+r
hcAdBHnq5D0zxLFOUNN9J9SbP80vBzbbSW/sTodpD3rkZAvRVDMwYzZl95YufMeZqWtOU8VjT2ug
2ilOMNoAXwm1FMdN0BPLI7Fst38S1x1lv3Sekfd/jeSVRV5qKSUueXt7Twf5vIOUHSgLLfzbqTcc
mEkK7MODwqXcGEkpWydEVMGyTEOpFaeSi8PpcjJCARkgbQNnS2C3auxPjW6ZRD7ItV6sl9Fm6gdh
lks7WxuMnb4bCvY/K0pCQe1cAAwmVhBLxXdREBJMHV0JSTuVJiX6Wu18/lhpZ1W6UhJCS+CAq3ne
xWwvgDEXiQTFG7CSAn+rModkV+QltdUuXS2gjSxxvi4fwud+VkKHlJvrHZeitb9A5Z1za32SIT/6
h/8o9SWlrDTZgmjVd8Zl1oeFBP2NuqsxOaQdE65/xfMWvnyh1cxMGWU0g775nBpDvyA7VhfSifyp
CPyJdXeRAeFeetoWPg/F8wTq0jYQ5TsWvbTt3J2/W7ylWqTtleAN3cSgRJ1B+XIsFqlQhq2Fd5dq
s2XdlGjDwwqlFCydxai0N51LJFlNBdkl0ASRngeUqBA+0YrsRNdG6e0cq6zrFyfNa5TrJUTOcAXk
JwqHopIga/XnWs23FDX4qyUThNQ1uLH4ucbJMducYcOKmsLYir59KdyhQLclMCkMnKsOivUDTiHY
5pFVbCpQz5G3W4KtziZFIwQAEyoTSE695WwA5SGgcnmCnuuT3eoOf65fDRrhPcZEPH6sNO3Edc7V
WugIjAYZz0N9UHcW/cydnfH0p7oyCrftAzLtBU7dwawPa4+yCVCRbtTqj0hOPwagsomHracrB4c5
SPZbfnQyRjeN0aO7n2/hG/wiHcFKqxs3zZngCyAgFsLuBRiaLJg10GDgLWiGPHYbuGsbEJmOdkw8
6kUHzdN7xm0DRiYN+7alN5MlB1zM06voZdDSYjfq3BaCa1i2waJrE3k3CGD4NWmgeUCzFIaAwlrH
B3HIhs6kjE9BCWF3ci2rH+5XS+6BmhrvD/BeMgZPRGcpmvRFZDEyCfnQSS0pMwshJ8Es7DC6TKyo
doEUZamnZRbWH0wwytIqCjVC8vKIgE02zuZPt0GY3X1aPfbaeuFsHZmfm9rAsyNAxtJP6PoIu/ph
Ez6UPTq/0FbHl7tshH8eflmfhDdKf7GghI0mr0MfI3/oM7n0sTwAi+Hj+oC0RX9a8Xp2Sd3J0654
heUENrnf4ffrRO/2hYhRBPqfbRlxxu3Vz+XS6QMxrXVtePSY+HyKYK2QfEi2sDZZ9YOPlbknLZ6j
hxVqCe+9GbccTFETJy2LPQBgGBfxpXE4xhk/xk5OYDNxJmf0YjT2Rf/vZm+kiqvSHl1peDGJ9eHA
BjoerYip25AHaWhHFjf+C+lPArAAVZo09viy5O/IZonDe/klq8vuONqrBLgHPAHBK3OaZ/yQZjdV
CI0oW/Obw/v+AJIrPXk/Wfytcs08hde6gMnurWOb+hxne4AjPYxsNc5PQPMm0kSNclQtc3UZU0XO
vSn6PZKrcNdAqKhhlvtIltAef1/lpf6/msDHglx4jfE5xIo2t2hEsJAMQW+3Gy1koGKo1GA6ET0I
tfnNlocP2rzcZVuLgmdHrp2k5HduD5WIz46eyJFpgGZ4gQJj10Ms815r1cJzkz48BoX2xpQ3vQGD
9+v3bu79PtalbCrtJhtDjB+695Phbq5meYEZL+GQDQo/EnMr/Ay21ou5Y8PRd+85StZ6k+9V2nAh
fCvK8lrB8akIWOiI0cBHj86UWGsj/f/2S0mQOT8s6GtkYcDwNYm5fbC7iLXkm++LTs21dkEGmkjv
aZWCBz49TQXWW7OrVXEJyfrf3Kp7Yu6exl3rGlPd5ONGqjRuScxhrjF7AL18soKQ6bOqdK46Y38F
7A5UDBlOvwA3M86kVFypLspPhgNnJtoCSWkUIwtIjWgGhlra6XMFF1RvtTZKR+pEAY7wz/gH3iZp
XYaGe9TvebppQjwUYOlw/KxueZ6mOrxQdTGiXzFHAjEtfyPH/XdGrhN1gHyKIGt0JtbI5ceCzegC
+FL6iANg3Dm5ctLuxwORxmFrt70kPLmJ13w+KH+XuNaT6zqnIu2Iknifd2WO9BgD2kl3aAm3Dwju
pYSarL2J5qGnXnXFFF3ZdNjYwXFS3HVQbxgyZjLTdJP3irvJnbOaQQQ0HM5s/StpzOhq7TZPNMQp
VHR8aI1sIcCmDmNljzpLV6kqTop89/VEgkNz0bBoH4bXC/vKUDJVPUAxalCu5kj8A3XeX2AWcKPA
d9aZt5tBHojXw9pG4FfPhZ9Nqt4mDLR5vMXcqTD24YFcKdDZSP/NP8gq1Qc8Idqq1RsOF5oJOBu1
RGSX4HpDsu9fY4KT8bQwnEF4slmEbe4vm8HIBVOnVvASD8Fhnb9sQd0NnYmAVCDnCBtqNvBT+qAM
EeTbKEOs9AB6dF5b/6Ymg1Kt8RTbIcUkALppejCac3S7jOHQjibPY0PFCrt7IhVL0ZEozVcriSUB
kAMFRbLTVm78lFGu3YFNOpBZMjDfbJBxsc1y0WqqcjBm5nxYlP7KqOhJdXW0Uqrc4eOKAuADW1lU
y6APtGUMPriS+6PKQqqRKKVPJJs+iCGX6wyJHWDiMr2riXaSinTHh6RNGaxFG+fjwtxe1/DBXEU+
LjGSulw+E2uccFr/IWy9RepjG5UiZfF0b/ZrliSot5gjVjOtM1yThjwynJby71LOniSOK0p7OWbg
cvjaXdd8ADXDVWZ1eF/mZwxYObnYhGhMReBuY7ggkNJeSV2muBCs+2MGpH16h428rJtD0j8va/gQ
XHO8ctO3vY/cjSuKHJRFc4HaWq6GObKTmlVTQwc5UvZXOmSwrSH2IgGbuo8tcgWvI+5XHsP6+FqN
ZfLRomD6VkU3jh9sdxm41a/qQW8vz3Rzy4l3uInZ0wC50huijD+46hSZS8uLcHuu53xaMHeunllW
GqcfFOErngwgnrUkBvprbzhbUF31x6U//BfmIIUn4Hywelu4HHcGjPfmS1D0v763CBMCkSVpM4xM
3DrwoKzd+dYe9TfZ3pWGJN2HYvRdLVJTLhmhjP6+QhHCWDHRNtRfRYBhpcVkUJMtUmFx/aw8CQXa
wtQHM+2XRChtW9wh7BA4/HHnjB0oV6sfJIKw4pPOteemDnXUhrD3TDa0me7ZM+yT4Fy+CcJ9zQvW
8lxQogqF8dVRYGRFTZH8s3+dg66D/iEpPS7Cj4hhMwoR/+2HfYBWg27JxsohfUeKUTHyO6P07Mt7
4F4UM2yypI8jrb/j5jFAUquZ/lt0vZduKhdliMHJJUeq966Cmi5LO922reSgu77n8m5gch+oG/oJ
agwaAUhCm1StKSESk3VMt1ByI+EpfgAXm0haeLbT4vn+BuYBPB5EuvWbq5eQ4UIk5U4Vnjno+nbN
IbR6r5HGGdkcPi77BTDBcjDI2ptNXllrgqc9sCi2I1dsa2SLOWG23VTLRhuQfVE1i3ZH9oL8cfDp
SATDQJZDBCF8nfJPRwVQn8EYS95dP4kZb72Ck/7exi5Yodoe3Q3wi+3LuRqvR4QNE+B93eLTmC6G
8wPcv6cbmaq9CWz93cFWSEUj+y8LOwWsR3+ge7Fb2vO7zT2aHcg5oUYakRVW8eXoog3ABn75dk/Z
VMNWWU1S2NJW2PqIyUXbobydhrSRjdE3bkp3tXtBoNE4R60ybQnaIQwupqVpltU9L0vmA1gFxJ94
yDZsOfoMa3f6fYQTh8IPHeJVja9WUsCwzyK4q20PFdoVDoOLs8Cn7LIPNVHbvd+KDD+5kzatVvpT
tXjrfE771wz1VqqXa18+uvH8YZE7tSQFxA0HAqYiI2G5hFPXenP1saRp/gV+TXcgqaR4xYQpLixs
XYVFLgjWVHBMeTMcH1r56qewzY5ww+Y7FtS2wknBxXia+m1tITEdiRMQQNMTMKaEbC/tB65ADst9
Py2bZvQojbJI0AWAy2yTuk/m06v9krEqMVnYltRbHmxo3AKh3CKgBnh8qweLUNoiES7vcdv8VGvq
C9LkRlIvIxrL6TJ6TrGFccg3ncB3vwRK9Ka2rLbnJFQUS87oZX+zH6kTT3n1ui+MF2AfVu9+jsxP
W0eR/b3iT0fyUpjaIM1WHwFW4K669nA5+cSenxonHrlyNotff/d+E51nFam+stD/lMy2azn3ghHc
XetQ0ASKolNOtuFaXux5YTp1/p4T6+FlXB7ZdYXPMEBUFptRvMN2us9746jQ5aqCRT0vlwsODg2T
Kdfb4MlxfUtCdhmdCttaqW80mRA9CgfkXjwfsbgIxBu0KPH7O4GjF815oA4iIqKKjx5slhTfsLHC
nLb7Yo5cucHsM0qZBQzdA2pgTu3kdZrwAcaQxa73w2lpSTegFByYD6GWNAuK3Lx41FialN39rmnP
Xdt1MuYIKXVUYvaVV3g1tM0k/T8dcRfq/u4rMexv0Hsj7GIbRSxR3yfUSktyWTsn4AhHCNpw/Bme
SJgK5deZ7bekc4LA3NGpx4lvGyWlOESMnZfJm0MF9Pod33RxcErXXjDl481D/LTrtnSY/Hwmlq3k
dVQi4sOfZxqAmsHA551zAkk/5Iuau4mSyPVJcblpV9iLRBeQx5/zQv4ApQTNw8JZBeCmdn3Vm0cj
CPmheRG0k1zuvrVi6R+DlUcjDItZ2aFKhuY0sfAXq3kR3t34Rb9w/gDEVzVZfebqBeXAFSxZF47A
8QErgyit/bAkLDJBD4Z1rq9TnIOFG46G4h1PBOv6eK98IPV6VA0zpocjPSwLlQGfzkm05RHwWnTx
Nmk11P+13pYU/aNjzGnB8YFk6G7BQOcvsvaACzcSjG8gIYI8mzlG6ymqnY9Y3eOpLRPP4x97oj7C
lx6/C3RNrYIYAhnBpV7xeD7Yv6/nU7KLTEfG5+OHtdKHBsufa7Z9mTFX2o/BlKZKPUYydhD3ByqU
DNHoW4D4G8HCYgS7vtSSc6P/uDEQMu/MTLVJEPPQOO3y3oCySBUUOoFGACTo2LOWLz65hfyIqDUg
E/g3mcnINGVSCiGwXFj6GI4WhnVxeh7d5hl4tFn3t5hbzml3evqICHaInK4DomsNa3Topw6OF4Hn
KairVWZ4ZVfTSmEJc5zZ8lCVW7R1Nr/PDtdwylDXjPuOEP4Dsp+91jk6nDsBvUl2RdBRF7SVR8jc
hnQQYu9B+s4wp3Q/4Coo8Hi3LjntATlbud2VUFReCczB6A6y1ny745sO+JVfrxEJBftJ28+R5whV
9Vny1UHRr6OhAUBmU2WU/mJ4MIgkdkPVnW8VID7T6FcvWeDwo+g5EQRFc5E2O3dIg8fD+SNRu7z7
7J8IWcjiC/HE55UcWwjyHaR2rjl1E5uH7tsH+6p4MYcCfdV7lI1bEftqfQJPPkfwSU5vR6M1TdNM
ROTEBmvkCBocaOjUbVoaAs4+UOPwPAclzZMwhOaN4WshmZmfSRngbgIUGPWF+n4IXLZp4lS2O9W1
G7LX97wxI2rc2uKUzd8kNu21AFxTXtuoMSZCMJVA6CjM9ZwLBWfrYC7HdW312C2HgeArARh6DAt5
ilgifa/Zw0EZborik9zLuujYSDsf3SR095JFj/nVllOMMIT0/mCJEAf4ZNtxOUYDsiBTGIBqEHXy
XTnAmTpgTpi0q7CRIHgXeTmYTmPugF6R/E2nPEs6vEkIN3ERwZNqKE7N7rMwrnVxHeiv3qf1iDhh
SGY/34E1BPaePyGTWxz/fioY5caZmkTGGfHgfcIGnvboc+adbmhXfEdJPUgAVIqURU8nFis4hJlP
qdRkd6kPmyK3kCfVfVx9WhOsoZiXemjQG8l6lqun/4qtgkhuDITvZBvU5SXat/AEpbgNA5EZwcuF
umW//TvCTtrS6EVfJuXtXatacrBmwd0QDwIHyu5m+Vdlilud+Z/u3vFKnGvPm/bLU2IfwlBbmZRp
rRAqtqDTPzMKDQA5TrSL2RQj4HjuNsVFUpfhMwYpcJTRfLlbwWMGvlmjBarQv2XPMOe8yzMzBQB9
oN/BFnz3YzU0Y5EgMF47j6wgO2xbOTlqfvHpC7U3wmBgkP4JLWZkTWae4HtJ3ROaPRtR6k9PDdJZ
WrpOSrAqzDi49VCTQIVJsH134pB2bwixqQmxCGvaNVmgVPgU96mwBNHBKR91SNecky8sd/6tYCUg
XxrtAZk40IQC+69pN0XJ/p5b43lxTRLmtonz2TvFaRYmePpTdMmQPnRnT+4oPk6BjBxmktxpiebn
e4YlBRrag2qZ60C7DIFc9M15JLnLxNalG0OsL6MBUXpUk71unlXnrA8hglRsc0cfCAr5EPEBJZDk
x2BNpHxT90Z9n5d59EMxeBA0AY7t+sKpjtd0dHWsw9+Dkksuytacc8EDnEAKsYvnJhU+pcvV5reK
Ov6qfSOkDjz/a/c02RaXetS/s2+FwkgfB/GtuPFmXYZ/7317ITAtUo6cECtF9Vl8FT1ER7VCcQQ5
kWYLM6cuFF2zH1Z2emQt2XoWTwauTJP1Pq9/nSX1pzuOUj+qYyXAk9ezhAEpb0FDLgdUGy06XNmT
3scHemY2yO1XVpZaLldhhe9y4LsZGyC6YomasPdwpPEX6QQmHThmBGa9fUtOY2/AxhNhPo7Dybby
2pvlgT2xBBUyjpWZ27t7axGRju1WE2C36/6OaP206Dvu5TilVxsmkIvVBjSZFqTEn8ItJVhgNWXS
BxwVRXnfyJ8JEvUYEVMJrfekw9y/81lSWOUozaf2SAEG3wrVaMD+jhJwLwst6b0QSCk5DWNxs0Y+
5jIgTKvp8Iax1I4vSNV+qjo6xIcKZsjsSmPCWMiCqiWmFq0D0cG76g4j8oVhxYXJNuEhWogvT7Aj
xFJrY1wjZm0MHtT0YaXM+1/8QeJ2k+Db7JVOK/YzmlA1/9N2xM9ihMQBElV3nHqEzqtDAbzA+Dqd
j2VojOn6oiR9wS3NTI/9Znl1wlDc/6/JEFWSuYWvwuEl1A3RaC9oQYAaqOeiJifqferh/YHXzRmw
MfU0j+ivIhYkWl8s9l7O6FlO7IcDUJmZ4W8ZixdUj3mb0tvkF0Bpi6Wy/pFesuNn8rc0MTwUxLFr
X7wckUu5Wa/0AyT85bHWoAZY4hzfC35MnuYKZTcsrjkVKVebg7xPG7im0Fibil2Y9CA2zMpP77Ci
/xjgG+BR4+BNEzGZ2X/8TGE/IppNa0jY8NA3aWZ9OoTou7lgSM6Dro5PjOWTEgzreMc7xK1pVr6u
P7qvm68CFmiwKjz1aZ9jebyC7ieIccpoXnWIMECsXFgE2T3yFTTniV0y6xKMqnjTVvJnaKKmcw/9
9niXFcF5XheDGxuusrIunBXwiePN9BqhwG/MdsHaxx1WY33TjO8fnGQ2lube4pm09Wk3fb/TvuS+
blB1PQ5Lu3Ym0Mqf//YxpOiMDm2ZucixMemKN0upn64NjVrCpEVV1MH2djBRjr+qk8GoWo6X7E9x
2SrrYc0xM8ZfkQ/BEZ6/bLO+IdbK4n+YcwkgwO0tENoDeW9HKKfzva2YkXek5ggHypuF5HEjwM0m
uDD+sE0BO8Nt6nkHJsWICt9z0LrPqe+okEcnOhvY7ys5FADDTxfLQDlSdFc5lpNFwgF8LZpDZgjn
0OwmUC5N+bm+fj44yUoqk0YRpQKH+mc8R+fGvpPEc00gHnoaKII+HlqcvkGyvWzTMpuJzE3LallU
5VhUYPHH7Ue/cjmEZ4P+jVE1NYj7P7FEgh7ysRy7U1KVfMJ7bRBTNuHIQDEqTO32FqvTvIeUK02L
uV2wRjoeINUYWNxZ7E5BtqQmqf59BkD7ssbX18s+S/ZpXHugKj9TdS1ur51PWuqWhyaks/YaroJ8
sflIg+4EWRWLgWifSY0MnaVt1Nwq3dTiiD2KLgq19Y5FrhUnqcJ6i4WxQ7kQ9fMX9bHY3K9OHUoJ
HqAU51BSL5CHUtoMqxQO0kBPXmIGULT+tSVAu9UcKuyFkCvUud14JhlzZfe4sbGLD5I0K6Z7K63P
rZEujTdBZWLvTOiXM84gzcPhR0yvP/b/dgq0mVuzNMgPDBtNZQGZMKFUatvYwAj/IdDLlPR0fYO4
1BGKLJ3WdcVhfo795IQNtOadpMbjiqiFr9x2xq91E04cGjdNQYzLNAUeXf8xzqFv59Gw5Os0aCh4
GwQoyhyuC++kVlwknzZwOJkFb+nJx9zl5cMgYDtAYBnzq1UoghU8xF490nX5oLTnbiWtL08ku1qY
LDbUi/Uejzfu7sWCfilq0JiV5dGWUurH6/ENRKyR/KaQQ5KvIKVOWXVzaivgAS3Xi8alS4jEo03P
wNPHFF6f4Z4UWEfNtGepwJ0Juz/3oVdOiUjRTmbBWSLNEXVlNCB9Yjz2zka7A5mzHyvJPn7TyMhY
AoOUzM+lsNWuv3wM4RnTm1ULlwv3B2p+QAul9VlnoVq2W4rBfgxuRCldusbToXURqy6siFxfsmMO
THReILmTMqrCpW9otGAY3OeQ4o2kiart51hhFhuh0X85sySKXJJihL9PY2Sn04+yQBHlLXoOanbH
2jpQ7nl7jJ5vlTsV0EFg7DExXOrfcAyvNBDm0mDkOu+yAbkzfNlMrsVbRkfKXwIIHWH6zFdpWYJZ
EqLeiBm+Kl+7A9fY/Aog+1qX9U2TIaXhfo2PZDMqM0xWsxR4f2rIKJR3XsRvRekws9qAicqn2YWs
BboiIfpayj/0AvyG72FMSlno12Ib47Z2P/soRZhOHMOx88pp8AH9Tcxpx3vI40r6FjdDeCCNVhCP
iz9LII/0Gk23lc06xgkKGZZfAPtnh4ESqXb+A81k93RL7jNQoF0gNKQblwUe3ct1KbCSiCw0Ii+x
TQlntVBRcL/T+h9ElVrQHyzMCX8uvtH6bQZ99TWkxb+1W6O90rqazJrHAQhn9c++TuNsyzwMm1qJ
MPP1HCMcOy04+LFShxrj6U9PqPZhhpfXebPsZeuAjPm0kBQYHlHBI2dgi0G6ODDmjIw7caDP6uvA
8I4Di5F9VEcN3lc+UI3rUa4qcktDbu7KPUc9UqfBpvlDB9hkC04RZuy8UL5+0gNLZA5dNdTBHGVk
wBxaJ5ftgF/67f9o1umTH1Cl272GZqVrCzRZiu18iOEb7+PKhckSJEBx1SAT391ao3IiO5wq2JVj
XTmRK4UzoK5E6iMMeFVxR3MH0a1KMTcspGuMpKsedyEHxuC83gB3uo4C1WcOyqbPtlzLePe1hJAz
AcM7PrsNFBcNuBoPTy+zEUkguvs48qfZ/gF8r6IY5nZXVQ75FnK1a5Uniy3Qhi6u5J9t2unFB8kf
3H4PQQpp1c3+FOzrxH61DOA9UwxRa7Du1iC6r5JWneZH+1y7Dyg/E+ffdUdospFjiNc6rYZoXEh6
PasJdKN6+3w17XpZQ6VnWUsnB6Q7UJYWlfzGGfkefLQawR3SV2bQVLQ2Eu1NIe/+3Fv7htqe+uDI
pyCngJZ9b62N6zqWY1aAFqU+lIhgY3NYO2xnxYZ5NitKHjTHTaeyvGOrAjSFQ+F/4Arb/GmcTRz5
ENPS2xgU8rCLLXRG4ii7UpHaTETzrx8sf+ewk2vGAsJUUlJCEi7rn8AdNzjzQBQn2IrSWfEMSNQ3
AqpghkcW+qM1ULPCaAb8QOD7Dv7pvl8Skrvs1VvzVV7nxR07RQuiUnGGIK++c2ztzBnEbJlqb1cR
Te5/5wJiPpICb1mqFnIhaIyuA07xupv0I8lL1404dbrrcauD7WLsyE01jqs97/ORzjHmZScWCFDl
xH9LxDTnzVwJjSiTWiRCtEvGZFv/8yc1MkDaYavD7bC5vgDyy+06sukmaV0qp5ikMU+4PKU1WK7O
ldwJou3JQYgNi/MAvTvMeckQnGB4sm/ouKX16Nlwh0+GFGdEdNvBXaTY3oYBhQD8EiVmhW948ReS
kugjUhMg5e5jz40vfBXi0fGtn6WBhHB5qrXzYbeME5JM0vXDuKu/ocNk/arl+6tfghE8JMgmjYcj
RDKpUayFVqFmBKYGBXQUEQlnzdLcZLOqwQIcUYdepFqFRSbEeZbOPHy4U3ADv0+/hI0Ll+Nc8tPz
Zjh4+ADmvjo8mrxwf4YyyOwik9epnpK33dOEyO1kgQ4+6Pk5i0YoE/qpyx/lYD+ZyOber5JX/gRo
JQaIdyzYo5VOtpIgtt4hdpYs8rR90TSqW1ubCkMX3kTkBkXWuPWy2aeVq7a3bvgPsBf+bgdy3sDh
qFDXGF4GvbYiku115rBsuVm9ul8Y47uDFIQDvlIwpPvYQAfwR1Kg9YQpjiwoluGAZW8l4ByiqCCb
7OGm+32Q8ffz0BKXw/SNsFT+CMgqyhOGLZlDwPhhg8C9bQrGQOymD0z3t7J+03BZfAdeQT/Ji6nY
IvHEKdM8XDGGsDOeZZaumDh0KaKFuQ6APASfwr6YEN93DwhENOYGx7EWO8sONHOZJ4xJwELxCFIF
hym4pmAN42gnGJYKrNO2TIZbYU5wLZawetoiZNH7ZNudwghBgvNRKrxREgMN5jwqz6ZCUKY3gqBG
5ofko8aOZCGUTYZ3jbpxUBG7iR4q3sBqrcYzQBd4OnivjIo3gcvVBSBK7wa0MTzGX+uJ+ShyQWmJ
kgfFDsP5vGzUC1dMxE8dmK2wpVNhpDuuP7H5o337cuG8LtSwoQVrhSZCy64dKMkArLPokXeeBGC9
5T6vYb/am5XFpsMDC0uBNgbbQJB53QMayDiS2KHK9d0hyKCsXuTj8qayk2MO4qSOyZgdVxSlUA64
/vh7OXtPh0vVd+drmcyXPEPm6sbF16jQeYrqv6gh/nNcGbsanIiJNIRm4gkHH6Xo2RvywkNtK02O
9tHZ1gLp+tILoZ0HD7WGtxQ/XpOPbVHUfaPI3hYXJG7tlqDfEtjtzV085jNJIbCDecZ6uj+LD0Dm
16SsLd2LZ6bRvhcuiV4byGjj3aVFGenYwiKXzr/QvHhTXc5/SN9g5tv2MZ4fcUWvE8m+Wdcvrq84
/UrubxzyVgyx8Dpv9zEZ4QeqMtdL4Q3maN63MJucS7sv0SIwZeOtATJLNkgHbh/WmV7HjO5fMOur
D80ib68EJ+/dX35T6ipiMbqD0E4/AZ3FqhcxtuvmLnIo+uMDQcy7AM9nve1Kb3yEgE/u0T0wtYmx
WMHowD5etvm+zQwJvZCDCX6adx8S2YDgg/oxlwQHfcXPu8bGI+a0NLHmX3ab0kjLXaUF0uQry2Zn
O+4QXk2ckqY4qppcMMgm9om39nbB1dLzxuOr0dMnm1rBEzEPZTCu17UjsVvT/nT5pQ/QpGCTGPw7
rtHeiT7/nPzWyXwbKkWx3fVOtxDKukjrlJzKYiy/df3RU8S7YTi6Io0FVaY0JH7SvTws6fbNp8gu
JLkMUJu0e+97HdLrSKbeto1SPwBlu2ZLd0rT6sIUBI3CzMjHuhB6Vg+MUrpqefsA6ErnSAQp7vpA
u55owgPuUGNZ9oxgQKajhEuJW6zmD2KLTzdfX9Ap8j9EAtyBVe6i8q9GbFekh2AGWkQ/iLm4hCAo
GavRbWX7tbeChM6TwcKiH+X9VpMK6Lq6r5dGo1ReIxYB4Ncps9rUKbASFS39UuywQDyObJyO7ll1
xTOrgOaUb+zDCYzuJxroq0G4yt6Dki37LI/XyuUxe7z/NbsavfO/TxchPRuNh8MXP0o3wC6XUZ2G
lVp+U3gFhs8DoMp/OrqNHhxVeEHc5QWzyA7F5JZmPYK1Z7JMbXTgZg8kekxvLxuxWdNwWTN0DFhP
ZQTZ7vtyXoujAhte231tGHVxzuazsAcAJe+7MMgriacm9ifZPKWlJY28QtniaV+UDaY+5mem0V/P
LFTsYYbSUkq+ErjQeYU0UNftMHZxwxlRJoey6oP/IDBkL0V8KAZU2KPMlT/SuUtNBrHIQ+eV1A58
1Qz4intcVh4mC8UJ953Qpi8+udr6IUeahp4Ns3XeTz2ZuVqqKSwnSZICtMj9kc2XoIkJNqJT2q6c
HVkox5phXkp0LTC7kxwXC2Rd+czU3RS4NpApkxa3X6wtMkbcNlkKvincWPO2A+RZpdGFaNFJHUXo
SPkmOYfy7L22xQNfEflWTkhbknyY1pqCSck/ygOeTd4riMrLQMfhT6zWi/tTj83AnrNTSp+7XOPJ
U4kN8a2NZnn640HOXLjBO5T8UIq2y3M0ShUiejni6P5KX0U+VNAOE6QZreqlN4SeBWn2ZtwD/coq
aS1KCJYWOd0A9/R1aIDmq6baFDKckeOmWrjpD3XxOgTU6GVTXcy2od/4zijqNQe6ksD9P5lyiVoX
uUnD0zzUweLDLd2mHeX5yrKGsGhoURVCZWhkTJ907GQTLEPXCLNHixJFyzTkTs49x8QYqeK7KB8L
lN8pYdDF4Hezi7rhHtW2IJLwk4KKZP3anEUF1muRBJJGBmUc5UynKRXRe5HR+gih/l7KdSzWk2KM
btmVCP2KUp4XHEKhdzpJ5PJqyIWjrahIKsOYCpYa8KvmZBRG8qGs03/25IbGHsb52hlvI/E4iHQL
ORXstnUAVImza16fap2LQEOa24m/490vhqUWG8W5rWyEchflQXzIwanlEAaJPH6UrpFCMRZOAVhY
Xw2fSe1WkeIj0XpVNzuKyi5fsDKEyiB1WzRcPjodM4qGI6tfdZ5xsEUuuJMTF4YyqJKs5hR0pFha
+zVbjvTZVaq2rkuyCpzOqJoknTMMT/Rr6i3+ZVbS+zbENIerx0Y88TXhhsfhpjeRpMI+Q3H9gRvk
5CmcEySX5RVYCc5IKUvvV2ojsr/rgyygeR7FuTDKr+v5lCbldyVIApNNLi1i+E9geUHbpvXzkhZ8
DSEBRjyKdMULqF7+zTuENZsvaO+kWY6EDwlElPZrFE0Du0QAtDIfV8N1JiQTFJoD6133dGAioah3
Ys395iyS22uDjb51iyhrKNvu7R3ePty+ydIU7k4/ETYNwyMqX8lbzin9mgPKkjlNXl68R5uFqwuH
hEvI9eFZNjyePJPV2q9wSozYs9h3IOPaXI9Cf89AaFggUkWnv1Ty/keFGL0GdiRUy/q+a6dOgZzK
9yemqL8y/jwvzANL+9Sq1meOWLvqAjrHTSxeoAY4vXgtayofU8cXtQtYusJuPQUKfWpdsp+lGFXV
B6UASmgqYBcNozS7f5e9LTXzmrrI4bGnQ5ckemGnq2cCa0NsXXsYNRV7wtnI16t6YfgA6dt1Oe4J
RBbE2XfO/aP+mODYRdoklxWTJ7plk81DFw0oOcIJD0XRsYhd0yXPXg+feovjtwWF9bEEX8dp4zCw
KJ37lvxUwGtfPrM4X7eG/AF7pqfo672iVTZcxHqXj1ZJ8qtzmesLkKf6S2K15gNbWmn8KfSwMK2n
jJyNvNWefJFq4tyLUyyGzoJ+LnXouLx7byNcITlD5UuXGz/Gkk/uh2piTb2UDTJLHNidou1T0woq
n82Biy6tUU2UykmfxozPA+qGeR72GxjTpnuuts0eoQ8Q20zkK5kYHntUSF8TBtX0lAa/IU3TsaId
zq5owzXnPtuGq5maTyvADNYH6hiL/UPLmWFvnTCJOoXGiBbP8p2pws+BI1V8IjpGSd2RW58+v4i7
gwkDzpXdWGCaSk5wzngsf91GiEUwMWSYT5Y+9+kJo2oMjN/YCP8C6TiG67oPxYA9JNsFWwaYvCEg
0bnIUl0BKTO8q13NNgTN1PadR6M9rDX0BzIx5v1gaAOr70LsQoy3ucm+G2eVQICa/DiPH6+6k921
JQvrB9esDh6Oo1BDkSmqBVYJHz6wVPvDSeMJcbtcYY62Yt3SY6KgDJF0eTEUkr4LZFy5jeJo+D/M
bIOQefYbFWTiWfUkm7p19mG18abhOxDZ/P/IqlNuzbTBdmfdJ1XDO2pk5skg+e/6ejeenMRZPP/p
okoWRW5/qmag+Wn26w3JgFFz1RHqk79FY2zcPYmJPHzaS+jWSTyKner9li4KNfF+hGfF7aJTIhEv
BqHpeWyz5/wBhsZBa6l4DZnVraSbXGBS/YhTz1t5vC+S/O9EkT8c/mmNJAbXV2GnqolJtmbqFZni
WQb3CyZ7CvIcYz4SEHCc0tObD9Y4Z0jG4Xg/kqPUI5YUgaMMWE+OJZCCyLQWOfsvooRZNQy+oOAJ
sQ81Y2YIbE/mvYixWvj8ccebWO09QcyUO/DCBIbVqSq+jGhHdcY6iK28LUOmX8vfMpJb5DV4xc0M
pnUnPvdTHyh/C9HIXMp276AxZgGUOvxBHM8b3dg5Ky5KOiFAyDpWOPoBEOKN19iB2nOnZlkvEue5
rysZjpGwPuChzoRVvKKYy1AWQ1nRMNhVo5SKgf1JqKWcgk3VsX2mKouPHtc7XhNe4V5GZvYNQokk
Ns42k4F364frIPslIS0CGoD4jw1NA42P0LJrwr+zgtTrWVt7R9ICX7cmWbL67R0YEv/XcnHBN0TY
ZEa5vHJXHjyrdyB7b+1+ybPv+71kynCOM04EQFsveN9WHM+T43sUOHE3NsTrfRhRzL0zjBzss7/o
N82n4aUGMhphL4XZkEL5vixxAyScdkIxS6pnRiLdcOLDWLDmPx6aGovnNKd0xEN2JNlCGk9Mq7WL
cit2VLwOyHbMTUV3jo8MyvLcz8/s+Ko3ze1tMEGYzcS7mIlo9pz51Td2R2+RqLkoaB0jna4MhjSd
RcxjxINJyLRzchMLaHtyWNdpfFpHkvIP8sRUW6hxQOQZtOQYaV+kmb7CUiDuOQ3e7ddjMyftoBM4
ACytFE9TC97mlFXCeQ8RPWxYCE2MKT8AcFKRBasKNTq5xlpuflFAmRk66qyWkE4eVi7cfpk5vV1S
YhFzNt/mF0at+0h8pFSTdpJ7dFcUMLqUeJCl7thUG3yvux0uIajbrOT38xyd9WnIA9tXSgoZ7PQY
3iPGkSD+KyOBW8W89qVneL4HnrY2Z+aWp60lKN7D8z1tzrwSA11ax+29YhPkiriUc0prPj1JeuY3
cLiOe64qbTlPPC5uKngt150D7m+z9qyZuXDKc6fKCELfqmPgXoOZRnS4JVnbv1H4VTe/B8xWOKe3
KTT5bgRxusagYdv83wll4NPFpCoyidgg+QqaPSQ5bqU0bYkbxEER8rj2J2Om/2ZUCi4Rvr8SudNc
0t+KbXtECfQnUOlSqftqr8T9NE5cwNs/jwSOx/ay41jqWkDvePbqpRhWcfVPsOqZkgPkr1/NPgJW
7nEE05xQFXO3JmWO/Bc6Yy0VGkEhXZvV5o7os1lc1GXH8j3eH7Pr9ws1D/XUambnc94ul615UotD
6Z/eu0fN1RJwscGNSMKq2ztJNmyIQG7FrL+KCjf1fW8Fmk0NE8nBD6yITpEGHHLngURmAPsJnEjd
yLgVpMZ0fzlzS0QcBVLyrIA/RUKXR8IQYJ+YDDQ8mdMRaGVgGvSL+1jA6ofx+8e/4yg7xyyw7uMV
l8WGyKoJ1udgqmBMgKixrwxJ06iUefxETtZee+ZLOSfiGATWkCmm7pjLaaq0YRiqB2OYFlKJV2Qr
TmbdlHsP2aHxjJkTCxRIfzeFOS5jqXq5z3XFo/hWU4PY74Wjg2i4YIGaD4XR683Aa03ak0uMfUbQ
cOmya7bPuhPeHgDW2cEawBzgowtskY02XO+RDgoHeHRG76HftlAD0XhO39i5UYt/bo2BxBeHqjIb
qYTDRTB9NZyG1uE98i1FBScDHP8La3S7z9QNfNY5Zts1uJ1SRwEKrM/Eo/1VG+FHsBlL8/q62QJ8
Q5oNXh4eJBkELyzfnGTTXqQa2BszCQiyFq8Rrddp7gXC2OZPh+zVUVHlLDg0+xm9KjlydaE4pnbE
7y0TmTkde7PLqbwwTQEJqr82uIVchL+FrtyxiBWKU1WOk9ot7IsqVR0M98gcfdwFd5CLMqkG+HXK
UjUJ8VPqt1ye8AVsUg8WpcvR9rrCCfsEv0rncHM+8H+AEbhiNtloghWL4ruDqtikWa1tgmZWsLfj
EFZkZoFN4XvpH/shzHAk+CHXVi3AaUa+NjYxweO6OK5U9YLkcz+mPJch27o64e8FG7va0i+rhA5b
DPNXFe9lxCxoiL2xTle7iYf4ylvRQnjPO5dHHNlTlj45Yy8bx9K7nf/L14npB2R27GjMazpNONaI
EeuJbkNc/oemLYANQmcqN5P2ZLDlqM8XEqS6jFKdzLYWi5eI/hoFKZs1I7eXGtXALro39sn6mVRk
IVwYkVPnRoT1PcmjwkCPcEwoW/v6Uu8B0NXEYpuRi8p67RnX03UeIiHYuhNk/8nbgx5J01w7AdMD
9iEYkBUytU1vjoQ3gTFpxKJ59uv0TsyJSX1V1dwb8g5sjTcvOPslKNos1nq4JNHGTt5I+tz+EmL2
UvnyHDFcgG8eC/Am36buLbWT1REE0kKcJD9Lc2tCpEiCG8rtXUqvZ3IdcMb+f7b5r7OYx/Y1aYm+
otDhOAgLpG/Pq743jm55vzv1Ez98FQAxlEnKWuKbtSC3zglp1voaKA9JvSR7dgqhA+Da0A9SU5iQ
HIlzkBrxbRF7CNqxqESRZ4v2fpFyZduGYAWmh18G5N6dyKg3TuP3GQjHKcx8kqOso1S6bIXhXojX
Pb8617NXL2jND3Jaid1aWPWSHJUoYN2CosvCsnOfzhEdTYtiVIFgOh23fH0Kgq1eXl2lA1QOFVBv
j9XVQE35cDmAx0S39bDbbKkmtf6IzjZJlVp96ZqB1JM4u3dRBXnOOj6K/mD3kcrHkCsPq3iYZa4Q
7KJPjVpgmPpsDJzn8KhD9zx5/N0V1Jrh0Ab4meyN5p9GpGwx9JrJpS6QoV/SOA2XFDyhlB2y8adI
9Rf0sSq2v++hT+XvNaWEsm5SOSrm6+MQPKh4VP/Fu3ReeXzGCjnMY4Dr6Uk/aRa1KDYiFF552f/a
ViGO26DZDDhpLmF3eOez7IWzZzzmY7vzniKmj2NLyQDh3Q2e3WXFi1YAymGRza3s6God/47Zq9sH
J4eb4sODIcvx0FbKplxlyaNzw/g6wffL9VjL2KsQvEpvjP4RsuNa+tudwNCttTSLsMlQpcnpeMv/
WCmvqWfmEL/+17BxgapvdFf6kINLkM9G829UFR3Hc5Gbiy3KewOkejR0/U1hJh2dcjMmLtIuik4J
FchoRACstxy/nviRp2eAA0EE97e8FnN/NY94/NR33R/iR6K61qauJb6o18MhTBm0NM5p54b5ZR2F
YG4zGU1SPaHistF+UUeIOwn8Vsyb54bMHnqZO6n/i39RQSq/tBymYBhF3SRevKaQ/ne4kY7GX9n6
0hJIp+xc9XgQlB/ImnUdRmFV2R2zJgWbN9aSbObjpcT3wsnxxWaQtFvDYSdyBGh+t78fGAEOwkMd
iTb0VwqeFQPttbYjPH7AhCaKXdt2hqnUyopmipRYWJ3FHItnFVfK6t4MuPPEZs0C1Mdh38cs5DsK
CK1cs0n6Lbo2puaYkEfchsr/UHAwoBJpAX3sVgar6SWUZBh9pi7vwrHxaP8HpQVZvCOwXTijq5wD
u5cRyR1kC3uNhYYVGhgZwc4P3uPd65YzL+QlxsMBvEp1tzGJYqR8MyEBF5FGbbtshjbhk1+zd1KB
OgZwmXvC+U4OVepwvz0IPSrLjCLcsqq/jw9a6NPr2C1U+vJxof7h+LlKHGNm/lcB+WYc/hK9/TuV
oAjRhkR0Yf/muFy76sZhG0olZQwKNSjxsGB8HhomjnNePkzaxXlCgav0P0Kr4QJuSWLFG8mI26sU
ooc9iQYbEe6IDWoIr2zZMQzHZVL9HzwA0oKWqHaGMKjZeW2MvPVTQ1OPYqdrLPAtK+H8FTKFb88w
yerTgKBOBHGUxpaWc4uV4OdOavSOXYyohD4YetztntrZ71LciKX4T3r5trGUeczM107iJr+SsSIs
Omnb2ruMFDSvOXJxr/z5fojoxQwX3WmYo2Cjpcc1Xe+iZVdG0tYPT/jp76TQgiFKpWYNgZCIqCjc
nb7Kr7ESp2VeWBzYwnrHNh7vcBy7KVSESuIaCPxyOTQjMrSkm3SiJaBgQiVvPqAnYfMAJ+aFMOjb
iH0IlbuBqwu1hLZTyuqWxOVJ2D2ujqxTfuZEhB3Bh+5ZWAoLNIFmTarWl07+w5ydvqJzR78yXalf
w00yY6Frh/5sMaQGMgdG2XL+FLKfR/ASgLo8H3JIfZdQebqOcmvQOwu1hAz9O2RqSXDN8zTrFuEJ
xmSrVPK0PsjKr2Ni0swKrdzELkmsHTKp9X9hmkt9olHUlHFZLgtgcjPqUyZOVpougcC9F1GOnWsx
XUme0crZ/es/1d/0F3h85ByCh1ot9tNuuv+LM7fN8Rml5HVRlqsP3bsm3YG+ZAxNt9i5Pd+vTG61
J6l62pJuxF1r5dBV6lRF8B9IlFMBz+7+4pdLWDzaBc9lX4YeqD196cF2mD/Nq+lJOtrrWBqd9UgG
Wy7vs78MDLVbyJR7I3s/JRbuIZ8AuI530IpQcyxNeIm2TDY96acgxieAaEEhCTBnnbfo8KkFhzn+
jlXDRHe1PPXwLejSfgj1srW71LVOTmCRbuddAwLaG6WX/6i5YgH8EUhHc+uwmj9GL/4Pn/25IkyE
2ODmAQbOzdwva8t680FCBcR0RS11x9vlIa4EWfKr0Vf2tW1701okMvMRmyIw3YJVPelgN+fTEMvs
JGMOLLDleBBjLF9qEnywvVdkAACSnHVNODVokDJ93l/HoKd/3FZK7kudlKAtGhKOLLXowzTpY3ro
HXCIPBfCRC0nui9CUcb72wosRi/9zQp9NnxN5Ucs/gFv/bKNpB8SB3/yHnY4RX0D6uUC51+OefMg
I4vQ1x0uVQ8TX79XP5X/W8BS97n/WyQhxl0oDNDS7Q6IQ9DgWICp4jmRM1JAF2hLMOr0sIKUIhg5
/s4Zj+CP6tl/Iwwmcz93ubP4yLGGZECvZCAD4xUmEI/qPmdF1K4rw0LN3PjmUx2nGBSbXz3OM3rN
GUWqYfEjnlBSskjJFvaXyxHh28ZvCBp+9fQIDqLxXVJe1mUtovhrehCUleBRpG68odROo1Vs3nL1
YH/eCGrKqt1uVRrWwKPtyfmOT/NbVtYFXmh6wjZWQj/l7zgoL4g4dN3h9bIVReAFqArGdjKL1MjP
yOkyGUdLsToSvepxA9OqoGz+Oqh47XltYFt4RyXmfcaYJAIETWiIyrOT/zSApwU4gjjOU8BLud/P
QLCOLPmYw/bvx3ZleNDyDj22Qznmdci9X/o6jdTuHOOmi8T1SSAgF3juQAmM6GSQD0dAqpAP/jJl
DBW1gcNJNV9/OVAZ8wQLsmBxDanF016cb9YR6vylGb9Eq8o28hbqOTgkCkDLnmAszGItw4tNKyoU
iT+qjB5rW9cMIsH6qb4rK8k8cC2p8yT9EgfOUhb73XaQNIEQ4J1orDili3nd2KgrSUg2GFj7wAXl
rKMdy8cdGXeaB8DwBgztBov2XljlYStEHdIkycJiFXSgHd6+oeoLwbIABoZXzwV7v/4FT92ZtTgs
Q2XsLZzzL7To05fG0icWMweQipn668C6dHhTci9d3OS/ue0oni3B26TazuTt+m9ts/pVqCitfNEs
/tdmhO3Jbv+ACDmebk3KBZCKJTYTtDFrh9BWYE/IpqkO67h3IidfNZ5ZkOB6XUhgW/Q5J+dop67/
DZJOXjS6jqjvqDgtFJdE1doAcQOdfVikDxvjGIWVxfolG2yJeVt+ZT83ko4IPKwIhiH0Iy+B5H32
G0qDysdzz0qYOFiqcyNF5/UQjckNwntfgqw1RVMMUoJnqMPUPWRqAXrMIUpQK7bomaVqJS0CqLyj
uCLE7CqncW1RvqswwxkF1mK+ks6Ke/R0EaVUBFsunCsaPXlo8XDx8PZvZsv2r5CBfMHUR69qNB8w
CshwxLVjmnTgxx5CuCrqSqSYHeGm2dYc52yoz2bz6O+Fpnn0ik/AtTyyUDYUAKzL6PeU06q0CjVH
sI95lpFhrB21tFEwCmYbH3EVZStAl9I4bIfSLl7hpEaGOFeL4SiFl9I9vkSUlaE9UridvRvMh14K
vRgeH7gtDHgyBM0TEnUawA7dZgggnJ/HYgd1E+kork4xbRGS8sx44X0nVy5q/0VRaJjn6n15L4pd
LndjnAbSFMBlQ+qu4xcCqNPUQ+hvc1WPUY3wOEQSxetO7vOK3b6heolsxh9gNdJaSH7pCAXokEz/
mqPkKNipTsSs4EdRQwmW7wA/Tvif97Z4CDK12lNuci4DFo/2FWsVziLP4yHK8kNLM1kUBfFAVBwf
TcZ8K536pdUdnrofcDxPPXTae6wEfJ8Ai6YVX+3Pom3q08B8KRayJVDQt21CBpuxOM0XJRnYNPeb
GhNt9auE4WNgqputUjGXD1dQwwUL7wIUKDu4tiWgV2/NmLeZB8lGetufIZ/WGxIH8mOL8yCT04FE
1SA1Ilj3bhQ884Fiq811IkV9s7WwkoaA4/AgB5aS+7a9CXDpCT8tgiMiIKTREu/ElXMchMynz6Js
emxqKRzX/ILQgePB7cR6rKrDgf9zm2lbtoPv+pBJ2ilMEBhAXrc3cJ/9s1GqgZ22ShM3gdFJVkcG
6rmXSPBL7lCxnYSW6896Eji+I5LhaHBSy241orRtraCepPh87C8NdQ2e2DZRhxUB34aKaAUg3auO
6NkSZX8WUZ32smgTT07pI11gpYG5qh8U6pNYMq92gnto9n1JqaCM/kl3Z1OXzGbNM84VR4HhC8RO
qfjD01o/V166AV4Jg0zHTqENPWyDcusAYYGM+XToZ9zzQdJOCZsQKcBniXoH6+cZQ9Y93TqKHH1E
2PLcQOrMDpzyR1mJwKKGGy58s3QeHqybPJGm+yWazYwpYpRvYYf9s7A9nuw24xcz0o02/HFZh9kh
vSjOOwGy68/gSb76oORjjn6rreUbaW8KygJgKRABEDGB8HR3BDE2QpXSPntupgiAKvNLMnylLRzk
Ed4nuzKEOKPmXJHITGEwlTftrOQj+eU4LLkwgTBkxFaQNY1SV0uvAxUCWlLDaM97S2c5f2IcB3Yw
8K7g4tq4PomSnyfB0WHjSZy96NpTNa8HiastIYKGHsS741g/oZDkQZbFRWUDhWR50R9zOQOBfND5
NxnqzV67Av7ii/zyfI36Pj8rxYcMD7FMuEUZgAiIIXk7g4PUu5DI7j0XfhGbZMFcfToNhQuW/zYT
6YwMNdw9AcrmzFODpw+1pFzm42LQ2WrYqbvclVRW19UAhU1SqzU+1yH44r6FltYhUj4WMHf3A0wJ
p53vz6zJgP/lGt+aIhDvAj9en7vaUZNJ6daAzuXlPVTQhzYRZFt2YU/lQNX7l5meaS2tFKewVeek
sj+2UT0JNyRhTAKIEnrx3AfTn0+1AWr/SzY9RxyQOm3h1z9r/KpbtySEUYiFlYX3j4yBA4yazSzA
8gEez8lx3/42qmy2ZS8Pu+E9VFxuwVhLhapcZ/nyiCXjZhOWJQ+HnigFq8IqHUe36o+xmt7EC3/M
hUS/Rk+l/8FPvCTA9rf/K0IZVZ1xQI6O3WvYy0oEaARLbKglzpjWfBY35LeLA5IwRK21ibZyWwYT
p2UtFZRFVb04ty9rgc/m4/4kMqWq0NKGAkwX5Z9mXZ802cWHGVslJoH/suWkgKaV4zook0XtEtK2
p7YRbiwEMG9eEnWUV+bJMuHagodqvLgqXFQSCOn4SHRKe2SD3JoP2J9nYe738xo76ru9h2iTH4Ef
vGzxKanlddNs4NUsnpSqZla5DiMw1IoLNTXSSMFHvY65p1K0umNANKVRxzIvNhgY9bBsg85lLbiu
rvX8pUN4FWAAtnIE+OMQi+d5QwQuloA6Ex8ejDQZ73JbNfKkY1e8EY8VJVlrYsbCRJy5zBuNVIND
JgpKEKo/6ID3Gm9x5yZ20kRgzIQwkuxj8pWqvBHY1gr/StpI7eShBvyF984ovE2dAAQ/hr+LyAA5
/RT6EsU5kDiWIBrmjgRMUYnKKZU30e28lBDq0sYddf03MD7S5akjRg/UFhctfWew7cblFfZ/7bnW
m67K9JQSukxaujVKFvJ+/5QRQSxaLHqAQcJTROv/Whe/wHBAAVGbL4s+YXPDOyx8sqxfd2sNrvuO
yZv6uXsi2F+9AZ0sEMbx3O+6F8xOex2nB50KhmkauRWWNsPy1xa1aNP4yqhQewZgV5D+V36nd38I
Wx6/4UzrbIGkfcElU1mVJht1mYLak2jjTnJWBgdvZ5ClshTAN4CiwOTI/3Anb3SQjMa+TeY7F3+y
4Y4sU5iXvgLetYsMXGvF6tKi15v20Yw0G76LEO/fGck8vVWGQSHpcnxTu0S3CiUUCzX7hXTnvRxQ
OL3qw/kEhn+Dbdy5APEvl9uIQljyBET3nuGmsIxkJf2IT0NYCOxP5S5TLEc+5fveRXG0AZ4eXksn
xb5lUKUVB0WmCjM5oVprqZZuFzTAuQStv4VCX73A9oECGKuH5jzSsXXU8F+2qQpZsyKg/z3gHHtU
UWp+fOHK1/f6EMvu5aSdEWVlEr/DLyz88LDDWepp+B43jp9MhqHNhrB4QuzfPfLkPc/sBJjTs5KO
hQw0rSml39SB6MDYr/HH6gzeHuxqJjUXD2mVUUwiOKV69T0qB9AHeKAv6INVZY8smhD0ho9PDjR4
2qpi/K35uiNFgYVTrlfhmkojqftQfEtxXddcnr+teGDAurWbXXw6MkroXYfVyThf+5R7XuLic1kB
D3s0vLneH3Ct13FDGQvxZwk0FAn8dAVvRG3CsazHPqukfRlPh4FJK3vmAtAParH9fJUsCE5+qj2F
G/YA97v4lMlCsFrbdcIhnJZZIZTor4PSyF4yCtTqfzI3ztXkwyVneg1FUqKno5B1emPVNyG2W7xR
PZJ2/vBSdzb4jNNyjgzelSWz/Ic3I0623UjJ8rdWsjEwXqpsHxoB69DUUOx8uwcCMKh336DJBjkj
xjZNfnEWhdICueCSvrSYa8rCGIaKOr7kHEy/D3FoRBhjGY6kUF3bHYuD9AeFeetUt9SjYCAoUIGw
2VKL40uttquofNW0hmmBzvJBcS/yq6+Apy7YQ28yyv8dzJmS7XldHZOJggV9SACTD9T3doFrvnc1
kZdJgjfpKokzmseJy9ZLv9p9yhtW1J9Mn9YNfbzTCO1x4MrrNuJ2vqpRinnYS/zRtNmN7G2nol1x
OX7U4gRKSto4ze6XpRVClw0BpzzX8J4r1dyso6MPOUtavAygDQg0TTU6BoadcILvw/cmvzT12JD7
47vDCx4Q2IxdwOs1hc+ubS9zHD78ebgojNO2+M4EKNutjA9Qwp3jnrxbJA0+K537wRKXz2gVQuGr
hLAR1NEJx4c587yGpGTVFFfL16glTQNrtjzNGHtpfQTpWV8tcl9ySTqVE6ZEkPqfaUy6PpfMkDYJ
4PIG0SwPP+Guy1m0GyOcJGakXQiFKpwL0KQwHn4kWJOsjuVvOCQ7mUDpdN+CCydGC+b2XK3gt7F9
KF8Vr5mVk/YAP06CtoG/XWaQoaUUwhntYMH033T2c/XHabXn9IHy3l6NnjMqTf9mYnkx60Ey4GfD
3vLWh7H+D7Pi6exIpWZZu4zlHj3ummnT5zRb6ZJ8zhFCH6sviVxmTH8TNhBnfceQ6s+j/5BUlh6A
UnLAJkmoUKsP1jSnpw66avEUIdNZm7WchnhOCKY0tr/kid43EsAj9oaQiPL7BXO++lci2qjgmR9w
EzyYdZY4+3V37JjjXI5BErydrH+x5OY1sSGxDKh1Frf5jPWKpVGU5boRsXXIAnflp6On+NkAvDZ5
j3rqRhDOeQAX7DVnfMoe3W2/bZX9RhScasV0Xc3SXN42AkLPgxttdF6V6XsR8BohAMpMtok3EMzI
QMLbEouef2+s+9wixsZ9zxo1KgtFq4A94r9aV/m7/BiuMjDqvAYhnW3r9hvQUwhng311K8nTUZAZ
nvskmYQujwndPoHvZ63VuyBWw9v9N9k/099BoKZ+rT8gAybmsR0IBxH2l0BHFUcGSFkaHW2mbEJB
Wte3IeD3QzNO1Giv0awBZrkKVwg/viqVzWeIvKooZ5GB9kxzu4MQsQR4+u/p9PIUEAOpAKJS7dUY
s2weqPfOzC99RM45pt4Dapjszlv+GLBIdEzvVJ2PNAP+5NtnyHLp173m+LSDd819jZwVbr6t//gW
l43x5Q+81ysLRwRZOIlt32Ezq+ZjbjFw9NS5Up75rxsd8aFagtJawD+9XQN6EB2v0cw70yfbc8W0
/otwi7cFyF6RAwyEiEiZK+mTpaaIJXmqUktPHqmN4DKdqJShMw6dsP6+eNxCfEFxh6GZysOOmot+
M15gkizBKUTCvAyM273rZThy5vTrBbpSLelJZAzKO9OhdXV8F+amMRPy8Gr+cxPk3mfxlbKEreA9
+W8HrTYsjk6rw6J/Wg/mfpUgu3rEarqxJ4cCXK+Upn4Ryw1IoNFHkCJUy4WlJT17PlSg+K7CN6qQ
ylnqdxMsgBCpe8/QDih8URLJXyiNDQTzaU5zqTbBuf01TDBj9hZ9SEsCYVX5k+04CzAFBnsvpLwp
jvfGGX+gUQUavahHG0ERlYArn+LbX98EwbLKGlCWM8HCEMMNXitN7LQON7YsrMcSxkjLVRGma6Wv
WneSU9a1YK+7BWNfA4xpyu3gQ/LacqWLkSPJECKGZQ9hrVLnqaEbw6vors57KF7q3ikbRVCjSYWK
aq62SZJ0T6f9YneE9MtDgrCCrOpYBRtei/M0H1Vzm/gPIGZnOxMtBvvnBp2ffBM4yxent7ceayHn
VrHmhtu5Ufnq22O5nugD3v1Xq1kzA1USbxtKbasnqnJBjnCafFJUZnwuH8cr+RDpZT4ZMcPIkSbA
yhf5WrqsjH2rLH1Hvo0E3sRsJlpZkH45s3RqnoLZEvHFkI06PVCjW8NvL7lVXRlTUsH2zjYJ14ow
oV1dl7IFCsfacCx9jx9DNUWAmjw8e3rdMngT53LQEDbaSGbqnDkB9Ae9TZAioYyEXrfdCvDMGD8C
fCByOJkT0MaVq/3NlWcfZI5Qb2UFcvhtozhENllBTs4mM/m7JHNKZwHqtaojQoh8UJ6qG+opSpCT
pzfTltuLwN9MYnNeu++Arpj5FIeA3Wc+QiwY7XbLV8zVgfD/CdO98ACDo5pDwyRJdQii3ZJGRW2d
Pz7mHnQhP3uZ80BfnZvrFhydPLja8UL1ZFfP8CBP2rHWZ4KeYhqookrYAxIh7cy68R5vAvp4q2P3
HG7gSyudac96/TPGrWBjE9W3dUzdO0/dQvFyJXMhxXQ4Ox2WoVCtLkSBenyK3WfHNh1K3TQf5Vay
cgrlshHg4HINayyzP4dF1qCLfeN3Uowr2jP/jpLXEPzq5RebFofvM4lB/yH5bHbsMkQIqahex8w9
aq4rse5yvXj7WKUWbOWtgmGT8DT7ITQMGoMJirx3EuoMDuutQdcvK/rUvWdQZibMxPidGveH88Pi
vQGXnUaGwr1gH+eicTpbixseepGKKJUqN4CnQkaBAXj0a+FZRH5SvecsYe9id4t3CYnNS4Vfczfk
61YmScwP5md+xMT7QOpLyGZfqC6DADvw3Z/VNsGU9smsqPKfVWWnKzIHiUFoPcBXckzS/r3Eo3RG
7xsIVesnEr1AEfF9Z3G2qRzdHUtrg44TQQKJDqhmrqE9BDzzg3Ycw6EHGgHyaKTmdqSz2mzDwgDw
R8XkPgE2NkbcDzwrJ7gFll8t/YHM759uMSjFcQsEIWCuAnGRLQVZb0WwforkNA4CRy4L1iTUtqLQ
6YEOb9yEu3rAet4w2cfAjTe0/7dmxqn50x7MzeofuWEafxqME+SJceoNO70M4wCa0WyY+9LycrTX
lUK+o1rfhbLwdBxcpCWMm8H958eSD4yUwlZeiOXny/9Jv0SsjKsFEoOmMEDp/JBSGKtYxY35euug
IHneestAeIc6WH4iJz8/gnYYvWhei/RJGM67m7d/cXSbs7ATwfHNMYJDnmndsH3MCrCWzcwoPqyb
AAMjxdDTE/2CL0CIejm3dcSstIfUdgdvHBeCS5E2fB/TKdYUg+dfmR3yLUDeCkEg36qCEgNDWaUz
2awtFqxt9oW78lAEB2deTD5l22niCCLStntZXuPiGI5gw3mVQKOkS1motcxNrOG9tco9wCIWjnQW
s/kGSH5CfQgduqw+kKx4ZqqfC1KNvQMmRIWbkyBFdjxWSSJUQBXu6NBDNKOFRdAGEiSqphVklfiw
kROdBoDOixB3wBjW3t31lP3VYn0YO+4LYlW4U8MJZDSlA/jcDp1zhhzu13Dtdvk4rrZiXWnD5OPh
Oufh0+G67+S49aTBO46STGiAS9jtEwR/IAAP6HoF/2gHbk4MuTlsFBSJV8kXNcFQ80ToywvAY7/K
3M4i/bRHVJCe1rIL3clM3c/AKRrRgGf+kSu2HLf6+Tg+S4BcGAdoDcoe9Mto9Rvj1WHl3UG+LrIM
94OJhwJJIuUGN5igCphK6D/tsN70+uPtG1gmj52KmfD4+VU2hUNj++4ZlHFtPDsnplDB25p8XZJc
2HZYvhEo/WH+Mwu4PL+k5uDs8G0mwcefTFkp5bZ/ihutaZm1prceXTqrxF0f/nkwrWiPxVTQc9CQ
mO2m7/+80gkc4gHFudJBGSMr4XgJ80rmUhOLZ1e21+tG6FM/AjvJaH1amvsqOUVSX+eWb//KK5NR
ZdXSLh3blPaNn/oN3n3XOKnCPHJQdzqB0h+hN8PabYzCX0Qi6ej1OuVN0pqYqL5mgx3PZGkm8vTC
rFsdn/kuUXIxMf1qJgnzmoAtQ+q/jA9PSB11uk/LR8apXKJTx5S8raI8sK+8BiRID2MKaqBDvRNA
MPM7eaCeaowcbztUM5gdQHW8Mlbo/1G22QWTcgNik7qlGChyTpR/yBAiIgcb4nY1t/m/SRwesMjB
lgbWzeiWk0p+oXosFM6PaTZS3c1JxWv6s06tv6moRd9EOnWYrJfKv/VRkN4o3Ee2rWkW2EEcEUdF
Z153Uq1h1B9BNSam/CQW0Qqn82F7ojyluAP8BKnh+XbMMbOLMpSyQdTRTT8dJ/5c7d85ouDO3K27
MlFeZXi+vM7skNjb5PbaVDROEzz7kSiaYorTQV/GM39fv4b674PQ47m//Qo4YWx4Y27GHRcnMVyF
s6TVurQifaFAB6K5AFa19A5e6DrtLUnnNwrAdFtsDPM8fO4y78vIMvE9oRqZnzJ/cFtpeDPHE4Oj
r9AYSFIYGxuuN5OTtspDPEhua+34MXGAYl2jctj+/DYf/X/c8R5zARX6VPUIpmOg/uhQii9qqQwJ
D1E7aHnSA8q35RXg/lRghiYbDULKvR85sRBbmxYqM+IXEFdpV01JqxyG9uvZhpUJOVZlkCAUBoMT
9ibW8m/wRyCqjTuNpefy9y5R7zPaWEI/FLxpYT4OMm1Bdz4a4s/y7s27BAsFMOLo1PrIHDjQmy95
Sc9LrhmExlM2KJwx1t7nfmpoFIAAHr+LxKMhAui09gdDRFAZJRr2nykdm6q/RVkJfIyGIbmBE/2p
iXFPC/oiR8F21PvrKbqopKYDUd4wUMn25BknsyasJSY4V4X7bQsHfcJdgcLNOJesa/3Nb1gcn5F8
ZvQdQPRZtIXYXhe1vm0aYJsvXvkQlt1aTCopeVRucjylKXoH8eGmtP4G2grcFbYtUQqEmupwDPwM
+gwYUwQeNqIhq9ze3BYkQWsaXi67yqnN6B/Q6BopJvOxlNIPDtPQzfUzFCPF2SI05Gb5eLawcGvT
ZmD0rLgG97KyXIauKBY2E6eJiZzXdt8d1MGn8siewuvPZSngZ6IbA7oMjDWoQhratka+G/5i7iuO
ODtUFTzF5zy22Scw9dJIgSMUNJRlAQoBT/5Gg5X8JOeD9itxNjU5VE95DlrJx7qnbirUwZLVzF6a
//HwuWqPHqraFiUfGyW4Lwg9vdkDO7MbHiO4hMoDKmHZ79AMmjtteOugYQCznLcURbSdQdvrENrd
vHspjoW0om1ClUa7wPTLUZOUo37CXFc51WAWj0cfV9Cs0tCZ0l6QTdr2wT65LPn5Xgo/2LNi6nTG
N9V9TXyvHcb7huZIb0VLuOeB7OO6/XjXRAkdE9oLW3IAj4u7W5EH+4+StUegJtt3WTylgL8ZxeR0
2VRyxQ+NI0qLkw0mOVpAZp27u2aHmLUDfm3OIrKsFSqjCLDGMEBomlv5JmDdu1qhiQYIRYBGuUpy
+/lo82gKWQf4kfSycYXa+pK+jAd8Mx7rsZvJZa82k0kKlbRcrSPFV2ljR+cuSB7e5ttt4zwCo3gP
Nn5ntYGQ1KPLNXkhlHtSTIO1ZZ1lfgvsvXs5zDO4lCe1BbDtyq/DaGDdxXfzRgVxZa9Q1wfj6cx3
rWpzRceWNo4B+lkPrSeFccQ1h8nuN163bOyo9oUFReVp+NOmxSz49rIt8MZQ075JyH6B7Y8RO95a
NYP7/U1zEFbdAjAJfNqZmN3Itk1KNf26hCsj6uZ+xVoB7SYIo3l3IrXTWOKGRasIa4PsF2jJiwUu
GF9+G+JD1Vo7o108LAk97I90WZx06a/Ve2d16ryQadqBrzVFlIEnlRQTJxzJbA61bTRCQ8AbTAgG
kbGRWDmBb6f/BbgBYWe/UKZUnBnb0j98W+43eYX5/qDEVMzEFeL9Yjg5OYyW34YZ24kgwfAHB6KB
+XHnYboFvT7gw++raSLgltoab5d+Ex7QShgltvVuBq/vsuZU0fRoPtAv/S1vuhCpnUpMCu8kUsNb
l8w+BwMCRsmRsbbw+47OYh8Dwji+jVFSmombTOi1MIsU6rD/yBYfCGMx7wLqhkZP6AUE7BFJTQ2b
9k0lPlEhXiZIQfKDWSnUcqOs70UV3R/ptytdWK1eTHXyndWsjnU0F0TvP+bV4i1oDZsPGOE3m/rZ
bmpruZahyK6oVcwV4DEIIdIbDqMBDhdFVv1w83Ce7KaMpEwGhzrEwRC7NwhfuAZa9J68HPkHwwLr
lHHQkAues+rNsNBiT2wPdU85PGeqUgaQUL+Mns63km3NuSTXqJ+zkJ2Ki/LGhUKJ7Mc95qODVTyC
cyq3hXqzLF34TAsplUKZf0Z9MpzMgV832TgY/zc7yX+0IO0wsId+kVbZjuqzuJf7ieBgYXVbCoPU
Smiq5+od0p8ad3ngyXmhjck8hrk453tKswdxs1v4obqIZWpXiDuPHbw5FOiNq34CR/9lE/+D3+yi
PI9h8X1P95r5RjpFa+p1Z6DYQrwcdBjtcqJgfCd9a29dt4dY3DYMBX7adiIbs9lkaLUbmTQAY0rK
pCYVQ0dpG0Oi34NHHvEtdHDToQDG2qwRuIHQ9KPj+lO69OU5YsErZJ1HqhOI6weB2pUl4R7Sumtf
DjXJAnLm5h7Sr/lfRzeVzP66F0mmmIFjiFZboCsDg+ubF/BKWMXy1RdBoUEO3Egz7ZNG11t+QZhU
ufrer/hA2GuF4UgInE3/yj16dJkQatCw9p9rfqraEafpDRw4vLG38yMmTl3Q3Yv6vyj3KM3TBmVW
Ltw5aZHdZnZfrDpUODrusghsCU8dM5TyObHCtt3GGZvCesNYp2uE+owk0hDkdVag2iRMAywKZRsa
2qt7HZ+sEzhvcKjpQ/5uKFb54hMbr8gkWd6ZmLBdXVIuYfQdjspFndlkUyPpGot5RdG6UF0BmDW/
5JGQSfifgbEZHjjQJC71eLC+0575Gbp5N1c6uha3L9bWQNqjSB+g0A8NqKfC7TV7zOEJwyOT3wGp
s7Khd7FLAulpMRKEtqUXDY/GBh6a+pEGlLbra9diKxkA9MMdK0RgsysY/Uyc8Go8b3wZ8X6QL7rf
x+OJZGtYKXyFID+PdB6VHxwNtlI+ojHWofjXYgjE9RLv/xaxXwKGX5Sjav+vm9q5gHEZM6B/p/Fq
FWWqR0Dy+v72X05XX8xVfIzmKE02cUkP5cqdZLSt+yMsTYvPUE8kUus1tsmRnybWv8G6T2HPGh5R
/qhPr1WR+XnMyrsMYgTWjtMA+lomHY93d4DZQGD6ID9tak+LVj8cbfBvG5xdSoeLPKxlAoC9utFt
BWpAS0vqkQzdE73Cy/O2Vlecg4JM1/nH+cIw4ApT7kee0phv0ZNQOqBvYo8KicH8iKthgtRU0Tle
0yI5YBubKNWqXjaaQ5t0e3M6L7634C4XjbVaOS5pqRIO95GRqC3JLYReax2nvjsXo8miHaFsTRek
QduHt5G0nFdvRg8U0wD6WsiAMnDvpBY0Jbsv6obEN3GojNf2HDbzpW/RvTOcsvqieyPZKikwTPPB
lK33HBbVCaWJRL2MAOOlG4rtLtl76/FDZHpuGslkQ6MWRuLDwTAzgRBlsSegiO9mAwiuXZNk8Ty5
fCzmO4MVZH1GkNztlPvGdMSaJZXaUKWvWwpHuJPazOVWv057n9Lbg6i94gTdsm3p5n3KbJgHsnMF
5N9L/Ut3ORX1xU4vVO7lLSpASqxBzJ7+K/hBtfyK7mG8BxjkqAsyMcLKGmQ6LlBKSH+c+wy+HtIo
7VGgmQX1RsWJ+sUrhjZqT3L7EhJCIsJ+k2OnIJ14Hifg1fRhyQ7lEGwCMy/DG5b0M0oFXdZT7TrO
ww09eRDqucf3vkKSBnC4XyQ38wDLAAqDmN+4VYgYWojHtkMAm4uobwSLV9J13SKka9UMszKi6UAw
uiO62Ci/SaM60a8k8/bRf6h9R3XZrHHWZuLo96kwYbeTfHU4F56YUSCOpgz/7hw1NPxHjPt5eP+R
2AdgDkOdj0JmlLfZM7bVaiMVzGMYuUqfO2UZqiCVxQ/H6Uk7POkZ6pMb1YwCvVbWLPXKT3VWpieJ
sIYUy6AYFVq8a2/IZf6v+z+JUJ9aBG75JiQgJmfmZpqz+EGTL6GCxW1mVkNGTj7smsFR97fARtW7
0XfLhTV8DSDDzh8pNm2XWH4dPdZtCUAZMU4BBgt/apKS5mU/Xlf/e5xbifYnw6BmwJWqE53IYvDk
e+vT/zSWRiV6cchx5JHoWpOtOvy5gg/iiHFIKFXfn3qil8PVpWkpD2UhwD9f5mFgJ+8XVu8C4GWT
QIi3L+TCbRbgE/ofwLaUaM2YRvIEikBxmLU15KAnnFRZHyB+jFjaQrKl9S0yFiBtK/9+Png9sGpl
NQgXt3S1sBVaox3stjhU1OG0B6+Q604U+HP5qWkb6f1t2ethJwZJ6UZ+LHO/iK8nbOB8l1rowyJt
TRtvpzgXLoRYX0641YO/6RbSvPlSzW+6hYMQUTmizZZMBL+2whkKk5ZzAjRXLkUGPRLz+bAZPH6W
yfHoULjzPkanqMZCfWbwhHs0CvTzsBgx6EmKWuSnOH64IllQ5AD1U2QLvxqq6QiOOZM3vYAJPz8j
JBowpzHrAba0pYqYU/KD1EvT3CaPrD/5Wti+f97d8uWP43CCM5QwXG8NvZOqgy7Lh8LnAc810LdN
6kOzlg/krlfTpvIzS3GZVkyJp2bnJSzLr3Gk7Y1jD4LUnpw1nVa5OrZpFIyIlM7CEru9W2ysoxk1
XjQuBl0TkFaLk2r9QwSA71U11itxMHkljVh8XkCQ7nxIFGtX6NegR2ZogZ71lTVbI+BRVyLysJ5B
Ph5UgUPI/bRch32N0upL+MZWfpesFuz+tFidbC9pbYtIOXT+gze6oPS4kwDO/d1+5irqNhrRfpQH
IGAyUv/O2Ma43zggL/HHf2jio9fnCAhsBcUzJVWGeMLgVVeVVqvoIeCnaKRfTJO7Jjwlmr2iOlxp
KLotvEqm8g05YolVLOyKy7YnaHMbqj9K3sp8XRNTNR+8iT3i52Q/eQJO1Xc1iVXdbS+KidFuCJ9u
oFlR39d3Pyt8CFRoF2yLfMu3Fu4uqDf81T8mcrC99OnM2LbcgmX/dpuN+Ysicw3PzX9HA/JJ16Y/
h4Jz6lPF6PW1UryMfC0pZQSAdub70Zia7M3Go71qFyYxLbbnCL5HgmZea8r1shVjqlic1y6Qjdlf
MsZQZIh24Pf91wUBinqKCIf+seShfrWNnPPKswJNj8/bUOmoJGZ1iHJ4SNq7oic6iyL7dCYf0ZNz
69RwizFTQ/wLBlY7YaVMvXcdegKUZNVbeXg277HloN5gRaSv01xyeh0LpWSeucDDKOB0xxGQR2XY
6uMWkSawONoHcvBYqVyR93G6lNBYaCB1u65p03X2dglvPHkC9M7ku6pfLtjT9gJr4mg7+E3fegkB
cwa/XnHx0GhZsaXZBwj1tqb1iAWNnl22RDeHFOcqjRUcBbLhwXCIlmzgTWYxS/uxu+7cVoAlT1Ff
g77cUVQTFtiByejkgE259QKf20Zxl/BHYHXLH1HT11ZNvFOyq5dEw07L6ikVHlM9lv3Xzg1NInN3
g3sIiFmR3yPzdLkHgExaPk3u84C+UhQk4B6BtzzB0fbUjMKsatlUaGHRe5ARGEfKtO9QCIWK3B1P
DaLGjh0Sbo7sjaxYzM7EAvWu67FN6fEniTeEJIQXMPgFUsTFNehd/D1bY6ynTATpRlPJcn80g9lz
azKQPcVamJlUaRCPM5NflNQZhNClTonXXj2zRAbBI65UhI60VUC3majNN0stX/nJ8MCVGIkjHJ9a
iqct3cG3tHpTUS6fxaHmFvTnzJednOCPGk6ozV6XW31KSOkLzAgFY1Rvf/0kTt9IAh/7zTGT9ijf
mS6MvjPDMAC4rfPhuE0b5a+YsBWMLcZ04D4EUqZvfojqXTzhU4nKwGZ7ce+hukHtcVS6HJYxQiEk
DahNrmHxS+vNBfXSKJSlsLbnm8np9F9kpevW7V3nCCwwdUnAZdoUrewkJmzBxJe8/Clp6BAd+vIt
SfhRzerUIfSeDeXth6Hn1lXg7vS7iWKgrAl3+DguNK74g6w6kMnzVMqpkpmqbYPP3QgtUmq+5NkR
dvALDoQ0XQG99tiOsMmaNcbQAz+b+NGtmA6g4/GbAE74Tqtd4MzKy/e88j6duWqmaef1HRW028xE
2fnvEnKfCgZcY+2L1/QksYYujArE9xD6BFoWuZEhR3EKcFr7nv+KRzeBY8noTbcuC2+TG5jE9Tj/
8xKQo5+fd5kpZJJFoFVq6xundiJzfHwQoQTvLzZ6wgQ+3sr7qsJnHu3Vh0LaK5/1OO3ENXKC505d
PkD4HyIWUqgeUquKkcWE0ExXCoDkBhMXZjHg/6K7PMgSnbVGAC/heVRG3waOBLIU1EOvHXxksI1Q
IY+VQh4NkinlCFqdtaK/0hBUCEjy1j+OgiQHuQxEXLNOFj9viZQfHmuXn5Dv2wTmjdwrcHcqZ2T6
pAfaBtJKo135gd5TesIhYDurh317a0dwp3ynMy8uLVBHdgqNgr41pkXTT6m5hNvAVL18fSUPporm
AFv6fvE96QbjIK4anYIp88Ve0WGoiz+/6tG11c3l/f+xWpazZV90+7gww6jdbMYBzHfYlzErZtdJ
MDFErr0vTIA2SKYqiYy32l8gp+b2LdQbAS0e2v98q0QrQmBnDafGgNhcJuxK8hPVfj2quQ0O/pv4
GN8pl4dzPNOF5ThQUOH45WEFjVoAIg7bfpNr/rnBGXo0IICU77zo2S4cnKOmqO2oahKUlgzct4qS
ILmMykVJ3R5nNPHvMrdj/dcWg83Mh+jcCO4sojFcRZ9g1oHrzFIIFGKcSG6kLmbT1yxIR//smeWC
9xS1Y0y86pLVa3FmNKHVbZkwrDmgpa+ILhFJ9O3eXQrBI9pa3L3qB/SfkLxutpWJmATMk68Wc8xi
uR5o8z8BYowa1CTSi/NjOgqOZdGopcbFteZBYcfSGnSqS5HS40Rdu42oH0VwTH9pRR458ABJ13o6
xsiNEMGv7aOPsGCcuG+74JmGqByY+bXjF5IFO9i9jA3y582AFxsUqAPgpbIdw/x8NKa85ZyJqGdQ
kn6vloD779Y6/iwhMJeQPmt9H5P8yY/09RhROoTYB6nhRLV1PcLQ/8xiFXarHdTfgX17KSYuDnKY
uE5xF9v4a8dbcqucNIRY3v2VoMu9+3wujXPNHx270w4eRslB4O0OGJ8SgN/5HTmuAHJ4CrvewUsS
SJBRkF0GYJYF7cowY9b1He1VlJe8c5M/yy7ye/AZsnW0tQw+fLqiDYAa00CdC5QJoaBsfP2ZaHud
TOCSywQDI32FC4hHMUVV5lE8oRE0yymy3ZTuFl+lrrK69OEXZeAzJTRAtIEDt38MTLG//9c9GSDD
jRT9/bJx/1hahGBqBeE1LyHt7r2YDh5BGIPvA8ozsk7Qp2eze2MU+PAIWMVSTaa9uB0lomfroskb
HIIlxsHKcayPvu3aco7csiw6xCeEmlOM1h8dpr4qBd0aD0bqFA7ODCX4lIA0eb2YTDK+2D39ccvY
RFJqLdf0jfi4MmypMK48VUsMTR/qB03ZP8ajyq/9L22CmA3kBTkqjWupVMDltm+MGZZHxMOQ9wEc
8EWLCO6g83f5MPKe/3UYrD0Lev/rd+q4GXAoyhyENEED5PfEuuNwNDki33IOoqavjA4mePW7IZql
ZYGFMyv0pyz4wkNzfXIT7kgJ6QQ7Z5lO6dkE/bKeQjz2cOh8R+snoN36QxMmJJcPOjU5AnYZE7fP
d3UBrbfFvpES0vZJeeMY/ra+waDIedA6s9exwRb1s5dA1ngy6F04ihk3JbdlUeWJIgWY+ME9VLYe
YUU1LHVAe45s2jeRZ0rB4LIXmJgax5E2n4oAFC4aFstLqShz2ZhgruofPnucEFzulfNW47DuSajo
2euQzU9vI/k/OsJNunt7jRHJLY7Nuq2MWUVshsa/vkW3/rJubfuTt9XZTUsALYj3/NEGBhcIoHb3
ZgHVPGCzWs6QTQrGh/5Oc8dnVZvebkmd3giCQStniJYrP2eIrqJbq/FhMbf5GRJpGSYuYknQtg+R
z+SDv2Dt4AyaGANjmGfY0rCXvo0gchwhul4SugOmjFg+e+YIw/bSd6kr5ApIhucWXJjJlWqv/qCR
toy1Doe8fM7iOBi7KQpJChmpppWPRctqszPXSV1O0+yffhdar0rJGemXih5qoYzW9mgGqmm+t+aH
6pltWPJ7miOJPV0Nu+W0tBQv7bf36gQ0gLIdB05OL7IoL1DiFnQWDyETXr5tpou5ENOX9yDmy9P9
haMzsJNhEBfuoB/iuGiLnhpeN9kCDhcQc4pFPbF53/yYrX9exkCFzP3ATkzVlLde1XLf4z00CjHF
Xvsbdu0f3eA24XELaj+xMrg7SpZuP49Ok++d/Kwuh5v3Cx2x0RFWgOA+ph6NGn1wEPsUr8Eo2T2q
L/x010g6T4QxasiCTfGIPpm/SUCWSWl45V8DSQHYma8+N/CVLl776Pa1j9iD4/j0gwjbmC/+Er/G
c30Gmo8tr0vng0RKl2Scn7brQneom6hCgSi3e5LfJB9XvUUeMS+TBPZmBWHig19m28D4yVE+QUzZ
4k/O9DOQyQDf4fhwJ33pICR2snb1WNL43WHk8e362Y1gcNb8GOPXsaDDEvs9Q9AJ6O3j5yHEybh+
k9OHYNcESTA5biqDk6dUy08fS/5+pXR5CpKjjYzRPKpzfYl8ZrhezmTBclnLOqpB0S1gPQDBfAUh
WES00P7DX22YWtAwzH/V+d6s76LJ8AhQadPYFbW5LNr5KqXAtItY4+16DblH7hlWjup6Usyst7V1
8x41Q5STk3R1JoMi69Oz9T3areudEPZFnx3LUDfZfIb2f6AbzOVgV1YjlqfvmlHAYzXzq3YqH8kf
7I3oDZfGtb/oFN2yoTRYfT/25QG0MugqPgj6LZ8yKRyRrH5zzmAWP96kpSPVeJzZFR/wRCFgQdWj
+4MwKlAkp/If1qLIJozYabqE6euu3hH0MO/rMmPCTeS+iivsEkKvPKNEdu2iiEgr7GExVDZOXUJk
da6PWwMuHOBfSrNQ4HQNnX/nNCCrZWenYLc8XG1xMT0RHQNzOE7I6kymsVglGAv6mhtRQ7jtTzpL
JkdnahNAJISgb4jW9v9iae96ksltwiqCLtbs2eCAw/+sk3sp8DFRpN2g0ZKCWJ26cZZtKf4nbZYH
mgTxg6LWfspGN9yzVXi2UK94fpmM/MwJBQVdY7us9qC4L8wN/Zc0YDj+YYoTA7uxmOwhNUxaRDjw
cAiwcyx/Gp8/eXczO/TCAvUeNlUtXfL3XbsScUsfISEBSKaxWFzLBtZOQpX4MTC8rXK9lYWXOMbE
OS+Opx6E7BSviP7NQ9jNEMZdl41Ye7zFjapYYQV+BdjJNLl4uIc10PYeaQ3aozLD82kgGLLIQh/Q
E7WQif0ufIhqe4nP+MdiorOkGbhHE8hBHxq/+vcFhKk3ry6DwF76OBWnA9DYQsN/9TpWMWiUyhvK
lBpHzjn21DfDjjvzaAJJEeTSj5+HlqsyZnj0UK/p6mb2C+aXPFdpHZMRjVkIBfarIfk3kRtQRpfI
f9keqTrW2zNMpYMQNK5TKiCt5PO557RboTPR1S8Fb5etphepmri8Cb2PTTJLkVJ90kgX+lqu9Ife
+MBib2cOdP0IHUmKiv0HuD5LeHR8Rb3zvEsrVtyWYxWtThaqBeuBrrXKBLTGxmvn0dMrKcVLM/td
DcZlBpfO4nUy9sy7A8t5aFTvsp52iO4sr0WuRppdtSZYCkUSzb4jmYspytdItsHXSnDLKvUK2csC
62Ls61/gRZWFNpvFnhtDM/+nMMmPbAuJ53qkPeKm42Q97Lc6lnV5Fqqa3bZhHKWc3A4Mf4cVdcKR
RyOCTXCRq0E9zqslcKff7fO2+Zrf7Rmu58oE0+8SD43S+zuyjH+EUSXxFiwJpueTp4fCe0w7neXN
hca0J3KWnaZxFkML2BsF7yZJ7pWxGNAp5f2TfjJGHNrff7WTyWMNZQJyjp1j4iZO38L12He+LoQU
E67Ta8bjgV2Fqb3k8h4+tFZohFsWB7DOE8o93qrYyMVi2m2AgYF5/HQleBIbJQwjXvWLJA/OQVxE
je3KKxU3kLe8f9qAYfSJ8xFO75frSZ2pReddNLx/6lcwPYtQfdc20KxUjRLtBex2/hXYQK8FcoAw
4YG0U3bpW1SfQ83jGjOzIILBIbOiMwNpP7pb4hFfkXQisCZlNvablTDZLb5ubenumuCSz3tB0Uv+
2jOBz2Tj7CNfYXM9iMPLFybwo1ZwEPPFnUyrMhaSe4IAzbn9g/DILweTd96u2Dyn/N6+gGZV7R6m
VHrFKvHPYKlDFfQxdKUsBHAXyFKkrYbnZJ6gKKvyiTHQuuTSbnTUvAxCIX9FBN1ob9aNkBGT37Sp
BpJVHA+/MoJmlNxdJs1N4XgiPdPg/IS62iMHup0mse/3yh72siqS1YUrS5wju5kMzk3/GtWtsBhk
6nkwhDNinRcT5UrTRQBNKRigRxDi3AU6jyg5SkrXXoOIZWGfohTkU0sO6mA4e6gNbwi4OF53ff3I
z9fSye014ksyFzg3FItFxUbr6ao5RnS92jSUvpwZY8hCIpVYUX0DXBYxvyw7WdRBPlBaCCovQF62
FtoqkyqPcsuRVL4xiqkVr6MxCFdUFLTLnPZLOQUunZUn4n94/MCDjsJekV/KWFKMBxXpKfZ/YV0x
uHKrOFY5WuRzZFUgzafAfHrX3vVgoXJw1cQySOO2ICijrN6XhTEk7GzWT/LwIWE/FirBiu6LJIAr
mqCzm3hLMip4w+PGTqy4DbRz/Lc/3EntdVa+FdOyS67Yf2hVkwmmesEAMw5l0rxVzZ+LTPTz40Fs
xzbCJxZdtCfnhVJ9xnDaDo+eesSuq27Ge2b9AHxbI4t+EaO58DhNHkRMUXVQ7Bi54kSbVmgB5XcW
5D6/sY8AEnNiasG1puL+mvYT/9681qdKUpowmaQcDaVtNJVAXleVsScKG1gXhgD8PtpGVGHbgtFt
wwmNfVTEX12fumSJC5AZsyGSGSZWAr9wZBuIwZSA0RuQqxXTv8DqMVdVgXhoNfD7JNAMKpb+2IaY
YJegpLyM8yj9eP/rTnr5t1dXA5G58f6tB39acZqyrohtiRjLjQG3inukOADg8bc3IFaBYstmlcdc
uZZV+AjU8glY+W1r+dibWmcUZZoyzJ1RqsWP+0++XTF+UxSz7e7pqJei+MXsfesE7M9cploSb4qD
XWpGbNqDt1/PY4+ZmnngDBmeqtx1IeLecOEfwydjKsDiPLAqF1YZgkcpSs3FwBkM94FlNKVJo4Vn
0pTxpYJqtt31doVCg2MjEXMthV+IAB6NxlWgQfovS7Pp2X9yXV76OpHtsi2D8Zpqf7KZOpwNc3+p
j2KZ3OkRIsYNa+/C9qQD7uFzQk7TAIkZQ35MYJfKFRh0Qp9KLcLuBFPtn3BmPeWYDmF3thNOIZ/x
GWLbS5fEYR2M3roE8YCBiEFmNSZsTMCW2ENAutiqWMtc+/Z3v7ODp2uSGMFYiTc6vKXTWLJRhoM2
DE69UWE+ZRAxt5zxrA/8yRY8QAKW7OunIUcSP8vfFejkkU3ubtLP5kJnvQs25KwKHlkvVEx2RYK4
oo5ggeYJXRhTYObczcYUgxkMsA2QGMktCaGN+BMQlDG9JETLPDWQpJukwxRqBEmXqW3hC4oS9gcs
RadKRpPC05V+xXD8y4Rktm6heomf325xjlf6HYW/7rVIAHKm8AB3KRIwpt8yFFByhbmHlm7qIXzc
F4P4wUfDykOgxz8QL6vAWtSpCJvQBsmTNrUcpZJw5LoCmlUbjbY6aYqRtRLcpVJefavCPPzPiZug
G+Qeq0GHzZ/DCWygOZy2dS8ur89SOkXjvBHV+GMGkLSK3vkpQCnPKGtVj+RhilJUAewuWrP+tb80
aiIw8cdLddX4GUF2tH1EqDhKUAW9RrsGotRDEtoaDSGBkzXTlJI72fjpbbIGB16U7SxrZIh9uX+O
6Nh5IirJ7O4d8fcNCBs2SjVA09r5rGLbQ1GNO0f7NnDyzBy9c2bk54Rujmlqrr/IF1Rw4pyZ0HDu
t7iNYojpm2/CjtySLKusmBuR9ftfJBCcFUwfhNZWlZ9wyrmAW4LaePGQN0UF1AAFdR8em4jT12xY
50yTFe4j3doW1A7GNbJcI2veiEBiDgL3nH0WDvzpKkDnXdbfnzzl3RdmTZXSsQjQC7i7rf5cwZd4
uz+jJQsQPlMen8MYQxAcg5Z8SiQBCyakE9Emhm2azgA0NUVINmTOGJeJpGcGEwhaiM27y5SkaCxn
NUQwQMqensVPAp4Cn6NIxCPS8cxzxsEgxAr9Hle358Wvblv6FMJOvU5V6GFZW53wXze44eFNO+9X
cANsf1TdR7eX+lnMnAZWCu5z8FkyIyH576KLlkYoYXOqYQ1OPDdrN/qvaqtKfMSF9gnE028zcaeH
SZVZhjM0AwY98l8E11VpMnWvB+7NLngskuPU7aT3LpAwLCE6Yrob1zSed5FyPlLFF9lnxhvdPidt
+L8iXmZhhbqy253bN8XiKZyHiExLuQ1xR9HMb9PcJ98OCkOaoesVobP1ouaUtZkyAqFp7qSlvuUd
lSWUmFnSuS1T/WOihcFbZqbZL49HZQF3tcgbuy/6UbozYCJ7e2UjhX9iuUP7NZtxuoKw1wYnMMga
wa6saBHw/22F8UI9t9ckDnAgzquZPXEpc3KvT25MENKk2SJgJRDoxvFMVb5j8gUg09j7Zg9M/VpQ
j6TbVGxOnGkcRbEwC2yDJJUmG1t5az1EpKKfsQj293aGafyy2aAlduxUfGHC0JNJA516//+DCgVH
3sHOhhcbX1nUliVbC/ZK+p1WiTtN3clQyc7kywfgT6sz8uvBF1Mr180AcWokPJNRH8AB2TF4/TnA
cfZx7gw/oFQzNSfg+ixMNEnRaEJZkNFVT648OPZ+oVu2f2HXLJ67sDCKAjeLHLbxdeIhCjo+qbdJ
nCNPlNMVUB+l13x+H1paQy0aSc9kQOR2L+FzHzKm8NbfEadayh46NBBpXo3BI3fQNkepl6+CST4N
EDs//YRz7eKYqVq7skGjW38tAK305vb5BMwj1vvpSxmlNRGSJdyFVIsy9IdvfqCuONucphkKcSN/
7OlD2BBOaqb6hdRxlDGRoKEWuwIB0plf8myrbtGHMnmwUPvMlY7h/g3lLRIxj9fGSynWC5p81CJO
S6/cor57st8wFRBMV6ZBcsyi9xc8N128gWO7fl84PpH9zvi8mEyOFhkgKHmdccP+7EtTF0aMh4gU
H/KSOnwd1OMGRi38wViq9gQNXf3qTMwvyE779wEPlf53agA/qr5UFDgKAzWIhNIW8pi1RKG5eyWr
YpdkT+MuLsiVAen/BtttZt2xxR/K4ldBClX51iLjCAxo7UtALVCOywMEvrWIAvsDZjWZBrMLCecH
rpYgGy/hwdgLX9+4ji38sScqpysFKNolVAGGO0/iIjL7IeLcTsRP68IFsF6A/4EAcK9xkzeKt7YD
h7bAbG/v1F4KbKpS+jTSGz3XVrURqzFc3rcRGzmsrWHhWgUH0fyP6N6jJm7RddBgKnboZQrvRZBC
E+RVrn8GekfJyB1o+qqOus91IqjhXY+1N/IYJ/Q9ceR6Oac5bN6qXtlgKMVGshycwHgJVzs/p3Aj
OEb3IQ5eWrjka23V7IgbDYcqaKVkOlO8+YfNnWmV+78/RnvYsg6JxaE7upk87VESu+IbRtH5k+2A
U4qieVeQoLTHurT6Br0aKA6FD9lqLic7cr18G1XNRw/VM5y2cGuf556FvHFA6PND7QXdsIhHBeBa
XcCDGxcxcFz138im7AX0o7AsyYm0e/6tsDAa7acw5cyZ79IDPykNkCNvjDJFJwTl6H+DMMvv7tft
Eqb799FVvvgDpy2JDZhsplsxsV/GN6dOA/86SV90Zp9RIop8iJJgSSS5Nv/LsPHGi4KpVMG8qvgY
sbe5b8AyG13lhs7g+/0ZOxmVz69CJ0viLbD1McxucVhYapA2BZCSZmvJITEGf49XLu2qu+iy7CnK
/cQVpEcgilcJBy3eC0LtVsVA/aJZBTmltAL6OuNR7YlfwoCtGKeBDn1LeFG4cUrBR2NWHm6x8fV/
ZMuhtofDGc7la/BZK97LVewVbesj3gI+PQP7mVvT+pof+k6YPMJyu8eXQX3QjklqHsjcEsK5+Mbm
mxk6k163JurL+17F04baNUtwB7J6SMiPTe+luV8dDdtBFISnHnc4AqRm3l2LVzShKmjgBbo2rlm3
mjTcFeqBaTijqg57O3Jgvtg2p94Q4vphhvXEuomL4plrSaeyoPK7EzHVkTn8TFsuZNC+kcbNh6uJ
upPv8fb9wNe9JVenh3Vpt44ZRFq4PTyJ6cdpYCPnknKX1Ylv2Y2eDK4BxD6ykvb0tkvaHhFABPel
PvM50WUtAV7uaw+9GwcsIA2u4kvbPyLY75Fj/4TMrYUdM4lFGlVZLVKOrSgyHA4Y1ZXbXnxo+7pS
KTGVWPNTrEX8/sfE/GKfMcErhL05HHdEDWVk27zd2zOUZCm+Yavsy6KhBquk8AKmPyTRjKwHcSMk
eB2QF7eY3wiWZoJJfNOIjiXFw6+FERlMKB378Pm1QCgxx67045y1bT4BoHGqficwkYgjmuZBEkNu
FXynrN2q1MhmZOgLa5OKu3wgXnzCOW8qO0DV3tt9ttpIRDjP9Kn58sfKljB9z95l7HKTvqXqANvq
La4YSEFpa83XhLus8caKpYA8MYd93g/b4mAxLXl7w8ODVL+cp+0VJgRAI3MCcTsr2UfgTjeGjDqT
G+WiRqWpvMApRlRi6S+6R49xYQzHkAyIbYfxUnUyHG3reXVBq+DUIYS+D4nkD4sckSB+wWkWA+V4
ZPwx026zG9JPosdPofMuEBkrVnTRznUNG5/Dun/gKUTYtIoj8xaC9QZUIJMANd5FbfnaPgTry4E8
T8kBpXsg5bM1m9CyrJPEF2oKhRLyQ2Wd/LflcqDG8d/aO7j1QfI1Y5Sy5rra/XIvnKfI/joCgbDt
KlLQH2t5dCyYwWFslWSVNxvz5yZdKuLLjb5XDhvLV/anFeuRxqERPf398+Zjfzm9/KL75p4ZaLmd
AIM1pIFfwewuaGGpJTMXTndMl4/YwTvJmSjijXOLFtM6k/GcbbcxwsEE2nveJSstV5KgHaW3KgvE
gMoxC0ozpqajY1LqqqTEL9j/evXWJlyh11u8Zb8K76mem+lc9LQc1zmMw65h5EVAl595tjhoM+nd
NFcoTvMd0BO+9VbMsEmBrCDyMnWQ04ddcDyfJopMsWjjBhmeuiE5oklfV51Qjij4/LFf7qrrhdJo
+QT15IiOUEoA7hrO/l5T0kWUELO3WkbqWkKpO3xUt0kA0ZoVj6HyeLPR63URN3g/YbfuCO8C/cl2
s4m2IzJvrDCohi0tR8TOBfOQ7v+TCV4xfmN2qZivPWzO6v/y5YJR2IvkceVUBcybJVgwpxwI7Zc5
QX6C4aPIYtSS81ECUNGuAU3BZbjO2n365CU8hBroDquANUhvpqZII5yMaBIM0FKiEHz9hvqVDc/3
UwTZ9sF1uSyW3cHC5zrCEF4okrpSpu6pXS/b7hSXIgBo3eAH90nTdWQQ/L3vLeXth7sYvUKX2ytW
AGi1q98a3KM2fZSGF8EK9u4EunjPGsOwg6MMId3vgU2zebHJX0R16q5gcD9rIWTJZ5THFoiFTR4v
EGdGJp6x/H6bBILtOx5hKbdBJCFbM70hHFTABQaRe322Z6YGl1lAWaZ7LjBbQIoF2xkqqQUURHRz
U+atWevc//uKPZ5h5XS/wRLbkwEnabQbLO/MMbDUMEzgSiP13zNKcTtYTv2ngxwgMmZZS4rTbjdx
3RqNEw+onJX+dVzBC2dy2r67ORhhEJeSycfNdVDVonlIwa0czNmxBZt7x5/+roae/IYkVHFvTaem
zI2X6A+5q5pI/JuiohI6L+kQguFXiu3fkw8+6ju/91CKVHqpUNjrVIQhrbFMqIGBBmJmSimJYi4s
ColrzjxYR+FoLbX+pNMbQw7hMPLQBGVKbJROa06CyXji13wWD+MSahKNHMp9he+CHVcHPWIM8Luv
bZLwTFT3Pi01QjVNKMcGgczu7OMnQba7T74vu6Y6UHiywc7Gf4b7dWqRnfnazMw0bqcNDrRA7CBa
V81FhB555nZnH/c0ve0sJXZKkJw+s2oSNdGLXqE9KIHpEXd7c9FnY42iuYQ6O9nO+kAD2Li5nu8S
8Af8zgCGQ4q1BoxiU8RghWbzNCIQOPc0ANjtI/BgMgJ/n/K275Mx49Z36r0EfqPlCHB4TH5fcWDS
FL2TIcEgi9ZjcgzdKX/lw563VP9NE9J7ZgruN4/xJinEM0P1AhJmSaqzD8v+t8QuE3jnWIHZh/fn
igyri233W8bJtFuussJ3nPLc9bZexvOjcpg12eMWX8ajdMM5TPUGOGGUP9oge4YueDcUzt2d5YUe
m4NIdImqnej2rqpAFAcDg8wsMIFxw5IJISIJ00DZACAopJIQbLsEgIFxuBDHGMpy2yNNYyGuYf9N
QmqgZnQLsEwoN/zfSQGASi3bbe51Hf3RLM0WC8a1j8KsMT+t8iVDrKkIYMP2z1oxy6+yEmzY/hmI
Ui1o51E9/5z44lfhCoW5wpRfnDQ+kN6WSdd4EsY6UMh6y7Lj8G+wQZk9v601MySKCYgd/BVr6eny
TloGDyFsfMKTTzmnX/cuKUdp3hKiV3kH0z4Ffy/R7OlcBuI/ABiQ4nE9jy7TY3K05WSMV61Elfc4
v8ZPHxOTRGoyNEdVFHe5ZyvjnjbJVM2s2UKOXmX2TVLUSYbSyCq+2VU7OsrlIDAkb7dhkcw2zA84
VgGNkX424lQp5OWal+p95zgzAXgAdlyWisg661wUAhzSLT+m5d+DZZOMoYXWL7F9DL8dw8lkH8Jl
jo8mOrOHf7DOKwwfmqU5fmU6xDrbnOb+a63abqOKoo7TyADuLSHUQ7a6YEBx4rnPcG3d7pp55sl0
cho78k6W/F3aBuz1Y2/3bqzUvzSxYxUhXWzafWc4GVZA17hQyI/B1QRk8Mh0A+fb9q+2sIQppPcU
ybx81B7yaHKUBgaZMMKiNz4DCQBEdTDVac83i9PkPfLcPHGPidiD0R4UVRBw9lkK5n5LVc6fx5OE
nzuj01WFWe20JGULdWqOCADR+juVDcwcbt92Y/YC+K90msWd/XanL9iFuqVkGYc/GgM8MjX1FVOu
oIwlDwdg+qXV6c6+BUCU7CZaZjZnwSoF2CGjkDEODds7a1vRNTCx4TNaeQlqukUhJUABkEj1+PEH
ZggCElebuAuDtalQxeU/YWW9K+Gxf9zFNixHIP5roxuPN3Lo8fvqGu49pxJ5N+IIoWjLrl+IDyV8
mZ9erIfnVsg8ILQUjoV4oR4YQMEZQKED1uZ1De7wqlmw9ZvBjkbkMW1jK8E/QPBF1UahoKCB/0kT
N4/aIbtPp9FsvScFL80SSrLZe/l9L0EdMB3t8by8FQnyWODIokzB44lljC/zWZyVR/r7oPDrX556
4e11KB39aSdkA5AfnzJUjtkXjN04jom09UkBUFSueNkKQ1ms/Pr2Ew4HGJXg/YX7VpmTKxSEMhj1
Lizz78NomDywsCERwCuHPKnERfOss4X+pXoCrBOK2uOvyQKKzeWNP4/O1Qg7tTZ/Dy9CjUWIJXA5
lH5yAy20c41g0f5qOvo3FDw9w+q6Bu5/2Cbp6nQIw1GfSbHSfHa6wmOY8he/MqKc3D9lseATgowu
ddbKCxGb+so4aGNNbfxmseWmvhN33uLfaAO3rnvEsy1wZkaCh0Em0DXK+cpzMnDsLmwfpmop2pq4
ZIUUuKRn+wvIC9AyDYjWHYL9rxpbrFJsJEa6fGA9jSUHV7sZc/FCMfYUNa64Bhw8322zh8oIEo2d
MylgiGZw+qT/28NakV75BtweVA2gPy/zGhD0UZaV/reuQ9mUFMhgRrp7RxcLSts7vN/XM9+dqOvh
nu9hlpwHhnu9wV6TlWRLNra0H+77CLfbxEwyg6KeLBgDTW5+VejYdLAzU+ip/fc9RztTIKDDjh7R
RsSP5W/GkG84OzageWdUH0GUxgtyp8vB6wiHOUW/v/ZbrTGNSejJe0SWNmJLr3+eMcDnET7yTCBt
OTQPi7q5AkntyHoSE9I7xJzUBV1K3YvLXdefj0eEhYT2IQ2SRKXGWrdj9MyKMhp8qak3Sp0mDsIh
oxAh7qmY02FehhiZml2RelUEdhm+u/BW4y71bna4JUwwDiMhW/IUyF08NUetSvxRIXIvQE66hlIa
Anv81ytyHsTo8wIq4jffQbn3bl0B2B0u5Ey16fZLcBl21442GNTUbE9hiReO4QCnwFflXg67PjsL
SVLELVYasNf7g+Xf81fBaYKSmyD2RJCCXmCsVl8DUvMptAYA/NxMSl4ceet1V4t/lKTn8djhCDMc
JfKllnSZxn1ij4LIdr6ehQ8vpPvC9TvfnRs/VRZcaGkJ9TZT0tTXDtI58bGDyZZRAsm2AdAckKZy
Q8DCVmXJjC4+dUjxoQHgTloKY97PBlp1ja9f4mnRzHQCpQP2HfRI//8/jGebd3lQdCrZuGSlLKZN
93tZDceSDsE3Y4WC3A82Q01D7ovS+aUNGb/tMBAROK1FpWAyyzghoBlK2eOiLcjynsuEtEWiHylS
Wn2HRkwK1qJVkmpvG6qVos8T5JXZX2t9hHtpiCOnJtHM9UQPx7lL7JC+8xQrzbanGRmlBZvjN7xo
FJZmNNZUJg0iduzafSXqOSmRaogvQACuSTV37r5ixOQV4ARxnO3HVB0EwZIjK/iQ0Os/5q2by/xr
3v++Ykb6FtqtCtjQViG+lRS+wEfKP9UzsF44hwTKyVIBCN5kZ9W6PN/w53FYzuv9wXPzPQKFNeKE
jdui+QA5YLjabsYTxjiS6qQaKtc0r3K+7yfZWaV3hERhyNavZsz5BHrBLlo7TgaXsWqwOjLGfJSV
q0ZVX37xIKoGmhvhk/FlrL5RUKYD888yRzGYwIE5Ufz0kzFmlSDqoPJVO7X1EEcdA3XHpY2Fgj1a
Jk0ZZFhZDzbTgtxIZkUSQq0tasqMuup4spWSKW13bjXwfaYXGX1J67Qd9alrpS86gfFwJBXvhBt4
Ah+p72t+ITEGmpq2jRDo5+1TikIfI0Mkjt3lpCAzFZKGEoIcIJS3eFsneFM9KGuLI/2oFkAq6F1X
rsGvlzebwWwvepGBv4QrGwIkodACDBHc0vVr7oaBmqhvwjSgEVhNreF/4vNOmDzqtP5xgKzvdTQr
lNfXWUVPxiqB8Ikja7PHE0VmGOpBF2mRGFXni1ExQs6M2YR+GIszEuLgUpxLcQBvUF+Yrg3KCyCt
OlCYQifatOmfVyEzrXTed1gMrngtjfomYIf2X2Kw0xyUb5qkvHIDK059tKAGf4t4j9d6JViUNfcS
vEfldvYqvtYFO7EPfDsymm0UW7J/kLTEJTXMUfSEywHOb2+gIj891juj+GCwedpzkHp62//jjgUg
/T+Qd0NcyT9YXbtRDZSLvxau2E8uIrrb/1eRxuIxsgiQu3DcR0Ge4c06mlNToXi1iFlEFMLA47VD
iMG2w+G7SM8mrSc5NRbaU48gbeso4J3yKX3LC3Hm81YSqKtkg8JWb2UYm6ObsBfFn4TSKnuGCNnB
HhBW3LPQt0JPnALE+wsHmFrAD7SN+ShNOzuQKYEGQaGzbsM5i4ySO0CdyqsUirZcrkioBH0+81B1
wLwtZcihDoQgDtiYDlH5w0Dh7+DWpMrtxrG00Z/9xOwmOGFt/sZ/PxkmBrPIYMC7CuI4FJlwdPAQ
I1+cxw+cbVBqHLKyxCZIHHcxCmdOkcKa2Q0UPg+3KqdsgfLtSoNhrNnn1Q0Ve6qxsF28q6H3m9sT
iVV2IcwKLEc7e/oDmexmtCuvtfcLsSmOa2FwbN6u/k69cjROTjABneW804Thx/npw/F/V9bJSqD6
Yi8cmGRKcyXwxxlfBLwEdVemrPDbZT1nvzJznvfqK+eqbmGFW26egLQhsK0J8SZhfifbvZy+bNoV
NXaV20Wum9cGYdq7TAls21Y9lW92aAQRiS5GAvOj90WYpHpH48WsMhCsJsnd0BUdrdgBlVRY4GAD
wyc+BLJ7i7llxMAvmafiim2v2lGXpna0pmMvp2OYM9BlVaR2k2Z7tKbCUemN+FFzmRlI28fS1dyq
boqyU7+L1Bk9jm5tp3j5mGJgF5ajwH65GDay6/+rlaCvpHxlxKDtwtPRU+dyoF4j9Q8VxE7vhXsL
djlysgTbn4uh8C8lbozfEXG14gLoZ8Xa/uqXfmgRYfIajeN3Ag6WP/b8I1VUg6I9CwA1+NL21i78
Q4EdWvbOUNcpi+Y0D1KGohCNeB4x6PDyHzaGySQPmCC6NSMQoyZOSPV3H5VnKlciGlOBiOIgsc4K
ZRdhKRXTU+chZ0fiXNpnc2uQ2haz/To1jnuHtxWGqQNpW62FQD1bFJGVAJwUg1Lx2ssdIcKD1Huw
In+FgebrWMySY3pMGU5KrouWFR7YElleqo49IPDeLTaoyBpGOoEOVfBS87gYQFYgaIRNN4P2Wy5y
lxS6bq5VhgM9Xcq/do7aSLTpcLDDbtKUtFbaiKg8V96uKTMOb37eS8WeZdoYJb4iQTKWDj09p+2s
FstoFwIqDa4Ci+p8X/aJIPG6PVLWn0S5rACf+46Qsd8TxzeOe9K9FX8qPOD1tghrmiObwKdWQYam
5iLQjn94f+hI2Z6MuztVvllHmwcBdD3/u+WtAmfpvEsZCHsOQCuGTdidxwdGYamcUFdkHApPea/D
KhAjcnrHfD8LREoHBhqx4ubehpWRMuzbvca0iijDjAeBVaCVM7rTnxh/+vWUaihDwn31bltEzHCz
XbodB9N34KndxOvsuVg+wpEMyeyNW1SefZLO/k2fdbOZcCdXuzTXRoITXW7SxD69xLWzVst1xpWx
S9x9KMYAib7KPM/TD80ji/NtJL6/IotPaUPwMc6YQiTTvhXZfrciLGf0UoxxhdEIRk+nHM0jlXfP
hM/qwY1jBUQ3TpUWPEfuhEBAJzq7rlA44KVdMQSxO1lJC9COe8buiGTENxbNbJT5ZCPFIKMglmBW
k1LAXv33NIRU/0DZpggAa+Vb/fIiuhnNjqZtX3OQQ3C2YI5n1ecqB8sTOu5tfZV++1bqmr+MrtsN
jLLlckLcBfVeRlz2Ru4u/DPqSAJv6QpWkP0vB9n99JolCh3HPqseq4ZrASyitqgJAG3aMiTRCUhH
asBidP/Ih+e0Qs0fevWXA9GMcjoExgbv8X4dO4uGW+QW06jizxyJhZB9UEz5a+7kbtCGWkUhbtCA
OumoN7lwQ3Tm3jfJrOT4fMySXIV0+DKocWXmYWihFzH+7+/btUBTd+hR84h5r+5B0oTH4spLDfgs
Xn5J8jnwrnV2aT+4les+LIJ7Ywht38MokswFYw8+qj2HlYVyUSI20j3uvk+RIZ6nNxaZ4v6DR7/P
XuqFxiqSJrpT7VfUbLghjkIldHW84j03rXZdCa0xOg/MOGjTq3iNdRStPBMaJx72FfMIRoI7SZew
WEeT4h5DNbU7g1U9XNL0JRFP8Iw+fG5YheiecPTuNwhJqJylMDAXl5s5MkFGhxCfWpLQXBBstGeL
i5eHlcWjxo63nRDjVUIwxMEZ0sacRUQWCMGcdUAhwlHp6Bg5QcByaFuE/JYH+WCAym55OYrNo2+T
Ske/f3Aotw3WygwdAaxUzWaZy63jG8N5wcbqB4vU/NFZ30AkkYNhKkLcrl3AClKg3WbyyV8nhLpm
luGdq4xAnvTpAyS/Y4Bvt7tQzTtB19SHZn5lasuWmWrQ3nKDXkcZAu1LNTDoLcbOblvLht/b+Jg8
x/LQetcxQ8a4OcXO+EzWqckldxYeR3xMGeikSMSaO5TBjJfS5L/KYAzLB4p8Rrww28hveBpOB/VB
8iAaFVK/TCO/8Wfl8AivsVV8OLxA0h7OPhta0nbW+Zz9bQjfP4MDtiWw3HD12AwkdMDvfCHiB+Ad
R5+wAMq8Ad6vm0RvlFvHSP8ilC2UV1t/nk+KBATvdCc9f03HjdbrNWClPJC5oNaCdS/ZfbPtuq4V
7vkBPvo2MEGPFrEVEZU0kSuL0D1Fds/rv1gHQteaoBwIhKdxSxJI8cFV1jvHJD02lPwxlid1/Y4U
fde5uE62gPtlwienIjufxJJJZGyETU2VK8CgKWTTFHUaFzhAXwMYrX+1alX9E6bALklGjR2il8kJ
+UrpjA4PJvmKMfxw/3CLoDBxYG+QRvMX/TFFQBPgDYxSti3TcCnYyquicq3xhz35zbaBHfocErwN
wMc8dFHKw8VNxpPOHO9CP0/LDM3VNzupDArKVNOxmrfz/gT7/XkeVD8po0kOuLL+uZcw6IRWgb0a
swzGYUL1SH64NYcJlYJj5Zcb4TvId0+PqWIAOx8tlzRNaMhCx3FCdIGszxCOzePROVjoiCDhBHse
7V4HNHLjV7Mw7nvUjKgk3T5hFL2XbmaNB6LCWMDDFucGd+bcqo2yOCtgfp4BVv5mM9qJtHq7cFgK
vgHsOOi86MzKIynZzar27dxsJMH9ED15bjgT+gWbiwMeLqpX4/YQbg0ZvP8zG09j5DEi5HtnKEib
/g7D8LrPKmq/ZbEWZpQpK+ue9wli1DTjmV9GCMsW6QCBN6Lv9c2/P7JQV2cIt+EjMH4NyoVGFaJ7
VBhe4ysD5NlslUAFAivsBDzasehMxvkduKeAn5+aCdJxII99gCddnSIAm1x2Y92OPWyReA/AQ0Uo
W/GC5xg4vSK/NHis2VLmd0xd+pPUa8/SGGfB+izyI1y8hrnRI8cKvPc149MhH0EQ1sh8bXddTK5j
ASSRpqYN9433yK0tpWozj7nUSCW5AzAF73eNbTseSPEfUzDCmPfDhLXmMzxorFWR6CAnrKcLVSD6
Fa1YVh+GFADky9vL/mga1kV8npZaILflVxh9fK5a1ubTYD+YGJn13Wzon1nmqk/IS4eGak+Dopnd
lGTotTPXfK4EsK0BSPj684EC+JI9kSfUq5mkGJEfxRlIBWkKR+6d8hBYCASnRqFLushneE1aR+2A
dD3QaOUiA1Va6cYoiAJpVo8XibyJlWkKkg3mnVYHg0a1l4vQbcLwT3dQVHLy0xmZpWaND/qkBLpA
FaFELHgCjIziti/3qOnS11AY6+ABI8lsdno5D/lyXwyHfmjWCSt769c8rTzdpcFmFQnbARcDEgkN
FoYwzulIw83ESUah9ABlsPj8useu3ma/TCSXi+T8VnDWaHh6gDT1CmkO4cVmYcJhItf95uoNo2F4
9ng/jj2EQqF1TToCmlT1oH3NYRKz6HPEiqDyB9+elg240hJi1qvf8F0lAstFd8eIP/E8eh3kQsiX
ZuyrIv5mcN1GwvD2gIiTw+57zwQWLUeRO1JQ6yJ8iXTCFT7YExhYtD0P5axYSVDLcG+F9CZ0UHGg
B/96iAOGEwF6NXuqg6LOKxvWhJqUFT3xbFGoORb1QcrD5eZ8rnBUkj/OnSIThXH9w/RIuTo778O7
hzrs7AtrNvSa2BVL0G4Juhg2VEFZQBvl0wG6DaVDnjVwsqTyaIgCE6HYOONIDJ0dmxTeT1KUgW3z
eUjbOnZzJORGd9WPzrH5efFMmH6wox9jOQ/hOY/owTgJa0UTXHp+Z67eKuMJqd/JcLa3fujsg1wD
TVb6AgRFKqaMUTXOmZ1wBLlDd+2BiP/P+J8wMnrCXICq3unkoSIVhYkzJfrPJl8cXmBGmq32nQyM
1mqYziEfPTwFCeDMhY1qUD20Kq2Za5TwQPlz7FQwFRN1y72n2k9jXaUU8FrD5IKsBYWR+Ol7fnOR
SBHYUEd5K/wKj4/G71wPnv27uQHnBN0f/PimH1sYotldvvMjspn8F4DlgDIe497bicpcd+bl1d6F
07SEUFeER744tGpHE2V6mWiqZ6R+ia9FMum7MuNKEojxYV/McPrbcPAV8my/z0uWOgKON0qcIH1V
Dhx0aLkMl8nFyLD2UxtWfukgAxCMrfWntNkEU9qJ0WhCQRToIjYqRfdka/odvAwuR0fEQcT0jWd/
xM2xaO3HtaAJyf3GMcXzGBn+DeNEZOG7w+vI+JKtT4tfUdsIT+hzp1pzn4CDO/DA0Lm4B95gw6Tp
WpYgBIUDvttyVD5ifvLmQfqEuvMBcL5I7sVt7I88nZliSZMBhe7L7+3bm4PsDSyVTE02u0apAO4/
HSvKZNsS8zZqkQBDiNk/dDoaA8rm4VqlO5k6wxpiXuHB7ziINkG85w+Km0tigt5hV6ZPGkD2zcjs
S9qPadJqQo/aZtJlE6Nn6iAeVIym/ijnj6TkoyYG+48wnauxqvwC7gk7QdWhNbFzxsZUB4ffIbsf
/vl0INEh6V5Vg5/w3Fr1EpNluPZLzDwQ3yOnX/wnaMQOsnotYNiMgOJn7cGUsEALQjvKILQ8dQS1
C+BtHlqXh/Tjr15Ty1nHG609hnS1IcfLH/I6H1tlboTFAmnFBqn2xcWmAXI93BWgxCP2fEBI7HA4
KcZRzETaFhTPGE3a9w8fVKl+yAk82J/DPJsQQnnmxk7rEoM/iDwnNg05AtbBqZzOlMTz2M59I6pJ
ALGNqn3tv7/UFiknsehZebYNBEV9d96+oAyHA2j2kJMV3r598rJX6iOPv8ys+xgceLr2drPDcSa0
aYlU9Bqi5BC4WkQrp1zCkgB/zEUOUbruXz+Vk5rebNMLut0hvO9GJqEgHtDQeLUOSkk9ikyYjPwp
Z3nKSTPABaLn44pciChh3FkCiDBO5P/s/X9PNT4jtwYEO2k1HJpo8WyxqRaKGY1STNCuSkOUwBZ7
8XnKkuXmF22WeQtG+KWjqB0UIeJgmUJ/VoD5bdYiDww5U2CcEvbfIn9/A9n44cMxTaSws08WtfSb
HiImPsj7Gt13yrHZr10pqfUeEHGrslaR2mYFboELmz6SRavrdXGU3wFRcCV34xbVL05nv8IfLOM1
dprgjiqD8rkKSuF1yxD6ecCOv/lwDsp07dfKkwybQS+azEvnZexZqlBNS+G8PtjjRlRCyuhZZt5B
Q2FRVidmzUt2+SzUFQIiZMe75dCsHrc0XPEIQeTEj8twPYMs43MLi8a3h0gGgJ9R1kbFgo0bXeva
lI2xBl9rWdf+GL9j30TZjgpWfvqohlnaC5/su2s+Jtrf37LhBuy5U789i8hMUAf4443XVqA2MD2B
RBpzsoJt4Y/0qnwClWFUU94tlqSd6sudp7rl8/Kek3iYvUipatijkPV4vqKgPAuFAOa6azlyzu2U
9Glo3DADLbp5Rx+z9jO3EHW+EbAOHNYHASd0kh3SUCg0e5WhueSWOywifNzXkLrpjpIH9t9cuawd
/EO0VA3djjierWY5v9m/ki6WTThgNw8IuLp9JXT5XLS7cyGMzyWFAGsQM1ZUqett2so1XmO/n0or
ftY9tmcKT6NXCOLjwK2dQU/IRXRpaf1+vt02KIoUm3r45fThvj+NLY7rJ5/WKvxo5orJBDWqaDY/
Kmsl+sr2vr8pM7vTmUKOGLUnaYmWJzjZpqK3gBwsZnvaYwLlnT+1ynj90tCXKKboWAX4L3yQpwS/
b9++IKC22nu94HjwotTmXueUfipGNzGulIwaEtLIzrltTmQdFeuIlj/4Wehr4PydssQr56s+JUhB
P72bVg6PMC8VKMwuYx2B3JZyJGenW0EkIFwbui31crtCApImjbA03FuW+kAc/uukIou2XYe4CivY
PhCzwyDkI0SDG/pcqnMrkfajd6GJYpQUHw7DyC3/D4o7GonQzoMP8PUEtaHJedfq/hDQYSdL8943
9TIrlUP66VkJXNXyNJGB8Lz0mV6KsbBZL0YrEpEtNd0UDqX5XKmiKa6LREe6BLspb5VCAIjNUB3T
wdqp+Ha0a6MHZcs5/xFGTKqJ/cc2G00tw4K5XC3znW62RIR5TTx1+kFoSgOfGCd+r51buSjxvUe2
9itxEd+2yqXXS2ENLvTIVSM73TDOvMGlZJDPWadfOlZv8wVa+Vnsvp6x4tet8ej8ACCSh9srphvx
iL+4Qjmov/anWXTIUbDNwu+oO49UidVEePDSZxu8Dj30znLKl8gFj3FIecppzEYceCDaspDQKZvc
O7H7xsX2OJekPfLWfwgh+/Xvgc9R3eD1Ac+sdcQXj1yoAEJLq19OkyUzgizZwOMv+5ytAB0HNih6
VjjjzeJV3lEKWfANg4/aYuUAeQBD8iKk0ZQFQs0OuBVgmGy8MvouY8yit/KUp7QXexYD5IL3lRnR
vMfeV1kmYebJOoycKideXa0J7DTrEdSDQ7PJa9R2xLNlClKXzS8cRPfedEZ4AKiHWK8i5N4opzTo
4a4ahgJZaW2cfOqWSlfacIAYKDj0bikBLg/BtMCOFvbqzzzu+YucqE31RMvko5MpekWD1bWtNgEc
VttahxIpkP9JJG4TbE1baC/0aPxkLMubY8uzaAEHenSCoVfTuvfwDjeqX4r6TX5xMblSENkTmVdg
2c56IVxSFn4iY/OAkrH+bwuBbrN2fzlGsZxEgTeGcRY0S37RbGHqC3HaX8seSkoIVY5OJ9ZT4B3G
KzaSgo2xCp+8WyRKEG14Vm5LB41nWP+iJJE+B3jGtJI2J3lEVEyPRPXf+lsCLwl91vRCZ7HRn9Ee
DaW3O4JdSgUF908zshaQh4b2Mwi4biW76ToqiILAy3bG04JtTFpPmEjrqVqQiS2pyNcZwerFLMkV
kAD1Tx+4HaWhjoZgMGKknQ7HOzSGS201O2A9lzMRQpLo3qjIFEmsdYJRS6NFrn9HJZh3YWgtOIXm
OGEhpdE1VNykK47hZ1jnvHStosRpm7ny2KgAr6p75UXfBsZzbD0G7y6Id4X1g4ilpukSso1SzWfL
X6fthzMNQibAMIa4rVMiESwDwcyMNn7Vufi6CFuVtDOalvV24ULq6MSn0kgPdSJihuuAaVhtxARy
mqf6amf9DVZVQfu6jGaN12deiW7C+XlasqSaWYdy3aC6kzBsDzlNbxPTM0nIuiDtlEvx/segc8gD
4edAQKoluatmIGpuWiPIr/xSzqOex/vjgSNz5/eR0WTvWzU8d2wwQwSpcFDo/Az3JXrbKiDGJerb
DJdpkgp+X3txYXq6mS6+yhRhcdn17Lgn3vo5+wMzgkxXIppOpezXEcgbcqP28ujJiXYIBm2HaoCs
AhGMHrJaWEjjeWAzwEw9zSetDdFnBoHKHDP82Fbb9RB3j79QpUcPElwR3hgjVQZaqd6kv9Cql1+Z
Og6coHEOdqVE1dHRCFE2ShIJ3ATAeBsc4djAocEBzlmm6pAAXIPEXIHhlObIhmudYyB874Poy+y+
0osY00+hAXNVj3oa9/WfTxCOKeVg7pvk6/NCw8aV9JtNr7+i7XFpYl7ti21WfO6M0Sk0hvOCq+AS
6TANCSy2+q6BhBMQ3HkFJGHqMh59L3eIICZRr/TMoX5ZyZz39EPxs0EUlYbMOg0z3FMJxlVVI3mK
aU0KLfArOwgyZFu2bXD0KtF2GFlj3TK+sD9xRxPnaMB5uVobTVJ3kMeG8HGmTd+ygjLOpg6dzXye
GF+rBeTzlarPn8Nhey6pHFzgWv3OiEaJ4f6aYf6l2K7kNGTn90cgI8NITSPV7RyK9/fGQqwBQo3h
4MxWrtpSx38VoEsTxwlOd5N0Mpra1o+eKwtfKTekrb1cI8EW1euzT10W2zG/5DYdUWGYmWhuqPpN
+sytme6rsOPFq2XhrkyRlvj8TLHaE7+i6uTYy+q5S+T5fe2YY6T6H+TmUc0rWsgA5II4XeKyYPLT
OUNpk0U9qCFMNEXjIS5ER3ZoTL1hTP8nC6JcctZci4WX77N9O+DEQwOyTf8tBh8q9ySMVSKL14DD
AwwNa4VyldeyJLrRzQeJx2vyEgZGdww1cA5z6YHkWlugAk5G+JnaojL3EeByY6Dck1BPjEm36sjB
ZHnvBmDFezLiTtZvw2Us9qUDk34EkmlbaCXUVxcA3K62BKcfTAKdTpKg6Jo6pwhkTqi2oxqGL+tz
2src2gMz1oN40MTAX1QM9y98sNCh5pN9SgxnVATN/89OBRnUXcfbKSwyYDTsv+jKczX4sLLuE1bB
uWs0Mi/4lXXM6jrafG/a2KSFGUDzp3HUTcwooFTxtm6Ic8/NSyU1P7SZYiKNb16TTS/poqVaMTsD
AywQ5FHZE7F/UCITE3oCDaoHaCcHLMsowNy/59H2AJ+Cg/HH5Di+rp3AwBi1cpNRggCoEss9QdUJ
2xQhQC2+rcTUKnlOiaw2p5sjoTViZso9RrQi/mF3REzjtl85X2UgPXOOxxofrAb6O1xN+WEgZ5Vg
vM5VUC0bRTd3X4Ms/O9q5RNCequTNjAXFR6WBjHlY4HpCGLPvsZVNQOcpnJvzeEKaEbOj1OpBS4u
mEkuvVdPc2thLLw7gQyWQgs4BNQtH+diB5vowlPf5LW5bef0VVZufhaq0EPx5+PTtlmf6soxKSXH
LHtAZzQEdR6M07qC1Czb9vvS6QVFxLZZJYWQUH8k/gnVSqAk5V5dSIJXstASs/i21t2Z/e5Dtibi
RzKiWms9ClHjeCZFfpV08VqKMOhfxZoxlPW41KaB87UwQ9Z/a6nbvUl0A+5hbJB3cdEe8HTcWj7o
xRu8IjEGPxK95YM7XHXQNGrGjfjGbhUl79s+MaKcT+OJXL2l28h46ZL1FcZ10DO5TYpdwcotjlwO
SMsIJnioCwfwtcE87nIOZcmlzOgKgdxG9uSpuJjKxj7Y+u4ameN/YizU551M+9VMCzIjN7XaNMYg
fagIPyCtAxIiUewaZFqdrMJtJOW41V+0Hzh4vBpsqxkrdP3z8cUgVpzrY0KEhi+1Vo3lNIbR6e+S
gbPw1MdvI1tK8kJjtK5J4Ldf5JaX5vUzDtGdTlASfxkVrGgh5wyfHxjPgEwn3LmeKiM87sK1lKH8
va4lH85dViCe3fcufPdlsNumYQvSpwLxJoqiEvJKAuyB2TqdiUPahCniQ3GJOlt2GNi0Qhjk3T/t
De9BcPtDV92IrD47Xu4k9FQ9D3Of3fopFfmH7pXCPHa0M/P8IFuWhnxz22OtLp9VJlnvF0yWlVSM
gJjKZ0kLjKK0YU8k9eCfzGmk1vAUrrPejp3FQaXhdEeTpX2n1qXzNbyisn3jI/IvmSuKMk4HqhHa
IVfDxjc3yZM8z8jswS3uxR9fONKZBJkKbQDS1ydlDu8s3l03QJF4zC3u6QZjimEr6Q+LwfRmFQ5p
ih9rJk4bT8FtUIaqGoFjG7wB/4A6wMEUxjwOzQMKjZouEFPt/KKnO51KABY+lziIXGhwj4dypbQL
EJpT1iKasnM+A/kcALYWQjgGOtaZBNMT8yW48jmNkp+D0NUANNhi8txa7o+/B0zmkrJN6JXVS3ZI
VHsCyZZ7WhGOLJSmFVz1n64sbyN1U+XKMYLj36DgMJ6JqY7gn0l83cU20IPanphbHcPx9UHHrG8s
1Fv+vKqvMTTL8X8gC4wbghRJ51ZBEQnHVKXJ0kU2CcFlp2Rid3ns4KoQEfkRYgWBBHDB6snGWvUk
1uwIfOyCPYWkdSgzmqRaE8UFmTTkbz/mDPrp7iGbneUdlAeP4OWXlCGnlLWc4zKc5oGy7A3kz8dN
AHRsuWkHrcu+6aNRp/aDYPN7KKWw/onKOijb7ze4mu6MbT1xwr/LsSigCCTMyPYvm40nhCpKng2S
uWTiBTDP+PACjrDguyGp2F8f2FWq1r9DqktwzORr8++YeI/U90V7P81iFVF32C/sTIg8jJpyBrVl
7AOsFjCsnwcWJA5v7oAURM2+nPj4vGBqOW0rcbNxjMB/UjElmTtwtHgn1fKn53ErIwnegk1RofeF
haTGy/9T++MS0db/vQvWXUHBYTAoPACwxnLdaaV6CjrdAsiGc5qX5uluboEYoscT4BZKau3rw23x
UF5fMIlFb0vh7myAb+qCkmtiX93XDS1gfNjvyb2mZeBuKIGsSTAIY9WWnJpSV+SOXcWvrO5ib57b
CNG8XhdMZ4t79byDCaybU/1XurBeWDELVF3J08TVWQ9QsNlOPab48OMigOleaHvuMmR4G0x3VcKW
wyfH5n86cZXGdmxH/VKPyXwSeYHNLFGrTo4x7ByIrut8UKQBDJviuR1GydL7g+qhXt4VwT8yt+XV
Nj+siPMx/RXUutgyZDFFwLTk82KX7Q9MMmET4i3wyCw4I0YdcPndAaBRSwfd24nft+2UzdWZNhfm
xzuNLkiektggOIyrSaLBKwG9MP8Ko9+wMKDxAD0i+w+AlfgEHUtOT+d02hkIM1dWG+1aPohynlrb
Vxqe+kN/o84CgV1L3r6Xj8BGedQt11hpL5psjO4CMYareJQ4ttd3jhl5ho6uIS/w0V4Ixyf2rQMO
zZsVyjQVTHzBcWCt0AGH9PfhqNktk9w98cgmRtLyZnDgfzA4msvDAX3RSUwvT9ABjtc+H9jAEN64
lSPXu5BjASqSAaX/agrRxcEiMmgxTe7NvB2/EH3zlnmfqwt3VYDGipZFHuPw/oWMzL3uW6Yj30gq
NZWGhcEXpl600tGECDo4B/mnjgASBMQ+mBxhFL60Hdsg8B9HtjKOhyAI1FGh5Jh9qVptuYHH5ZaN
HAyaoGZqwaxJR4Pq29tRIj8zXLuDco8PJqqPc2l8CgJlMkYyz0wBq8GIMTr31HeS7JRTDWsjXISN
8v4NF4wexNjOZI8cRC5HMzbzY+s6KH5oN46on1g4Xig/21r17hDBnzqZN45UAEE1hKBmZU8zMtDs
+X+wsHAcmI1pAMvP9sxUR/gt8EmUZ5BpasmlMI35a/n+Eih7UjPOtBXaErbjMLjy27i47xSOV3sX
owhDWZksQVgTmSNSBthQlGFbstkiySxc77CeDWmVWvkG3tj6c5vPanNL31szV2V7MAA/39JF+0S9
AvuLneVH1HAHCOpHi37Ioq+AZO7DxGfzcHrSwytbrlOz8SiSiYIqa2365Pv8+XBELy58amfGuii+
zvAwvCj6eLW8/4j12wK9ddRVsIoVlRBqDR/++OF7cR2lAJg7N9+/nc8ZjtqSnwRJW6r1puvFHoaD
Iff9ftM76jfqnui7F1mQgH5d2B8AxCHlzh0qlzxROgObdTq05REcxb367/Q6Fdnkfb+EkJD1fdeM
ryuXAesTnIUvJPGS6f+8NgLika69yz1h8ppTHDCBJIxW0DikwfTaAJEX4hzQv1TM2l0f9/eRWKHQ
pXCD1eJOhhZ9zlTpNvtiAJUzpGSO9Fx/kJdttRTXhd+3uXiqFdYQLM7g7A/ZDadet0ruOUiWTzye
selQ6Vf/lBz7Z/emglHK73oe0+gtioLzZFVG59xhbR1zcUVF2djWyU2oa7B3sDZx4p/vWNOUTRlJ
5EjdThS6B/tjSGaHc55ZXyTSv2uKV7VP1PWuOpq8SKQuIY8evZnbevGEfurbWygQ/rWNEJ7Vqfdl
Zdne1TNI4k6/Fwa7FjHiQXisLrVaiClDJjHByz5XA/H1+jeTmW7QZU13Mm6f6mrOCMIjVrvSRTyF
fj0FYBwbkHa5noObHJE8gf18yRhDSWN5qLVXI46hKYFkjYd/eaJY+f35hc+ZJdIiZvp/dmfv1I4y
j36WE6BIyZeQBzoNdB7rTT+WgHIxpHCEhXteHxVka+fvr9162U3LRWLHz/Z4C7XEzaUno2vXLvDG
v7WgkGG9V0dwfc2ftSr7DAOUVcFcMhMZMXY/v9bH5+VOedVUQnVJMwnULB0Dfbl3+b6xwyP9dDiF
3owzDICHLLYUIqUVEpbMw4lXv4pe7jdJiNK4UWqtDLiF7UZfcDKB2J7JbsA63oqkxlWgXgV3EsrD
U53YIC2ImW+vhYT8VdDUatXfUsI24e0MVGRKBFS+uYeRcciyBOsmFlll0pGNGY1sm4OZUifUk/oT
vyYQia7i8814CZeZrK4f2E2RQuhUpLL3fwAbg0zUIvONr2DTfcN7SShgHwqBxLggpLJnDc9rAWcN
NcAKiP+L02AQag6ei8WBzt+CUeS3yoW5AEZxHr4CiCw8c+Xx9oHpItp7kCmrDy3jN8lsLcbrMXHv
u6PHnkZ6bHwxHm6Ha6MXvISpa+gOiCX5RaigE8OWhFcU24kCQIPygQYxZjTBVPiyl50nh5dOeHB8
LsAXRAMO2YHAYKHNg6lZCMLxnF5+VzpB4FJ5OGo/fwOsiits42vLU977i72B3q9yv2qKGq2PLoad
DiTwbcNgNcekQ/6q4jOWRXufbLw3XhHcGvuvF+zCo6QxhLgCBIKWYd3L44+IviHmd0eWQ3WZxRp3
/ue3VEzIQfdkocdH87GLcQpv/G8iCNiQgMSh0knRvGLXGIblRGyQQLK7vkoj6yKMqVM0YkJ4JOm6
qBkeSZ2lC7UM3a1kHaXlsuKGhG7KTyhvSdQ5Kg2XSHiBXn0lWqHZ8c1BS32qr4KyBFP5M+Hc91L2
atMOK7Jz+e3EojWPhtJ9sxkkdNnUjNID1P2tWcUkzjXAmVfadgmL+NYCxUJuAXIzXMJRXWwIRZiI
01ECHh7+bXMIzJQBZDuHH6+OCI6EEJaExPuxLgyMJ5BNf0HvKZ22zTINp790K6/O4THBC+m6TESY
7GcN3FEY+HZh3XB5sO+2SyqsGUwjoR7j9ZrvpZUdM88WTGhUwHEuGJOxDZs+AstwVtotkyuLfggY
SxSlBwMjM3XIU7wxSKrn4Zmsk/hqmQryLZTQTEZMNTRaErEXQZV48ACEL+yzuO9geXDzjL+gTmEQ
vpwB/6M7uE+vgnM0Qo8FDeo9djJLzXrOUP8ZQzjWQUx45jYrFIxyqUrc0f+wGw1oBkSTjjL6P2yT
tDbAv22baArWIfLzsBIIgeVqZh+jjENJ0gqQTFREN3jRjJKe+cCHRXsOwRBevdrkGBS4vtZXr2jY
M+UmSb+mJLPXN4RYyfumhPPX8hzGEineoKaJ9LyfXwu/as+mwK7jNGAqtYsho82QR4+MGJq9Mzmi
2ktqdBdnbGhjwRgfdF/b4Azm612j2jAWR/RSkn652VMnFAPOVNtV6aUpfyiVMtVrYaJ0bA+YBo4M
z2SnZPn6+sON7RAfaBo2vhnHpEsKD+eAA7+leQP5aIcdbn0Dp36SC9lNmX1p0s+nxUFHi6fAP5ow
M4LOUW9UBHSN0ouUJyYO6xQzgARak2tm6ioKve8mp4sx41txxOfj1cYrgdgaKzpa47yGZYaOoItl
Q32o+kdjMA3mI1Lzj6L/dRKvfRwLa6LD2TZN4edarX/TE921YXZcdb4e4hWw497NiFjkghI0vItP
jJaCH11BZtcZvzbeg5aYBZuRoijjmKSIPFeRtKiMJ0qq/BzJy5WXrOdL1LJ8IoODSbI5w3sBlc2j
L8E0ty9/4oVUhJqrVkvJJdPLuKrBuqGEuVIDXCG2pkL2W5LGAkXPuz5VZqp2sAaendZQ/QL3Hg+a
Rr3fA0EvxIB8QvTTe4LzawoPzh1UU8LLi6ldHFsQkYlLgV+irPOZXooHjTwY+x49psmxrY0mkkIO
JwQUKeT0uoTYN2XLe0c/t8Ww2c2wVNqqzby9BS8SB40sDRdH+J3Zkq0tgrbP6vEunz9H10bWTpit
Ffl4gVCiEOwgXGMV1/4u0RIFCFG6O9eIQ3jiNa+lNyD1p1KH5qS1FIakksa7ETwf7t9BTrVovmHa
RAgSjdVSCFBCwh/BfnMtpipzdtuQUMCZShn3Glxr46Nnhp9puWrQvvr6a2uzNzpW6afKDy9WHWi1
qO0LhOWaM6Q+u1fcuwDB6IKwtzvsqMobJJlkK/m6wtNnf2aM6Kdyl1fI0YAye52dek3/T5tyskuu
yU5QqKm9wm2aGtyP6pniPDOb4BJru3eMPaNxIQHOR0izX5xiJPiB4Mlo6p7FiUsv9/frbEOViyeL
IA4PkQwZt+1aFeyq3Kyhj0vXh2Pw6hO/hjDSb8oGrs3FbLPlQ9XHew3qz3gW2ygsmfYjhYud8D8o
fs3JhyQavIbhShGLquPcPHBb93oHgbD37gBtOpdD/jPk5CRl7f9vee9feVNyqFkpHQzV++sBEmai
t6Me0Mto3PkFZoTxL4WpmGZcKS7qFZQU/BRwnjvr2juZ1+xesl5vd+ibzW+nvb/N7RiQNRcrmho1
dHEgyZ/HfjjhsHMdxRhj+saeiUqG6WAwq/o2ESbi/9Zx+RF7Pa0W4APTPAQvb1954vFdizlUL3Y8
B4DGlEiZVuI+v4QnYQXohgupQE/7xHS3W+iuMgiKZ75ziL5xrYI9fPu+SMIL+OMgMuIdr0v0e5+e
KfOQ0xZUBZ/kPSAGE7OZQIfocB7IZ8XY5XjDF/fukTkUbPg32IHwHwxkK6Y3FKlbaKdSfHgwLC0I
+NNQus8CEZtEcU18BmRTnkupphudJXDPNyfIZn9DOt2Se+B0mOHHML6/+AcGBkxduqVRY8FoclSg
1LFLegY6zkUVfaCeMA1ckO82Jx+J0Tg1ul0bRmhejEWflxBMPi9FH8MDNLU63MtL5maYYJ9pYQMB
GGaHod7AwIJ3NIMyU0y7yxJQfY2a2SuspKrk+NOIvG0NbAH7JQPcfzC7XemKTb6XMTNELSxljkCC
d4ZNkxo2f63fTCz/RJWzYlvpqqlflZzK3or4krYdTNAAnOIGxtvAiuV5GfrJBzMz2rW8CggTbFDY
fyCbt0hg2ie4SgSMubBt/eZyvHh2j1/AociQuOeR6kW6pm6YoOSqRkBCamTPo0qaQ2eo87/RS+fv
KqfADuewITfpHjbSf9iI7aBhAABKjpzILkA9iUdRdqQaBf2dpZcvrN8JZT35eEpx9Km8KYfCm+Pi
soRtq/QLmX4hnAdnXyre2akw60SwjNLF1VU9WASFlZ40Int+MVb5NWgQ7SbdbuR5SIaOGxi3F+g6
n6lqzJMjUtJxL1kDIjGFlWn8gdvvSnBwXhUmru7SWGvwcWmJpKEOw24JpmzVQcSsVi4ELwiSLbnd
kthQoVNu5jT5CgqJNFzprm+kuuuLerey1pPiXrn/Upj9DRh0w5bcxFYCJpCfRmpLrpZX9oVKoKpC
BQvKOf3C5hWJt641xPH6VzKb54Q17UJeJqh/lyO3tn5CXlNeF4R0pz5xdMjCJNmjHDg4heQ3oKVc
Tu0HJRfeAgSpN7rmP3DpXh6Gm/OdkBAgbmL22ynw8q2TYWOBfz2vpyXDlHeUtWvF2Zhkr7LQna0u
dxjuz1o7qBB/rUKoEkjhvT/q8yMFYvSPiNEGhlrxI4Y2yfDlZMrImF1ovFuLnvCtFMHYcxm4XR67
acpgEiuKY2C957fdgxalV7wT9NmBO3so8SR/GNNq3J2vgGH5DZ0uejEi+qaq3pCuj7GZ5qB3Degn
dI1DaffKQPtCyZ9ZJNGkbMIDjdZUcaB8DbhoVLArPZsamcMvm4lSHA4QabWE2VLB4vYqBYYujx8+
796wg0k8PNj0ze4uICuoR94iXzqALhbhhd3/Q6deTJUOzLlySrh8hN3QTeVV0K1uqHrzH98un9ni
fZaZPmVSjPSTurhaSwnm6PMCP7j1AuQ5UEDdDI9oV1CO/axufiglH5haLxheON7Q/ggHNkzcYRfd
TMJSROfsrlHnQzb7JDHCc2qWXFZiRoSufz4RiINte2lACl/SpPV5gxRk4PLZ7tOhNKDRbuxaBhSv
S+FYaj5qSE6wgcNG57O7E7D5oSVKjGhhODquRYcsgFu7TwOlop/d23HlJI3sAAxN5VzNIEQXCCfQ
J0eZ3/xFWNka40LTvCYuwP7Y53GboOhAjIl2zDqvrmhXqUJ/mdjxPCnDqR786ZQgiVlhy2N8bw3V
80SgPKVgTKgV12ptyKVXuJGtwDc1Qm3VfjnxtAvGUyfx8Jjze9gHosskACPGjI27FqDfrlWVrwB8
dzQmCsDRQqIqpgjHbDbRwIbzDPWEOqrRDoJHovFqa2jebkefshiO2PnB24HsCoIRh0RTljCv8x4+
XjA9GkbNuyF2RE7zM8NeA7dInRJL2QDY/BU+fo0y4i0tznaIiF4au/ZKPuNsMh0OMeGdiUOTxefw
dzhX6xlYsCo5i0jNVcs0DwBEfPL9brQtScReQlrhSOu5eRPX6N5B2N8u992VfS8JpduNXZCX9gVf
2020r+iSIRR1+0EfHQpnCWIIwdz8sPEGd/LoybablLhJ0KAh/gNvJblrJ8hfleqs/IycX7SLizPh
AechZ2TrODNadconsnKb5usf0kr+JXuKVafNbrneKka3UkrM066J6D48F3IcxoiwdAPV2umjwA61
PtIyOkWnUZPX0aQoAFBpwzGIAna3vlQaxa3BL3VFUffV45qUKn4W83yiYRWnFjgBz/14kn4klwYy
X0iCz3I81Z0ZGIgJN5OcFn7z6Aclg9gpTRnPgE1hRUZFN+QZEAwYp6xA9QTdZHQ9RJbFnEAXLEZJ
bojwfozowsW5xmxE8Y3w/4glUYZCQeZn3o5NWzdtFy2q0RLYvcuQf7k/Y1Eh5pM2Vm3EOPb2EcGF
ZN7icwd5ohQr41oHx8tHWZvT6ucsZmspd1C8i3JbJLPcDvpBXlSp/Otjr0N75FFbmiRs34uMt4ly
BgyshiDM8dGkjQubIfGHpkE5KCgnkDWRAP7lcOTj1ebsxq+eN0hNoMw0Tpa0DPV8+18WllNbuz+7
H4Jc3/VHOmXZYAdSdbo7MoMbeham/GH8UKqTHTdxaY0eEKp1ANxCBZJIlGrcTzDwvj93CkZSHqM5
02ILGChzMs46B4bHtl2JHiz/4oM7Ho2WSA8R5PM3GGDtxLH6xHYSAf16jmjFVHOxpEQVQdxJz+pW
uIAvnMo+m3Rp1+S69oeQ3E+pLwkH4LjDEgE9IPz0NRhVsQJlV5zftWnNo7p1u51+EOGwKjTpaEUI
ze3m0zrIYQAWs019zXVb8IXtsiLIzxtbiqYWq/bT7TWToJGJgoU1z1j6vDPKgvGDHhY9M31j7lxA
Hn7sFtDsTDbaB4BuqWjLtfiJAAexvxfQclflkvgv25mmj9N14Dx3PUNZvvuFl6Bbl7vWRaebLrvy
pWrDA67orakKvKvk01lSg/5YpMqz2V1QTQFzk1KYY0lsIgsOey3wNVGsIIjCddHaRR11w2XTXAme
4jnW0C8QWbCHYqOJV8z1jx48tiP+AQa1QuaY8K8ftGok5iRlg3Ce4Z8L6th/9tPsKCf2Sk4LxmBY
JI/RQsvRHincLJFAm536tkNNpbVwt5/y7HZ0pDW0EMF9ompDpAkuxC1E8k2WGRMxtsYQvb2URBWB
y5l4KHfZPyLRdd1Jp6w2fvLw1R7bK95r0SvjO1B4kTO7PHV3ZAAeR9vhDJzL13VZHYamQ6T9Fy2o
k6F44FvFgSVLbICIyyQ1RJf5xPimVuA3SIugNLPy2vBYZmgCG+Udc3L2IwttZTm6sFUg7swkN2eq
Wa0OxbEGMrHBgDSl/Pnu78hdLAWsaKNrzRQvxjTAkYlTOVBhK68VS7nm+o1+FoN5oWlKF7JTr0Tk
roO/45OSQMToEkpWpBAMWpu4UOFE0rbLnhKTPs0FZPtVF9uKPsnVgybzAQhMTwvf9PFZ9wOUpSMq
IWiwKXse/VLDhZn4B6IoFBgn/EQYytEVU/N5lsIyhMivBLay8sMk/py0PqEbQbj1jmyKgWW2Xi4w
AZW6+t9SKzP9/2e8QF4gmMpOCap0uK6XQqrSPs3cDg7YM5igmfOjKHiO/omV8U46J38/P3I1ubJk
E0rNm5jJTQYb1TENodUNdajElaBjORajwbF5EQAsU5+u0Iy3PDt3DzCuaqJMbSja3Npm74SNr6eV
VfZg9VGUBxeBoZ58GKlV6Ln2hLNc458YyW1ectr7w/v6XrFNTJdjWqvkyCdUAvzDnf4oX/As7mog
gwdPdjyJ28TFK/O0l9eZ8tdIfNp6YGkhV3dXAUFV9in0vKE8epNXTLTyGCcriCxiOLea8kcqe6jB
DNJ3tf5H3UXRsU7CoqcF1LDfUXIri/glqXSAE7RfoIfI34aaESvqpy1EzwZ3WVgGwvBtrXKJ8crn
ezUzocmm/ies2yGWLIBiBP1aQLdT1No88tK+LVgh4mneTi1ihyNS5DqSmsvMUK6Z2myqOGv1cp7j
lf3gOfotmCnIALj2YlhWD+QEL8eLnOvVPlrVD6DY4LoJhKLGai1cuTj7JIQ57AeqOZSRFh8DzQwf
1Okyt+PXPXxhj8IYPXKX9hYqPzpDJzRHK9TuoNUiRhh7EU5YghC4gdaB+AE3hMPxrXCrB1I+KyyR
P9GMAgcZQ6AErFLaDRfQVfknwWrwVsmdfj2X6VNvlYT4ZL1HYkgx96WmLaB1nniQzyIK8vPotP7g
ONanG2XbET3oXuWmiijvQZB4bmN/jgPkvGfepUMs08q99DgjRWjMIYTD6zDKsFgcfdwAewH427BF
VaQl5YXJFssDSX2c17kR5oZlGaiaWxRhebW7YUQOOY5gvYNhk/ty0zTJXzkPQfOSuDxRuiCLeeuO
v1zHq+6qeUXcsV9ATY5lUwQNf9nSixvPYqAVukmHLuTgxIwF3rx4vvq3WZ3Jqn1b7dPeoqpd4LdT
8km/XNXWcfL/FOFhjWjnUim3zcdXgag1VtzgREOrWIQ47Dp7m+span7bRIdT4s+bYMQXdd3QIhGR
b9w+nQhLHdy+80VgJZ2EJlyc0qpzNLgTC2tW7pPLtLp76akKiH70Di4QP5z2OWIXUhhQYt2a6b2v
dtE/MSV5m89IJ1JJ8HsZu6UfQWLryhYTDEu0KCP2nMecEjtmRb8tfHpcmA83W27uHzta5hfT5oxl
v09I1tO0kOSveFJdJj3s+Vz+m+H1KcWMl++0xxkpD6grkPgSa4ABqcqIgmG3bcs2DRIPVrM/z0Oc
tuK6p9JdnFC2HKI8WmZhLwcDUGQAlnenvD33KBZtihyX+f3jzuWKCP5mBgOlpT5we/EmEbHuXymT
QbbxlpgDqOXITi8rP3E/Tf/fdeSiswUfOBlmee8DLVCtThXEN7yBJg059ijavg9sgj5PJuEE4LeY
LAOBRsvpLGuRp5U582+U16Sy2nOznVZp/jKyjjezUpufD44BxEjS8ZmsoS20NxQjW2HfIX9PKT13
ijLPlINZ2GqRZWa2AvdwOu+dJovTTYizhOArop5p61OdX+ZBE2KdcF74UTThBcBaJy0aH+eIRRra
OXdablfyLzf2ddqdzZuviorJDfVZ5Lz7B8pVtg9XwakwUGukK5buiNFpUmi9q2mF4XlfMfGbbG/w
P88UhXIaTL4a2HJpIP1VDxXTDOKTBeu/Y0zpGSvW8ifQYpFgIKpZZk1CfsUWEzV7EVaFbXNU0phr
fNMBL5P0Co1uqtP0cJWd9jyTfyRyGB5Hxw/z8WEgdzY+UhMoalJy+tww+c7eTgOTZAF2LJj5+4N5
fsnJ+tzHGo0gcmd9wzxVJKlN4x+WRugHb3YzkwWE1ezRTlO7tRqD6FDPfAA6KdSvvSTKtm605lR8
bCbPDxVtQxkSUVS1FSN4XuVauX/kGhinu3zN3u5vyg1ajasjj1uw7ia6a+nDy8irJ6daqucWQyw+
Tf+5qIDMvnEcHOCQYF7VfQqIzaza/4uj/jAWVjPFZovEsFlYmM9JkgcF1bqa0hsQoZEpp6fK+VJm
9B6fw1tjkpBfZ0Qmr2P2FGaz85zy1JwQaQm8cGs3uWvTaeeVP2KaDa91HWn+msNl3T3UiEyXh+0m
aFFAVrGIJG9Ci/3YdxBjNO5OO66Cl4xIl48OQn9kyQNouKvjCRLj4i24K+jwyqSt8cE4TqA+VTqq
VNd6/Sg5ze6hPP6Szy+hQBUXUs95Fgp4gOlTpFl/fEhBLrJdCu47WeGDyJGR0BqH4ve9BJiGngKd
ACR5E6RKfPJDJ1RkTrPO/MLyIu5Xs0+2fyQWEb5vvARLLcQedG6NawtJ+yrkxa9h1bJwJFZQB+bP
AoHiQgGjSx5349sJjqqhxc6a7+5p+BROqXVcBfsK4FGHR9Dac5/E4RbTNnvyogbVBzgT0gO96hJS
o8WRlIwAf9GQpQROwNTmacPUIOfsTbWnPgtRNS9jJN+bBt9wLANL4DAp5mSPqxKJt+Z8aPHb2b/p
HF3TRxR3guiUvidi8oG+SM4xuqUB+g2dLuTeKB78nhQzwacFmM5px6+zHFvcrHY6MiO+p+KhdpQX
OSNRbuIyubSinqE2J8nYPCnoExSsatzWW7IkKn6xDSxUfizst6c01qcbcgffIUujrm5d3B3aiZMt
vPJyGeOthshYwtkMGsdw/ONdKEWIVZVgGHez3fUoHdJvRyuzGr927jXnLBCbKjn2B7mJ0URilD0e
g9/LSwTJQJkTqHXrI4aJy+m+BqO1aDjQkNXujna2g2J0WBaAuPyRgpUudAl0E9YXQjiaEuuGjKkL
nyBb/F+sXpHR8h6YalLe9weFJcmxNkfdnqmu/IcbPcBUk7laRVFGiXkJCwRugXOK0YMwjrbePIu+
dV6g1oKL519iAcpTk/gXid06w0+jOq8tXrIZo7RYpvDu3rSOQaXuTRKzxi6Dybd39nnf0P72q/a+
WmTcBQ20z0Dm9b7Us0rrsDLpFdUwsYaNnR6jGaJExfLYxOhZcp5dDiDbCZidQxGeoY77ItWwaKVh
8PXw7OcSM3XEMSnXfib6V1QwDZaU+8RqT7kU22z5zCWVbugrctDh/0OQty0SGAiPibRiPjUtbd1z
e+A5PETM8u4JdHSQUPhCG6rGrVIhewZD6SjGjshcAlCISVjWuJPIc0/miboF2w1tg+dXQOEfL0dr
Tcc614qWqrPXpWAEAG8/u1EB0VmQdStgFZ7CdkPZXSBSEfuOBe3dOlYRd33IUDZNRwFAgsTiBQXE
thZl8mldO1lx5VUQVJ3Kcu09XlzTdmfc4WKheSDlAH4LGDOaQfeeXkQcI1aeb7PfxgdAHnJgGwN3
k4DI3z6IRGAxXoJMrtvMdQ3o36NRB8IekyHxzfcMNjZS+E2zwq5YJ1xR/NUL01SD/1YbCARv9Pd2
dDcfX/Mkwh5m4FMDcuI8ucX6YpyZNqwKY6nq9IkUymJuBqq3V0ulbShex4P1n2sLBflDL8mO3u7l
+SLP8ips8BxAq2w0NPIvsjAaGHBe5uBKIjAJ55f7w5nJf4Ni/pA9zW/G0j+3ym6flOEGvPkLKSGD
sZX4recsHoVJdp8UP6pRToB/LgCgGBtlK9ada6PDPP+FZyarz0l81MGMI6dt0Q6g83QYpkkoEDmh
U3XlcQNtKOuVTGIJaxGTbGHZ9pH+Qkolk9SjJWwjGjrwQN5NtVd8T6oKXXHHmHYeVs1Fd1GT/e0T
QiVEIU6Jwg5gmgSK3pa2nI0FLeWq2vMlhX8PdQ7Nz+5tyT58e5OQaTPu3RBe439p3qeETmktkiIN
6VtFXjld2igcoVYMUELPzEE5q96Boa1Xa2GZjpakfpJpRMdlo0V5kYYZ935ZMBruaPYhxBp0EK4F
8ShfE3TmiaZQF3hwDC7Uwn83tv/Y7xjHOszTB5/rYt9cgJIrkWGyKeJ4T7EmNaaw/tvU5eBiyEXr
j3+4i5vBUqptA1Wz0dRGn8SVyTzAnkjAMfzSG6vSBrraMOJawYZkcYiHKudEbmGzkfS99ga9kefo
MHa5nPvBfeLpVDaf8+HVDq2cG7ehpLtgZ7RWcL4e0SbFDYrF+waEHJyeMXl+jZ3MOGM1FeZPbBEh
KwHRCC4jdvWeW4IJsI0riMno8nwOrlcTBqcEZ0OLqhdr6tb5KQF8sRXiFwa4MwtsYy9j4EkrNYxO
Y/N5uXyG0msXCNkwr/gn6k55F4K72b8sk0g2Tn0CWPse3Lz/485tqkYkk4OPOj7SlB0t1Zezv054
f96/upm2BhTk/oUBBP2sQ9dlfexeuvpXMUoGp+7Am/7rw51L651vqui6vE/LZYsKMbfY66kYGfUQ
Jf7ovfrAqcBFGetw8TlgWsjCnfBmyOIgmXFQIynQEi8hdp0STphYu6ZM1CYyGzZ7uUbGdrVgDg8l
qhOX79IISDIOYPHYZQI9XGbsF7K6P7EQdH9gBR/tU0JzqPhRJRNp3guBEf4xVkv/BLRcDgwM9s2X
kEsRx89DzmEyoLn+3Q3hKyPgvfS1rrjrYLjXGduzvHvb4GTlKzSLrQg49h4sLIXFTgIezTy9SRdh
Io1+KRC8wXHLZ6Eq0qIYud0kn2eQv0MV/22BFSftaWdvfSa7KFuBHxhc2AXqdRITXYugVPBNgv5R
eBsnI4WvvJvu1Sie+H6EkaIKC9TyQEw9mq4RFesUlGykitUN9qZVhVGXkIqLtJdxeBrPeAZ+rkMw
4mMT+/iGJBJbHjqmRLX79jA+ju9ZQusHJwkREbhxMilVlbiH8Xd9sSrgMazym/e7jLStejtUHDXw
6NJFG1D89DCoWgElh2rpsCAL3zArQVgB/voAxG1BxsrLaqdzuBT6RXAnX8EK1gttKTUjHWxFDxAZ
3JEikbSSK0XZD2lMYYensM4NccgzFIxutiaaE8YwUa8jW6yTpXRAqzY8vfgh7Mp39oR8BQCtKUrB
hNOKZ+QWQdP5W4fnJpM2q4c/CnUtv0wH/RU6BnywXdougl13WiQsG+XCSwTcJg19x7O0+oFfC3I7
115mfFujsWp+6BblG88EVLsgEXXYVR7O5R0Wwco55Lun0WF+qgbftsVhNcu3qUXgFE9bnEbPvEaa
wCeMcfe7jhEPCGw7p0Bs59qfm+CkX7gTVZ8ezW7lABjybaiuyb8Hymp40ak6G8FvlCnQ0LCMOhVB
/C4LxYNoxKx2CqoDa66JZWWzjRQ/um6CfXlSKXJczfvl1ARIgeS45kNcjT/Y7lo6/57gUDrq1VDW
29jZNepWyx2SrzKsCLx7kMpsWIFWQWe6Tt059lSz3OMnSFsJbNYIpehUmqURFJyMxhMdZwcKmGsy
ISwkuHZB79JKjKLn1+ikEMi0Kel1/OuJ/iJgqB54daGTSW+QXj6vhP+6eeI2bHLzVaUW11m7rDiV
nJNpeOqwcvkCJute6DQZWYI+hoSUc5nDdJWNOVpay6WlcbRiivAFleyN0JNy8ZJmxhv3nGsPHVWA
7Om+AK9v79Uu1UtoUzF3Jjp6eI0iMOc5GeW0A29lJBwGyrHh334YfQ7/9U9kEFh89xD9wO2VgqjP
/qMGdH0Mk/DYGj8QXY3aYRqMrdIIK/Ud4oXgIFLXlJsg+hk0T+l1Clj9aJfqdIDwmL3+rr4oEHOj
blaghiFJkJqW9k5Dl9iUocs2NO096MB/8MwS/uNhxEbVflqNEQKXzXCDZLdNulk4LvOQwy8bsTOj
8k+zaso8ZZPVecPhiTNt/g7CpTvoUXSu2VREMiw87M0X05iRINSQJdi6g9ytMqVgPgAFU8y6nNZf
FLH54VwRK1pgGidUOzVRnrBQTlKA97moORZBB1PwNRY0Oi5dPSwmNjBi9WKQSgoSa1KH+x4J0CHZ
/3u/YxWLIaX6t28yXeq/yxPAvp1ub1JU1HKNkyuj4bbVURYmPqVzDWncSUfqrM624osjAfRu7BQ7
MTloXlgH4q7KTEjupoubSzFL2D7wbqjIOXOXmW8BizSAX6uP/TeEQmkan8ft5Mvn152cbxczHtoA
RNQEG00gKMgvJSzGK8EItHjauzJOROXC9NZylntYJqLyI01plg89EtHH18BiatlMX1jzAje+rbK7
vjA5ETunbUsIVGf4/0pdKr5WJFyeZEVRG8skCs0HTlwYtssuEVD4fNTRY98BVvVsOl3ioD9E/MIc
F13maLYVFLMDRuh2joWWUAg3djk2DlDiu05G8i/fVLNg5+8q9VqeuL4WUpZprnNKQwL5spj0I2dY
nPWDFJ0tMuenUNPjFkBQfpE93Vyx59CmdIZTqbSHNbR50E4FhIr0eC2QbLP+ErCClNfdbyEvbnF4
20kVEEiLiYKfoq9R+GcXouQoNopx5BMqyjYke5vc6gprb2Umvp21AzT35Vcgsib0Ji7d6PIVif9X
CIp9c3jiUo6TbUga4qHIVnGu8rZHj0ViaoeqtvTXkOutrgwf085PrqeNIRh6o0cHzKsUmCgOriEq
h4AUV/PibyOmGDcTGbfV3rpAYDoQtMb9q+ftQwLSpaEzg7CMHMqzP51s92nibz/JPvTJnjUdmY13
XbGNrELXeYleLYX4++MAQYFnhK7vdCaW/8u/RBNyW41H+zGbDHdNrEUFq0CAG15bYxBdILWtaXvE
Ez0YxFl3L+dtFBv173r7y6UcF7jLLkEpZzL9vqpAYSYIcxPGWiZAa2QUUyo6KZSnPL6BRp8dht2Q
lUcwPLyeS4guXH3UgaUBcIBa6/t9KgGd/WYKNZagxOkwoCBWTrm1BI6+JtVRdVKIMrHoV8ZyVbtK
HvEeM2OASmenAke+AnGjMawhfdqrubYQMG12o6dUaIdhUAgZvU5B5V8Q1itg7LRszha0o94waxHc
Cmx19KJInM/quLNgITFMm+twWWhA+RZGEMggDjWsDXGYXbBEFYGRm2T2ngIfHib+vG/NLsB+dinv
HRYjUh4yXoZRn9TEq3jFGh2Rz71oczYcseXWpL/PsicwTQ2u73MoNynxg11p3n2ZMflqeGZK68xT
ieSSAX5vbIIh4J1wr+ptXoWx+CyiK+uSEdQk/YX/S0dY0V4y1nX2tHbZ1MSP+6XzHvSZI8BWhOR2
LUK3CGCOgG1OYVQgXUO7iqesOBEXQujYg9l7PN+DqPJRiyFluRLgyJPRgXEEeWmfhatWF6EgMejx
iLwq7TofIUsqIhjq8dp2DTC3q3TaIwph+mYTwlUV4VYPhk/W6DanYrqf4Xw2KR4rtJ+4a3dBCeXC
Y7PJa6AblTkSPQ+P1uwGvsP0E3xeJ0CVi0AKRcDPDfaJnprqV2JUWBU3MttGOpBsS0nXweAvX+L0
LVZgRcPCfs5Pp1/KTCDPcsWmITGlnhyeBgyNtwIwQCtRjxcTyY9RPqqT3CuImwMFvtgAjQ73ZrlF
4pvptlJbNmJ0SINhP0cqHt/JWBU2nRT9TYNoU+AVsLhWNijZjHpV4USg3gsKvuhyaT5rmoH36sX1
UKZjAtq8f8UpJEXYaVPOHfkjTSXmQCGcEWeX/i94/6sOhvwEZgzgpmBhKw75L2RCwFlpSan9d5p8
ThZVtZB3bW47GdZLDaf8gly+AwkMnUMGcth4my0pFA4BaIbDkyXm0Km4iqTD3ajdZbGMO1RDtfev
uzjWUTKd6ZTXf9Mgp8lPh3rPpY9kqmkDV42YNtlz0QvlS1d8Z4XPThwKnXTFQCtiSiHsSm3Eokxh
KagwJwOZzB3vklxtcx28CoDiH+yvsZb4KkYpP/uAFBkdpQrhE/1w0xtDJt7Eb2A/MMOtfZaS+5gL
NSNy3FpceZFXF1oZBklLf93C8PZpwjp+QDftaU3C+nPk15tmX2KAx8PvwcF7U6oF0aWsv7a9jqTg
qF3ldGAlMiwH7Cr86lTg2/+nrSJW0KyXWELA3a2OzWaUhRz/xW3GLAqtBlO0CQEj7ZYyVeVXZIas
hAFbmQVeMHMLqUu+nwDWQ+VJy/wyuuPrInsDm+8RZISqvf6EaDQm2ZUnVk7BlUKzdEGqOpW92LNI
3opGoc1HBiGsWHi+QSV77cjxP5dWVrcNWnl9O0cYHKlX1S/M65aA0fQOLbWsJud7aAbUsmqS6Lyf
v7sexMewUxB8V9qpwHeHCEm0k3L3K+lKQvdmtCAKgqQgAQ4bj1hY88MvnRzM1nzxP88ou84yARu/
ZJG1RmsXQQ8qhy6FLm2ghkoAT+7kaCiaUbsfeu3d3sZPomUMEoS2fasX1YMpX1dk8OAqRhj37E2n
HRNV23CWQpLWOmKCYDn65f8Kk68HLBYlToBzj+gKEWz8jLA9uuwPAffTazjnSjuwNE7r15z3c3k9
xIdZfflAzZNNBAdnwOZW2adJH1wLKULUgGoULjzCVMqXIPf0Cb5Zbq8MSdUnNpR8KMcDYSzbcn4b
9B/IfFUMAg8jgNSwc1qotPlWzlEQZpZisQcTVkm3RiQkAb9qBG3P99ekAevtkDMzVFeHhPHGjl5X
I6YnMHz+ePFiG/q+ZZUv2CCcEv7Qq5+jGC7lqv/3xfvJYY8qXOsDlUeheQzztQ4PoO0/WrFiPXn3
eLkaTBX2we/fMOtjWpRnKsx6D93/ps08ZMZrkbpQhVaF3CGguFet5GU72LRph649Xti0dyRdLbFr
mCBDCZv3Fe8tyxvc61f5pmQPyFrlFCI744SL+Kp6S8J+RRVTopEGufGtgTg3TqiPSGu/ol6JKCzK
689CvO1he0cblL60sDzkeF8wlJw0MHd62XVpTzb9n+MoFaITdvs4wyxqnu97K1Oh1hzGwNcvaBcB
Qv+FZxFy8G0Slo7RXgZxBGixwW9Ir6CUbabRet8hVVkJFV80KPEO77IbXr8p8fKoZxc9mQUgs7aO
LUM/f25jdWoRcncbZ0rkAbgF1ftc0W6lR19vLpl1htGvG6hJMyrwgTQ+JD92jIGeD77d3Q5HSRvX
YXtlKDzDaVWnVIhPkqI2Jgl1db64O8m2aF+331LsNoNrFsnPCyOWn+qJrCJby+B/mgE5pwqK1lbZ
+7vX40+4Ui33ff3hwi0IkxjpBpoSLw0Vodjk67XINGhV6j2WyJUoy2oxeW6TKw59MkLnqT90HS3Q
TkORE89j3ltTotU2BKTDvmKPPBtoF5ZeWBB1eAMihg8PpS95VN9stSjHj/CM+gvkm6w4KJ9UE37o
zXliMckf5YRQJggBh16l+JrP/NgYkcsmZ7q8mJEyOsxqwV7idLdvSn1NYwOlQpNPyIax+0qYF/L4
uSjUoK2zJZDpaVLt8HVqKjuOwec/srI80f6QiNhylpLnID8s04kS70j/v+FzvpVWKr5haIyUYvJO
wNzTufYEiujL4CQpXwt3p1dGiIjmIOZEFwCOyGtNL8lBqc7gF0FpxtgLyZ4WXw56nLg7VCbqx+9r
bwsZ557BUUk9x2vUVCViQLjNgdU2oHB5q8Ydc+QoP4l3CnWfVkUpo8dvealgija8fq96RZ4kIxiO
J6V7LUuZy4pFdaK3kyifYZXAA3ChQXolpmn7y9lXlZ4GmUm6SwFfq9/sGwNMBPIZQWBGSliXPDiB
wgRi83XmLTPRA5hiQP4P/PrSdviD5Dqtjm2nBFafSpWQonLAzOKKvrChMMzOSxZikIySEEKUP3jz
+aJKchV4GRZi2OJazkMB5x3hcymM3yDAAO83Y7beEKTGH391BfL+QN2yB1GKxJK5GEkgcp0SPnE9
/bp5EUqUiqcvmJJ9wrPQ2MegqFIzzJIqtWWNnJDQzb414b8N7Vn4CVx3o/3yBfuNdsRasGVnTdxv
MdgZMvLjj7AOPwxoyzas0xYPjKquaEGNj1LtXoTS3BP3/ouHDGTDC5bkPAbphwLYe3ZNKwpX+FSl
Y6SgBT10ceV16WFIvUu9kv80EMW5PCb0ya1U49SIocfaO1Jhy8FnPt0VH48GhoZ6B17hwoZn1q7u
k5b2WUJ714MLFEIyfSuWAnIA+vtUMazBA0iAxSDz8d3+VogFLcyzvFZJLlzUQQ58nG0bTq3GU6yu
vqAq2ScGD+4enkGDlhZXdSGfprODM7ELajkD2OadLvBoXFy+YiH/kSzZnqpaNRa4UVCjFQZ6thnM
cGdQbY0av6txBkHGHsw+peAl402UtNqJvKnUXlT2g7/K2+79R8T2JhWP0c0Q7KWSfYOyIF655REf
Fv/gYQxM0T82wt6RgQdQQKyU+2Ryvil2o17S/FooLAnoN/NW6P7oro9ypAIz/feUcZdPLuOcG66q
CyCi9b3RVHJB9X5GdTMBEEloZxtHyPnOPOCQoYSf/gqLo/eCQ+WF+imB/39nik97NUNOH40f93TH
9cTl2o/EpMsCte3wvSqtNuj7rR5RnCPAxDnqwu+X/tcl5poR7/PSQU+/1wMpmWFqaN7zDc6NdNeE
j3v0ElN2Xj9GIIwOCgUZJeBfC/JDnJGf4mTjzGRFhT5QqicJ0Khch0g3H3AupJzQ/z1F6iMijfwP
5F7iMH8ofHWu3SB6S+LfQ6XanRR3yBbmgCuyvp+YsxQI6X3clFLm7vv94e99fIrJgm1twxHcuVYK
GqxFUs2J2gKEhKnKRP+hJzk5vx3MlPRhZIUTOsoLUmIp7RFw289e8uf0Vkd0wn9xixZ5VbUstMJL
8GNx1pY4JsA12hfSMJhz5UHP08+p8YfUSEOGKjnNio6gdb7k2NkjBnEabMk0JQ+CO8Y2UFW257cv
k9GOL7DisGHgblAlwfMFBctSx3Gxme7r0oZPlywMh5Z4Y1Dw1HK0wYvqGy4tvPJ1kaEKPmnUO25M
mSeznscdtQSaTceP80pTvP085rhX8I1P2OdrSj+KzsRoPSM9HazHpoVQ+qoons3oz4zzuEUd1dQ/
62syMRw/TTd5O16fN9cleAXFihz7Gs+U/m2j2gZFZl86u2JYcot5wHNSTezzj6PtJ+f3O5DNVJat
5jZi2KF2qhiXsO7t4qH6euEOzRrRX4EH5KvV2fHtEgce+Fs3fulTOk8u55edCptd5oMWezBvgS1b
8saeZ1Sznxz4Fz0yFR53OE5mh4NuYzu609vFYfs/i5go2sTWTYXLpVG6XGCONd9xVlsJHqA5GvXz
vMvzZJWXO2byKT3CXhXqFe9wU9uKxU9SoRyJJb73nZ0u5AG1/oBt/DssuG45YiYtRs+vqa39ir2+
YzqRImNwFSJZfeIwC0bqPahGJB2sUSQLovhZZrTW9Z0YNg0oZH7gjfyxh54TRcpZAafQNZf6B9cT
BDd6cpaO+gIlku/G25RqcjiHal6+jNiqI+aLqr9NmM61Q6HF3rIF5h1vYt2Xifq7luDTlt2YvM5Y
Unox/iqzhVI/5mB8Qim3FaDXCs/ZEXdkoJSHEs2shya2EPH1spzINDq7XAQBox11Ihs3doBTwTJG
D8Y8alata6QCggnnlpTfwxbTpjiaqEANy6XdlD6PdTJBMZ3yq7V33zkg3ncitwW1pWQG503znV3F
Q41KUrJPXmepZvWF5F8BA3mD0XHpiBF3oDYs/rLr0ZbhVMG5Im1+un/s34EhF++9BdpZQW9OkSUD
TDlq47/lYL/gLq3zzehogB2m1QLxyZroOKW+xGubBjQmwLhYovRkMtTiqFN2fHuoC2ma6I7ZAbEl
9/nTdCWNb9j1wqpXIq3rDZG8D3k5C5qSLqGaoPSa+u4GWXmU6PkVn1TG4AMJP/gTI/PI5xbCzfgF
KzNyBtEBclFdHmpZiXWEKLt3lNnASi1IEVmzp7h9hb1aSGLTyrw2Vj3H9KcoqX+HfAxYxd7H2FaX
cQUMjsjftxkIV6OzHf7iXo77gT88aCXYG4Uix76l2HrfiCWRqIiNon+QbATY37J21lxAv031DsSB
pzDgg+e4iwjvSDb/GcYE6IUNeC4DHAMISDbhpBOuIVyhNxss3fNLjT4eQMA7NOyPqMOZNhJKmyLi
d3yaj9Ia9tj9s5T3tjr8ov7uLGyKkQeTtqpEN0j10YOjOvznN6ng4OWz4UrP2lH4Ta+RWFvYTRdh
P2F5kEiAYjp/lkjC32F5klZKo+aXJmA5kb3/jvGtksW0Tb77oGKG+U5izahFlnb1tyxVnRUODcYe
ZNs1wfbvNWmlmY9WX6Z6qCyQQ/ZxbRBT/JTFon5dT0tX79ST/8IBmxgNf6CXgO9MK+LnOyjS7+O6
IQ/AjgCO5D+l01Jwhv2Uh1VoDlSi/z4aYuu7/rrVsvLfjFKgGnhukYODhpS6eaMlbnyKC5h/6DbN
lHv27TCTiFAQvelLUimfmYswNc49ubWtoCPm+56PVoOg0RC+dJy4JO5j+sZf6jlWOvCemHM8DMLA
LAMDPtVIRKri6evvFAqPF7j2Le1meyIVMSUNVr47N9ZB6c3HY6jsrC3736eDJg+Uz1iEvgwwvLzA
rgqsqvtHPdufz9uIVKJ771SFvOZOICNKAe4+kJSwS/fGHdLzJPAQpXLdDWhIPw+/ue0gjAEwDy09
pbscMKZwUWkBhhLRy3Jdf2fNSJmdXYYOW1ZVrlSM9J3+YPPK263KKjOVaaz22Uhn6USj0IwbqHfE
eYA0qqvoQkf+rwc0NHkuzufMhLUY9b91FL5b61tUEbcEEFHhVtx/7PwY0PqEdTy2L5lNInsolqGE
jbHjiTIIPJ1cxlOedlhy2P4ETvqH2bdI7qss2ZUOWrkCBxgkJnSNMbUFK3tecCtCiVrnZlZisa3j
Lr01//q5T2ARh8PPozwJneA9gmtFaGehbxOMdEOWG7jmJwz5BGV3gLJWXv1XIe7uzVwC8Bbsm1vT
7C4A2FQIh6KdiFdpUVOOouQSchO3S6piOVVIDP4VXXb/wqV1wVvJnZ7apk5AleTwisoATONmxw4W
3vwQBM/5KGX9PrN3Z+p5XHvXou7nwO134tEWvCypg2eowujzigpX6oTVKliDrtkM8aSJWRaVSIQL
nbI8g6TH/gQSSm1HkNiJceUCje2/KO9G8bkM2lVDY6+A2+FrQYaWzL6didqEZ+QLzo2V2gipZ19m
5L02jTTx3wEIh+zbfKaLkTQJk9K03vVANV3ZPC2+q4VUcR18ONgyKVWdu24kArzHM1BhTEpu8QNR
Xzy7MnVwA4Ymp+JxWfmui66nwi/9tZ5yK7MSOLJMGI6yVg94XDPD0MBe678nLmAUXGyhsoj73bxl
xFJECf/VkxGO+IhWlHMulX1A6SmfJuBmTBbVfL3amN0dJFO6AIq0yLSOFINbH0Zcd/uXqeItxmUh
L2/xHPfmhnzMX1BfYTJE5JHizji88k3obH/7EYvMP/d+25HvDuRPFe6F7ZGWAHD7ZCgCByvnuZkV
y0stTfqvE5RfzqrQ6iCinb+FrYVLDlV+VBmA40ttNl+WQshRpyUaJRZKP80Up5yAmpTDSy3VAVnu
tNjXfZjHPGOgwcuCWKLDiP3qY2kvR5Kcw9ISMQUQvvIrY59sfNY5IqeikK00+yzCf22xiQI2/Yhx
Q80S918nrFX9PbMZizcflwxfRgW4esZ/j0blfDMt0hkmYYyqYx9WrnWiYRLijK0CG3gTi9irdOb+
XFNH9jkYRnqCPvJBStUeKIfLfSxNwR6HaTBzldbiEK1OdFOChz4g0UtGWv8sGvDLHdx4AZwO79IE
hOPQsHJkM3Nd+CfmZmz3wPOLOLIy27aZMiCVuwzmr7TUJt83wAJQPNslhnqhc3hqz+WZD5dCcN5q
Ka5niVXo/CuEiy9cqLyqXEI5fK/xJqUhciEOlR0qwzJnWbydii9Y2TtyEnwJhliHe409a9gsSjE5
qf6SWzHVbSdVr0kDSnp7nhsgm2ytIbzhKc9EsP3tsGhzfez6P7BRaxTOTSguiN70kebi7rFXUQ5U
UEkSBX7XuFcx9pPIa4UjRSKJrdBLRcv5V/ZJ7xS3dCcpOdyC98JHp2okMjUkz9CeGYou1gtNn1w3
JzH11RVNBt8qLhhaaNyJhPApxMUl/HKpuf6VHy+vIWiHlHQA+KbAWxU1jT7UPGdAH04WGp//6uVF
yhVl+lI3cMc0gJlGhfHThUkMrHqBzSiBbRkGjDdx2yACzSmhXqjdgj1GzZrhbx5gGbk9DMTG0APY
5TQLvLMbt8wxX6wW0x4XwASypALMOf67UuxTQjxMc7nMYWvX2H1DgmhC+SG/EC7RcY/x/yM6AInL
o+TB9stVTfPsV0wbtqdzDdiEMhtfqoTYiL3EAO7PLixHNEY/Svfyyu2scb0rVK1wVbFtJgWHSLiW
JP+nVYi3jpJJQw8c8MT06cf3hYV/DL/fRtlWyiDp5ns0D6Qc14JMRXAMeVsXBfvb1caHe6uCl2Qa
5la4EA22hh1939ETa+ul89bREK6fNP3lk3wf1dyXS45WqzZGK/K2RjFVQirdRSBZpa87IOmFm3B0
N7M25V9iAGXp5VrzX0WctA2TpwqcPGUDOwfU6t8IT71giujzvYhhqW8TOjV91KEJ5ZkI5YHYkfxo
mS3UrE1Wn2b/aEGw6IDrlQuHfYWea2XEMTWdzbNG2kTwiDHyrt7RGlzqkftufwup31jGn1QtaSTL
d+EJvpLcLzWrREK23jsL/CPJuDqmXpzhdAb232rZijRCBy9Mum5lJgjVuidyE4ZzHoAy+hB7ueRn
R8tukKJSSYlLNE+4lQsT2RtMfc9LrnJah8GomFwsI/46kxalqMVd106QtFqUHZR+7m6ZWFle7aD5
WQBLOI6j6VDn4g1Y1rGFhj3UNIMl2Zq0LusM/0LIR1JLNTH9sPBZtnbC2bXvwNJrKvZrjmbbNhhR
bHJBVD+EQMDOLL5dO90VLTpqlxlcMd/ixqyPjHASroegXQFpj33w87pSPhJFMGcDQVJiUbFu50f8
5A7sno73hXMRxvZ1vBdjC/jUj8MxrjPu6KwgwzQcdTq28TFXio0VH7mB/54jMSGC4UTERmmKMTMZ
KnLfEan8RFZ966Jv55cfYdz+R/bAg1Ik77ZE2Y6Xc7oAdD0wzM2CU7yjWPjF6yVmpLGXaLiFCMa3
5Kd14s62KezlBWVPZhS6UaygVi//zeISL4jNYe4ZUdMKHTMMxhRbrs1q9lhUd4HZme9FtivGGLCJ
F3b0nFBtWLxMXSSxL3b6uGDNqbqe0pqz5o+epArx/shpPeFarnyjk8UNhCGT/E/x6nN/wrNN6rMW
/GH5q/GhMK93EuoT0XzLu97HOdI0yX0AByLDxsudEeVuYwoxn+4xR5AMdBjATU6RJ5wXMDSHUG3V
WgbDpskF9XJnqqKlMjkp58nfLynlLQRJwe26JFikeTb2/ta1yEs0Zl830MkhS5k7x00uTcOl3T8T
EC1H1haH7bX+LHSYB6MjpifPEA/6t4xogHL+xhFAhwFM9TMaCyqPahdkUqP2x5AEeXlWTxvRiird
CQv5SpL/J5Xy/tznx+VF1PW5cuMrWgjJwDvOkeC2dJXnbpkrDmUWRB/8K0hI9gt4xeqcFgzr8uOr
km5Ro4WovZCwxrZ5qJyZjNBCAL08tZjKgBAeivN33qaIr/rMl2AdB4R92deejD/5rLZRcmo6BWyg
eEBM9tURjvLVlSKH5h8ZkNF8q5VGHlAyft76XOkg5IGVzj5eJTGVuegJ08EQkA5o4RhVvlKcMR1x
K9mdHHIfCcye8N9eWObccah57k4nUwLU9de/grjVdO+n5W5c5N1aHGO6YMAuSVSSXf5c6CSUQDT9
lnz11z3lUKX10jm6SY5nXEP/QCf+OinJWc/f8V4yZJnqXgIDsRnxiEkoKA70gFJTcm5suX3NfBRE
8Nq7vFn9JWxV5DizmdEEtDePkLZAt47kN/GGRKJGG5Gq2eJfTS3WJOxY5GG0Y/BkMVS86Tl0h3fL
0YoxTMSmUwjsW9LsXChV54vqivCCqLdocNTki6puaLnloQGoHmyyXw0ay6GKobzlPox1FoZ3S2+h
6cUo5dsXpbd39oQvzrC0Y/T2cX5t2uIsMVhuCNiPfmGIxSe/kVupRw8+/Pz+vPOXhQ257CNtrv9I
hMN9un6zfV82ErSzn5DlKMv+kZUtFjdaobbLNa2B75bAPsuOxzcaBL81RItsNNJ5Q6vFkC8nOH0r
joud23tyuxEL2YssHedQ/q2UzXPSpIFp8cykzh9a47Rc0C5ZJ+5xA64DJfJKghn0P2AoN3/Vp2E7
gC3e6T22X0NXS/+eZEhFUVhI7+i0WxBOTssXGuD8jidxHzJOhpp4koIu3TLuiCJ7nnLwweWULZHR
+Q1HELWOrADDjvG01KlO2YPPmM7vkU1GV33fKeex6I+ZZNiKTkqDDRgvCavpXEU090OgOwPtj+kz
Sih6BO0/wSLeKV4e8fP3m450Ean3tRsGqQ+f5dTRhUd/nqbIvtPu5eAy/uSazp1R3F5acSrLa972
YSzPEaAlsqInVYSQMxRUX5nuH7UycZG4ZaELL7VPy1hplM+HIQnvnouvrHKOOuN+ztpM+TlQcikH
NWppTDfARGin24L4f6bBDl6FG+iJP6A3rZIwhNCewCGzGMJxCa6tgOrlX6OpQOhvC54Lb0LGoMWS
Bw0FMQu6tGroYrMw4ApvoJHNEEhvpwxlOaUL9Z6pXVylzmYczkwu4JC03gLkEpfeoDjuYkIFu8Z8
P+j7dXJzuCOT8tkd99xeIzK4qF98kCD3kZgsLrZV23as8e4Tk5umNt1siZ1kZWLtS3g+nbSv6vZ9
3MqrMlUTvp7vUKgf6D6/GREEQW8ceFUV+YR8LSup3gIwBlU0iK+kgymXWHrsTeMdVGksqnVTcz7N
r3jq/fZ9KcxEulMH5Jnsl8kqjA+kEVCqJrOIG9Pk1eyl5EBSUb3ZLpJloJu/pynkFrWa0cQ9BwxQ
q/RHdf2FOVpiONYh3FNBqIUc5pafm7wLNihzC++Bvt4ntEzJvcOdg7DIDw5cYD522FfxtwCsmcGF
813jCpRcUEbCj7Q4zlMhWyc6JgFAZe0Np6Z0Qt52fvyUzVlKTvt++zs4HuRKhPVM1M6jQmet5KQ5
1HN2dJEfkDs3iKwIOwRf5E4r2H51MC0U+BsjxkAGKcojbIA3mPo4WMVEoYmmkjWQ/g2q9EiJL8Vh
S4nP6CdfoGWI4r/N0lfJzRaJjkXOzlnz5hNdfw9wA5hGLlR1XGVoko3Qfe0rTBFWZhdQ8+DYQ4d0
tDDGRaJRfzzH15RIbhxOzGwoy+ZUUOIwkPl601bvzycfkN1dPD50WfJOrgNSdfKfwN4qWLDHO9zr
JxTPSoef6fLZLituvEX5Xc+Y6dXDrGCPayAlQtmOZjywU6u4KCE9A6S1YSfkgGGeb2szPo9hZmNB
WBxvkQMsGaGBEY6CFHK7jmrHoE//HhIPKxZISw/6LNS2cAEPxlC2/sgBlzWShzQ+Lw7qRIuGuBto
YiX1syZQQU6Pv8YlMJ/ODcwcN5kJ0zYQxHaqPDYZbVX2m8aGClkKM+PYDgTqSPr0e2GOs1725w9g
yYJgq3pQicjXZRJPy25QWCovkkQR/177+qq5GAMj2OPStP0+nMDR9imLlCI7Hsgx15uuf9yUXobV
5GG/F/kiGToTdsSQGzvZVPmSNnGi+mWRf3LC9T44OuH99yvxqAffsePHGLCaHIn7lbIPjmWUtds9
Y7zKpRI/u8KDEPVZ8TWIblq6N7DPTjQVFKUu3I3dhak8HENxcPT/DxpwRVJ9YGk3fwW1u5Ge9ZCh
oSEgs79GW+ID49GYSstJLdr4lf13PHTuTuDrmBtSgicL1EnCGKnUwznjDs+1BMi7sI51cO5qn+xr
q6rRbnTNWtjBnjkCcaUj3wFVbspP6qvqbeHRtKQSekR03//CNndGMEk5zACBh/lAE+SWV9vGaaI3
p76bpAwHGOTDZrWQRCN8u2F/tPqt3c139V4qg7VAWxROJbmuqbPDVNSNr7Vq3DVwqbUzujjH3N1+
LdyGnJr1L2E7t5n9yXgZ2F+sB6zbTENEeI4pwgbJUvpaRogpRpx8ikVMVS83yN8Zt/o1lFjy7hG7
aVN4sbLqgnzTVKrFcnvJudhhelFPPXAxrr2dNMVjSV10Q5WTXmJYI8nPcz8LJ8Gkz6H8/2OZMgNW
9q7aU2egjj0ScPmosDS/teoF9Oxm+LKbkj9I9wq5sUQkOf0wHLm1fNHkdCs9l7UFxjpc779HNmNx
Lt+oDhlu2WO881zxCGpf91PhA3z2PmbhjP9ilk/zOuKv0gmDIS7uCluSbGjIM/97VSZLPurRRyuA
WhGA9uqRUHqBirrkLa1/JnEHf2cWtQH7keViuMEZ8OrULgHOx0fXtTCktMgPn4tDtaXlvp93i7GE
9YkquJSOlJtRAF/hkHRRSAg7GSkw5fp3N//4JYocl1SCX/oZwhr45dv2lfHqz3p0GvZFDcE855It
seG2DNtOq2Ju3CvzZAKbBBIPk7hYDuSkzXkFp+9q+8Mv8ylkDEn0IhtVmCrZvSBQIeEZ5uKGL7Hu
BQ3cYk9wC085LTUXVy9EQ1ma6pGsIYEkbn1LCgkvBb/jxlcQg4RqfdX/MnVMT264xco27JM9Nnwv
FIG9RrHLenr01YE7QjdkCoB01BRLB3IXgq+1kno+mo3qlw82U2YeSTJrkp0QzIWZ89ea0mnB9AGI
aHiGCwJd04a7+k3FqCGsfpXUD1YgXSy7E+O4GMpw8IDJz4D+IstfDlLoJKAZ4qqjYD/6w4I5H0+R
B4O3ByapIe2tnSO2DPrLIWPzN0OjTdc512FAEyi4PfsyE3PkmRG/qNgl567lQD4LolVuxM/bbjYZ
62IGeKi84gd1mrCSrLYMXWjINYvSsxABBhKWWeUrcbp3LvJuqykimIEMCIOR6LRu3goKKlQ5BQsp
N5XnCOlh3tAgCMXCRvTAnhkC4PlKWLLkl6fyAFnC6cKPDs+ylq94iNpshI0uEwBduqQ/lgQZtNFW
FHx5F4WgXqclqBiA/wsuQE3D/vKdotScx9un/q/PvBGqVrVS3VGktIJpq8dY2Gma1ANmU8E87jrh
+cFN3i+h+RbgHwJ70KdmM3rYAmMLStboUvi1b9PgyvNZdqBkcvhoneQ0oDT8tiEyqFhG/zQ3W6vX
A/cUF1kfITqH2YSbCDb0tpKmMHQ2aC3Ukg8AK13cY7Fq2SzpFWvr6eWGvtlMwc9ku7GFEaK0nze1
wtidmV38aolGDqffWepXuyMDD6JxRrJp0p4bOe9fO40iCiDeAzU0MilS3jWf/+9Lw+UjUhb9ITWe
LZLXokAUViFDZ0p7VFzDFfjeUXp5P2CWkSSjeBu/QwHVsMobsY1gCBMYwuvwAbj389W1Fh6uhVQ2
T01OhybzfAF6QondCHVc76+nuihvanUoij96sbC1Ezyom3Zz/c2exq4Mz+bpDG6w6r6ivHrGbMwM
A/dc5MnflxG8rOPjFcQxJNU7Q/HGPApa3AcLaeGdpsuOJ90dzYmIEubjUMXF4uSYsa0pugaD+God
1BbXAw3XoaeP//Sg1kBYv1fXup7xUkH6AraRWX8QWrYtyNL/7l/VslaApeCaZrnEZgrUghV8kELU
t6P5J52p0Vu0r5KSa0mR2Eh6M4trAkwbqZhh5Tio2vUYBoNbKck0eUgFYN+9kg5AxKfYyXzCVzqT
hqxPdv2RcCMgRDM6I8aXxZmYLoH88OGkldJL9VNTPXooGawhLJ377zLSWiGvev6q1kVowflW77J8
4Q63MJPvBzBaAmwjXLjvpgxLHR0zkpaN/Vb5/xdeWvd3fYhfRT1xih/t8wxcHz85ezC+VDZ4ifIR
n5JJtKHZbDTG//Y+oc/eYlRMMTDFi5nGM7v9rI++3r0vzBDwAXVadLeB5ZBL5fD+OKMN1ftKLx/+
r5bTBnSuZLaac42KBTfHLXqIydN51I3uZwNA3Y01RIrL8Vu2p+LBXoWqDkyIgSl66jKUCKr0XadG
xhub5KsGMUq/MeimqXAUGzWplEqj1/HNadOYara0piMfDNVk3APBpn8hbXNlno2MqnrV15Zy6WfH
cr46sWrHqs/xviFBC6mqDdHjlbuKmP1eZjlpBp75OYzGmh3ZuD/M5+71FXUmbNiIkZh5fWH6dQML
AUYbh3uI3xJtvX3oRbS+gEPof0Hjnpo74wPL6YUVNSUk303TTRZwm/lRHLXu5jcseHCitd3Am7gB
aEh9u7NyojISCx2hIlmvbR93cqk84+eLC4YXXpNH74K+Z8Pf23FfHB6WKFih6fSbsDfjb5NvOawF
DY5OWFct6wn2Gs98IZ8UA59pwAZ/wLWqQpzY5cm49hegPQZE8NFIS2IRQ3yYfDAhuD74bpFyeE7A
s5jf3/9lRv5AOZDB0ek+W0OGiHDRWDlIbw7SXfJlBxWWj7kUZWn0uiAEdMyudlek7GgSjp7WPeX1
6rUt7tZHOeAg93Viqd95TPBLJ83xM4h9hDe13SZpXvhNhWyBMXvAwQRA+rdMbYmgrAZr4AJ78DLH
PNhWaHDKDlEtKTlqBOIOnOJ5VEOr/VezWR8mKwltHurAuomQ+Zd+9mmJKEoKkzKxQ5AV/6vUvt3O
xGr2V8qMl4o3HX4dECdRyAvkbKIjG5F1Ct1BOTHv4rGDVrsf5Uc6vmMCWBOQ2roYB8LGOsVwBvY4
vn2VnGdVtsnjAliAu7NKILrFhalBasECmE6wmUw1LYTE7ad5R+MSQP+m1HgDnyGXLihl65Gr9IDB
H0VXdrlbhfZBs4TcON9eIW6e1rZRJyrAdHwKWXKfJt3BjueeLgInkgDzAAz6DHFXJG7Q3/o4+CqW
nomvo9bv1hWOYnVCdRkZVdvDmoMx8tXE8l/8NOaHJrSOi5paZJF9PHHwktuY4AEVjJuhnmM9Y7nB
c15QCOsuJn3Yt6XFMPkzUF6r7jthirjfD6CFINJ1L3XH/KKgtnh9uHDH2c/6dBIDeE+0/Cg3Y0cB
sXCUVi5eD3Sjrx8j/LZzOSLqbjXcsjrFXYOfhBqdxLbJQWWYXTcik1qFtH+Tj6VscG1Skk6sC+99
SKxh2ULi4TNhvLQmixvuj9Hhx6GtVWjFCYjokbAif5SzcDlbHgmdeZsO99qQmTkP62wCPSLgk3dY
2sxmm+PhLUK/uYFGEkEQkIw76otX6Fe2jqSIx1RrzRXRL2YJnwfOFNfWCwfEF6ZfjDpMtNKGGAVO
UCfmSGPXQOMmEiUzwryXxnWwwqyL45fCk2sL6rjVXjTEy9XtTI0v/lX76GC1VS4kt7OeJoQfzVmB
Zszfb0cx9Z+qf6PEbgZyjEQ+lSpomwVWw/OhHhQTuMAXY4VURO0lf9DF+Q0619jrxXw8CYWLTQo/
5ok+nv51m3hG4lfA/ef3S5+ddCRfK1T2yL1PDPxS/E2LxNfVKS5vewNy0uBPrzECX7Ucy2M8RkPa
PplyVaxQmGylOrvbeVFjx7n3fOSTkn7uVQXXG4inFgDmyyvJ6tFR2OWwtUsQ70rBplURQJBBWDUX
M1tuKCf5LoFTj7d0ikiGQFa6FvcKoHDWpvaM+0zk59cZzdwmDSPKJChzWYOAguYs9bx5GAR297pS
3UqAJ2xO+2onvXTCk/Yi+VfA+i9Y4zSPt6TUDE+dkRGhI64NWmX5nFFzjhu2vV6S+zG4sHZpLI6J
rjtZ46oetfO9x5WGDTQFQRjqqT87x1x1KzSDGLsd3EFyIaxKjiX1aLfJYafcZbRJhHPzWtnLcT2n
40mdZhTTNauZO3M4WG0Nmm3jwxTvxVe0dXkZ4310D8fhZxAMT1gaLBBtTgkeSxkDnunlh4Us26Zo
Kb5WCXPPYk3N7/WFQzNwN7nEtrUGDNA/pi/Wwsvgjih0/vTIZWi9oU2vLLpGnPTFFCZC3LUtFDvE
Cisx9PXc14K7nu+rejAaBApm/aL3NL2eF+f2jvHOIYCJYkQ+IZw9JoxQT7m1K/k8kTnXUNciKjXp
MeA7OwnjjIuq8mREPMoS0CLQm90pDdfMDQfI+G0nVJiUHFment8qrhk6PRtTEqaE0xHBZpLOPG3A
W7yN/pAHzhacTTyaDYsAG/od+rsYizL82bgQxwm7unGcXXA6kI9asV6pris58Q5ytRK3XCuaSDO/
C0Lb4ffYAkD2I0KT0PtIeEHVLh0HWZPPHLgOn9XzSe8n7S+j1mgL2C9TT+jdZO4BtnGG68LSMPzs
O70o+0X3eOWvERKs74SF+Yi2qj4ikS7/3MaKRCD2ijPccFa2jR3su9cHIIaS0elV6esPENXUhEnD
eX2AMb0i5t/oWKINujJALBYCd9L3cTfPPIaY3xM2A/GhKQ6axc9jHju0aJWQY+r1VCBAOBMIjdI3
qNMDZLwZSZwhdIH7w2o9Zdt966izbpcmzuRjvmM4dveS7bcmVRDJWTuJT2D5e9Pf/oRLnFBZRKX8
cSRkr2tatBOQDcUa0rPhDgzM+bHHOW73P6yO5iTcczuCHjMQ5Ue01U7y6OBpoxEc8qmA0sQHwONQ
FyyT94F0uKGxwN2mCMXbqGE1eQhC0nYDyaUvYhSHFAdarTMnPj1QpzDcEP2p5z5UWsHWOkxGEDdR
+G80Jz/eHL+e7ekxEWVJdruYtL2varyYLaZ9HLwWnJ5TfB5n3bwlG+LsBHylrKdVOUtORYTnzyVb
beY5FHm/+dZqrPICbT5Q0gG8mxKKckzv01XwAtua4avf5yJJH7bpN0BnNe/5MSzp4RjfbjP5LqiW
QVFccHldoqjlf2zSmfSEr6VudjqP1K5EBNMO9f+p/LGgc24czIOFws68BtM+fW+wI/WRZGW8FTFH
YYqa1Oc+5Bml6YlT6zjC3GaYF6XJXOTocgXq5K+DnWNM1H+sv2m59YPpsrKXFhl9moYO3uo5t2fz
ctJmYTjuZB/njU1sc6SWbL5Dy0nOlnbTiNLiZEttg7Yx/C7gsROFJNjRM0CA9NljWVPknf4hNczs
C4bcNqD7f/o0Vwh1Nt95nUAOG0upB8QRRi7odTnEJylmdPfNu6yhSy2wBs+hXUUwiDXLgfEOst2G
VCq5+R1m40ix6/SgncwkMin1Ko7cQ2f94m5kK7BxrkV50BoCn2NEr84ym7AmzV+90QzvqJj1noGN
y1upwsyBm+5/QhPtUUal6HZhpulfo3ZQjT3YL+Hdt0ntcOH4+nDbipshfzyXRPUanuJqz6cALmhI
lTCXtHue4ZSRoY1gWZKMyvZFGeol2/sEc1/DGwO4bt3Z4Xa/N6PelAd0RDs3s1+jiQkDATBZ9kBC
hrr/hn0zQBirqT3iKnBEsl9DCI6A9dbIRquAqBSr1UuI4WXaaXCEtzJgrspipoy7fSjO8XgFSfoa
d+JxiCiJRyCAGMz80Rjo3hjeVlDpGDZJfI81T4FK874gAJ1feDXMWuxf6h/vwt0Nybr2WWIRN6Ul
B4lphWwZx6d0lBOaEu1ES5LtS7/vhAoEDdNqWHijSIPpvUGmVNNKapQwlQU0Xtf3ChBv+dGqqIEb
i1YkJIVcF1X7ZQAzU91ajmJv1REmtH5IKwxhqHEzSYoqsIJm+jdTP7TktNK1KZ2c/Kljl3NN9Ds1
iRVdtZWao9+GiHAYF65KEm1D4zQzk6HxOhzmdzmXKDLAXZ30hahrILt3dwIIgQKGRXx0EAxSQHkn
pCJv/cktiOlu7sRwY5/pToQZ+a3PoLAcxSScHd0EliZV3JzpaGFTR9j82YT9JihUPkCLVhMmbPJi
F6CQmqBGt3whUjyMjFBeaLxHWsXrBTirHZ60BFZ0xLM/Jk59ea7Nlic0Y7RkxeEa20dy43EcKDF/
5ULVAa7sCyoCy7wdpRyCXup2A1mWkg2HOEggtbMSEmphwFZTFY9LWwnNWvH7Kikner3FUGX9Z4Cf
dGVlsvR/cPehS6jLeys/vyy1kjblGL59BGXKskzBRQSxMnmXtHWAwN3S5KJJQGsGHb0BUibjrWha
n7de9SPWQratvRDyFjrTKgREV7k51lRunqyOzojqLJv2ZNnIBPaTyP7CNZWdPLPRM/42FfQm8+LA
noq7OZ5eFN4oUBsUP3rG96jxxM/rs5ic/j2sEE3UU+98HctBx3P1bmjDLQzjGqK0lJ8jTGkqda9D
NFam90S/jEt33xsAzxIzGufuIjeg7NKAoB3ErHzwz4xZ/AE7soOUlg4q7IBxCPm+zHHimF4Fztqs
AjEfjAzRE4WPwVKu0mAnML6MXZDfV9fizQTZFkQwYfYGgvj2xHUcfhnl7cea/gLRgV/uVoRBZD8R
VykTZkXx3T2oG7IULNyg6J/Fen7RERCg+P3MOlNh9dGmbC4xE1b14kip2VhHtcrgEsQcOlKlWUUU
9ow/+HrW7eUjXV+2DWy6FawFY0vADqAcn1zo20bpw4Pu8l2EM1GgdDaMqW+68xzP28YdzSqV90ub
DCY9FGQON8FImU/6h1Vb6aXCeBknKiJHewCGLKhcmfv23EkPkBBrXw2zWJkfCbOg3HlzLPIZB35K
rcU+fatkggLkpUXZwvhZAsUDS4rOa7PfrKl/YIPRlOGk3/2yDVEBnUnQq1U0fgxPXO1VYK+NcG4l
/TnU9vw9HAchwaA7W/ZFA/PuzvSy7dC8q6CfMR26q7TTZ7tqaDFt08cAa3l59FJ616snxA7W48Vz
Ppi2om4QsL4p97DWUzxz3VMrY14Kjx42FjtzWGIP2/9auzxMiBkOG4/mlF8WUstWaa4QgNrJR3eu
gXfybpSJ3rhDSrVz9wS7PsrH/irmEyzcyioO2WGZ0IZfog/1kwAnrh1c5WPCelX8BaEda3dnukVp
rjDbayeSGCoBHFUx1VMpnbrCcPoBPoB5C6+w2HlbIPPYGJPVWF9AREVcF7Ckhjh9uWIcO5yaucEJ
M2MeNhv1xsTBEZ+cO+wpXD5etSPC7KxNtV6h/2gobEAQuJyB7MBvb54Ogk/0rvbvvZPm7PxWwnII
Kx1HgWWgUEZQGPPtlrvmLNar49lsJbOXR3mqF1UBEmRV48xtQO/5cD0nEev+L/1F2GPveg66vOTu
4aaj5RWvAVnNARnXU0tG26Q7IEcBR826SJWMq9eok9A1ZTmEoaHbyxW4t4iCV8wyp2hWopO1/HWV
PpIGWW8dzr3Dez+bE5iWpe6WnQmBdyRRx9tTXGNN6OCFf9MqN5bpQfDmICzBU0rMnO/Pv00bBK8H
34qTCc8GfY8swIUHmdkTL9Y3wvG3XMSKvsNMuSa7Pc8gA0lPKyISEVY1BreQBSBZaCGBp7yQIUcJ
48yRx3lQq41mlL9+6+JK50NqPhC6iwpekD8sjYSmBj+VryuG+9qDnWUFkkHFS6Os8gf+HAvYRBzd
1cO1tk50QRXqE5dSZuu6tgIwSb/QEpnIbrLbjeTHCJyImVlInfcdJrxOO5/pzABtaCALo90zoTSU
fb54ZYpV66Ki3esSO4ZAayOwmQ0e3TYAVoAvPloaiVmwlQw5lpjf+QCmglmoRadRLX+tCOFjIvAU
Pa+WF3WQ0k83ZytgEaiFMLCERqrS/9bPaxrJcSdfXphVTrCJewZtbPuoxn9RYhNK60oBcp9lb4fH
uAWZDRKY7Mc3R7E03LprZYgnrvhaU9lYL8oiKtA/Ufp5s+nyx5rgfUsgTJA1sp8vWu4M/Vn7lxaw
uAdj2A3tnuCs0rRFcc0xs3xmw0is5t5R74L4xhzQ6k5Xdx76D8E7bqZuxTqL5tJd5+Y1QP9eizUJ
OUqNyikQxQSeDqPzuQs3iUH+nMuLaqm4T4dzrYSn4ADTX3MPvoDmwxFdJoa3vZgXyt51QbfMeYA8
cLpcJPlPVLsgsHmmeO5eG7hXrXqwJHRKRYNimh8SItA1qyRLwVH+wb5vlpGjmiHhcC7Rpnnl11vS
Jtadib+rgu+pL0jZgxEJ/hgCuxMQ8eIeWF1RVET5i0fyfV/1ui+IWi5ycmvKbrDMCzimIcSrl1Gb
R0I+k4VwkNt4Q9tAtBfZUuSv301eFcD/5hrJOyQat2FJDyntmxtELzEQlRFe4jk8lIDyiti2X+RB
1ua3zMoJzrwKAQO4BhWSSV1Q1qXZuXoFUEKCBD4wqPU1qH6PpPxGLnitvGnQPeXdOSEVbZnR6KIO
hKqLjHjnJhw2EvLE3D3YGZybcpHdsnptQOcdIU1kILevRQXOBPe9FJjAR9B4CH3dKm+XSKuBdJGL
eCgTWvp1sXAHRa4ehhR9J5QtNM4DcIjibgGSmz4xdxoJdJxKqPtmkVySy9jPdTNdmN6z/bhhcRPF
IdIzKUOHIjRhec1YWAceRGVfLTAcZ5Asc3YGST7oR9hoZReYLx5Pg3W68VDPI0/bB0ukkFmC1PmY
J9VK1ZUh+XAXj4Z/UbnJsBSU1f1HmGRvWtbHlwdPOgZDa++6DJFGh/7AOVZAIWa5GBXy25WTSSCJ
NIDHW1e2fDln9233LXIBoR6JWtq5Df9bJ3kRE68l4uyvtpO9P7heWSX1mpOOCSUIkF3edKShRQm8
8ewWzLdvXEicIw91QauKLON0IpigJYTOO50g6SUDaR/9QNeWs1jo+9kw7wtXZD7+G33cQg4ciPOg
rgfBJCFxqVjD6/70fJ0shL8to6m5NwepfUagLA7slOzqiZV8SrEdmi5I7jMex53f3mLyR4CwUruT
SafZdruaU6J51W1oqFo87v+qKVcWfVDUGBj9nqT2XrqOAgLkGfRv9iuYeA7KoIx9oDYYbFL3HxoC
HRMpWCfX6oAT4ojPZh7+3y8d5rMJZR9d4piTVnaWEX8qyQdY1AotBj0k/ytWf7oQ56phZlbwpIzQ
3PnIMb3psoB21OisgZxwx6T1Ww3T3rWTdP2cOk+7lz4dpVb6jgTLv0COLFA26gJX1Qnx+Vys6/+/
D7OJ38DqOQ/lKgpcYkPmJx7bx/ir3XORcbtbkZhZR56svL77BNGnpk6h9Xbq7YdjGyG4iAPOHwFK
epKjfDNTEfFHV/du6TtfNkxvaUItZ1Uu6hN3fNUJWtI1zYtplxd+gyfEDlKEnss9orz4xTGq96s/
SOwOzyP8VhC9I3fu/2Pb1Vn1xgsRWYK1/7T6wXLjDR1kpt2LPlf24eLSlglI+iDk0hgqZ5Vph5fO
dVcF4zkNqouXuaF96SvB/hvRJo6G/6gOZyLS2VgSOiA9TcNAlX98f4Y7KRqUsTSpP2YmDtvnTC+j
dVLQVAqZlDMZBGbBYUU0LXWR9ewBU+FPuBRm9hL6EJo6pc0M4TWy4hqoNV6eis/2AVF3rJ08EK2Y
7mY3R/EZHufcYSsy8sq2DanKQz2UFO4uoqiWM0cpb8pcW+O2zeGFK/Ywh6PCTrpuF9rFENo4S/P4
VRzS6itr+BXKUr9AxNZWKxMZZ4u8IHwqRgrUx/9mf6nsGZb2H/OmVmlGzdJYlG3IDrUi9CJ+LLL5
UIq7IZPNANTTZLiWR0Bn8TJNoTsnpLXtwhtiU3HfvScarlukNMV8U/LipqsIHJMSIPCl2XN0XEuo
HvTOuVReRkUA9JScm5xFcAe5qV6IHIB7LJ+qR/obwmSLFhofaq+h0ttYWiNt0SdX/EqsZnk7fMMT
MCxZpQM1vJAz2ulK00k1iSlTy/2BLVn69AeVZzcPWxheMPTxS06Gi3Tlcf/ui9US/9F3V/DMZxNS
OVZ5e65vlH0JwkpBpKlu/DjgzEctKwxV072lvW3QoC0ditiAbSaWX9mi85/0YGIcnPNyAoaf12qw
ai7mn4eyoU/ckmF1HlUi0D31K44BwdbmWPhb6vKXyKEwOm5QuBk2KMgJ7A+K2d5PtacvDTLJsUUu
u2FFFXTjb6UEttxGpK9a+LtvaRdSp52wrIsDZ7AutCEwZX/ImFKjjO44aTvd7SuwdmFB/xYQWN2g
COj/BEJTEMlWiqgnqasMWzcOudAwGRd8vmo9LCZCw6FsZFsVmrL3DGPm3UGOdCBwU9+G96KN+Iz8
s9gjK/eIHfJryykw4eeKTbDlNZFZVTVVVIdGlNP4y3g8E6dsdHmWEoQ6dzcy1sdMRizwkm5Bp4Ia
I0aZc4mvswziJ7wSoUwe/HfB8+RAvCP7QgCBtll8MdA8LGUs03eG3hsmQFXJ3maV7+lagfTRQd73
sc+eo6k0iwYcCIoiFIXkBFgZ7c4d7SV+YpWXyYmOLMnHZ8bFBECjUVY1z+klNA0JejuWLvfIsm7j
3XQnIPyoxNc/2HORYRdbASgaRYEhrh/cyhwdnKzIv1R1xipW977iHvQbUQXn73D5c8KY0ss0WrCT
fnSfvfvTUUvTl3fxwrL+AFt3gREqOrSfqcC/UCawXeb88rkOheC7S3hPvVy9+ZlgR1R3d9evSwkr
H3uYFLRUXJ3uF+4K40dahtSkIrpdwAmHtQ9dny4wzVmSK39TC3BgwtourpbDr5hRteLPmRU75765
vFBPPsCSS1DiVHA3ZlM8VoMXwyuBt4EGpB/t8b319r4ZC9QNaCzbb1IZt7CRSCxKs5rMjr/O5dXu
8M+pMiG0Z0AgUu7RGwaXx7dwpkAlevXIpF8EaRpeOSMGikxX62lABz+HILoFiG8tdN286fD69iYZ
CjAGV+fxlamM8gGtWwbvpj89zOeDlOQa3j0FOT8Sy6beOIGk9LAIE3Z665bTC+3DM6heNVYr6KRA
5R6hUYZqKXOpXL3MwOQUQRmHaEBUGTcIZnfo0zAPWbSv3GmPVhw/V/pTecGqIQRMO0u7LzSvLaxm
5NLzEsWB7l8kTJ64dV0lg71+5kYdm0EqRW3kaNi4lspZpkqC31cdbxPcenP/GifY9XZ1JKAoLDAO
bbfhLSycPdcembiB6qYxrk9OXv6jBzS06nafWrl9pPUm1XRXuzpeBgFOhpMuQTHrM7QI3h2O13TI
eOnZy8gIdMGAZ0zueVJpeuN6eDeki5guMkw6uuv7hiqlj0lr6D6luDaInSKKpvr5GxKPZQVkYWi8
iCNzH5aDHxv+2bRmmoN6VQsgPmJnR4cKXZI+uuM6vEu8DdX1QGscnYGZxYiNH7SrVEWvZ4Z6qQpi
eURsB85anDivp9vtxuhCRoi9+H3GhmOK1qiLgP4MiU9Kq9tGRvGDye7PdVuKzIJ/WbPhhYdV/ImC
NW6oNiMWcGeUP63ajFQFJ79yAKsenQJYISmozsdCDa6p4fyclZWY5hHS4hyvCzyShobmEZJfPEun
sU5M6tvTN+0fZitx7F8+rUMUXMXZdXIBFs9MBVjAXMOM8WMWEoGAycOy02c2+yTspuSUfMZJ/+Id
knY8KLEJaqDd/M10qQXdhPJADfI4u/XelCxqoj0XQwzDfyT97AdUCfHb2/5FINfADbZtUXhe0V4g
+77boKWRmeTod6SEPM+cZW2k65R+iZA2afEB4Ks1AbExFZIhA2rXFrenWjgaDUWo+S46221Nk4+T
fr9kbhjCxP8Nn00jm1eLChCQP2SidJAhnqiOGsgTE2dcitOqpfES6vD8TEV6H9g8tFoITFLuUHgP
cenJgXfuRgZAYfg0EbXyRLZ60fl5Dg3PYKITDMJlPfgYlW0yahMIafTGyw5nfkPy6sU34hDfPt7A
rSMsBSR5e2dMlAnfMNxD14IMR627KacL2TNpn5sYHFYMegwZ1wHspmuTMNwKUUHWTfNLNpNqiUne
S86fEBJSlHuirAEJMvxYP4aXvfUon1O7gHeSlp+864Mg/ghC5f9b4qzjKP1/WX5el9GGrvXgqjg+
PxqPaVM9cGetJN3iM7HLfRzmejbaLOn+zkcFbc8hnaLnmxIKAttlsung2IWVEH9NadWcsXg+crlw
rSxTUPXvwPa2hxLcLFsLdVCnJkZOhTK3xM6JbCSj+tjPuZA8gdY4M97yU3sAW/RBuEGU5eURtjwY
3UdymBQ+uP7Hgn0D4tJKyxmxA2sSIZo1HN8Ut42fFwK3+tOopqo83QmA9WA7x9RcjB8jkK9g/r/c
QMKjeWIuzxhe0oswsAQuuVH6sTWRu4tpbbgbQxpu71rjOYE+02UTn+/KuCmc5CT/0vtlc1NZed3d
/4QzvVlklVQwc6+yQD0TkQOgDNft8NttcRHzoGxA9JAiFjT5Ow5zGMtcL2bA2QuGTjBq6g3uxMIj
I2iQGvP0lDM5Cm2FgfZOmEQko7C3oTN6JD2CAbdHQWeSn0xHrBkqNuyo9OAGyBi0LNarGhHbB1JC
WFnUmotQtqWcvvkDdN9E0N9b9z899kcnYQF09CKM6FPpYokEJNOMgcBH+0QPfzVB++ugyFogujBX
Y70kEfbhAGBp+28KoXwDatF0Mfdq5DeKfNoAhlmoui8+gWFg14uUsOO/2oMMrq96O/pOFxIxdiKv
xlPNSqqmPADNawNVJ2nM0uHqnNDhxwe3fsUpVLKvMhQITE7MAM6RdT4xjS/B9/q18bGGZhrATfWU
IyULitsq67xLZ3VI0CCRHH1B4WGsElF5UIXb1NEnix1rXKgpDjh4cDe+wGt40E47+jxro4pS4X7l
91H815o5BQ/Cz5YkxHUtMFReKrS1Y7GclDyB3slM/bl9UA1FkBLScJpevq/RDfV5HRNk/ZSRRQTu
UwqlZ05Sn78UbyJrnzzmTQFRwDQcqUTa1+zkvuwD/nejifUd0lj4mbM0VQgd5qJ2UtQVkp9Y74ga
ynKiQx2YsWY+RZobM4nmugmpPcseQkV1Z8HNdtPXqKQOOqtsmTqLvwGzjtaJRnp5NNWK1e5PuhbR
CpAgWDNslQAAlqFBeMczB8NKmC9iKrvhXcWfdjT+9iz16n8uwTWsSefldj7km0kOo62wbUudEX+0
EPQq9od5VhAJMwh2vBNqGzZvtTbyP1PqdmuSJBXG4M/1kprNFenxT4ohP1XLV1VD4UPubjjZiLRe
Y4EliG43aCysqnAGe5riJKhen/R7m3EHfayrzCyrRiPuqrC+c7HQYRE5CYSyxEMQiE1N0JkBMt/i
3kurgo2gHkZ0YhDbbNVGTf8ECwrERftJMjlSQ8x8ge/QxSHsHFnFL8AcAzDe6Yed7ue7jmM2J+aq
QnmfZNkUnuURGrEsVTxkjAH+dYZYkaGD6wDQEWSNIYdDkeLQQ53hFC2CP0rLM1cIZgbRgfq24d5L
xNk8+8XJfpBC+EkTKQAzUBDPV2Kwsi3PO8NICk2Hi9NMF7Wqor+qBhkWDHFxCbVizJAH6czbTGTG
t9kxPnRmI49gHEGiz3eUTaL2RBlfpK0nDR3EZFWAs/i+GuZ+RtwOKOIabQ7JZob3xseeQytgECQ2
3VTqnAaxHBh33c5dzblk92nuk5/0Og+/6FyLhel6AVPokWPnnyUzPH6svesW0vyXIqseNqFOYlsL
ZAYTKbPPwpl7Au7mi5Tk+5b2Ku6te/8cwYdaMAZhP210ly6l5drjx+q0CTfbCuaOBVkG9VArupz8
SCg92zF/gaundyQ+SYBlUfpTIoMBypakQdJBd9BTmk9krlkdcFfLJ1Sdd4eyu/9auxm3RF4hKhq4
A06Nr/yoXNzN3tmhETcPcNtthrxOJp3IOpSGpwGoDzPS0fYxTBT1TlVHF6EvHwJ50sukJrzWktJN
XVrD1BmD8WT9fRQ9mHd1RUGFW1LbaS4LRSo+8t7Ft+gzWTqwek/YSVOfGCt4EXW2Pd799c0v9i1r
wjEFmrAivrkxLo3S4cOIV+rT54cy4ALPqyQOvbyHaaTdDrpRmWarePQsGOel2Y6vGUfcHSetlVOS
87q7bXaAHYYkzQQgkFtdw3gBgsn1m4nmxi+k3LU+cdFwJj1nXbVt0/E9bUANl0ZdupoE/0BgWa3E
PCQSFBJfYwsrgGXWvg/PJev+voQytrxig6XqOeQDD4QXYLw6t06+UZ4Rrkz1YcV/nIZ4rKl+7DPf
OvNuB78x2y50EJpBJF9g2tc8Vg4tOBSsKQkSdaFGLGVP8RWeNIHcI2EdJze/7SP1H4BxZq3IGU2O
2qFsxt1jBUAEOT9DDrut54SfUHiIy9HngaW8IEdTTFNEa8v7RFfX2rRGmhysBO6OIHQiN0FTHbVL
QZIAKub2D+7AHwm0YmStwdCMF4JvrKX0WAPkCK8FiF6yWizJziRbrg3fyxQgiKVqNI+xuybufQsJ
HvGqSm9h5ab9IRAI2URRgFSaksPGmuTQ1owKogKndxyMwkyHe9yLezpxZz5lxQl6gQI3fucD4UO7
0fSwEMdgvX5OvRGFThHIa0+AhqzsSmjoZp5aUY33l1h7SYoCESN2GJ74o8ffsbPEigCVD5lwaKIY
96nhFlXe0s6ELkU8e6nvqjQLoPfme9+iXApNsiUpQziBuHA3Bjhr5wreB8VM/G39SU8r8nKHqpN1
b+vPfoY3G+2X+kSKXI+BeUiLv3jQlcfymmUkxlQgMT4dsqhXcqLQrahLNepI8dDvRx7ExwHkkltV
VwvBROT1Ezu3+ZY/tPUxtqe5wiYDZ5FypQXjdl9Xp/pvsPGdl3eXAgcq9ACm3fvcZBBlcYE2rIJT
vvEuq0kGNanlEsAKJoX1kkvDlx+zMcGPdh7bYehOxHj+4h2geHVAgCXod/rhpAcCrBtg2zh50oNO
4LUlLz8MGL0+ZAj082xsWjGphVmTGBfg6LjgEEdWH/XHRf8jTSb5TeRCD5Gao6+enU7xtTK190VE
wAdQefei0nCJJ77YpB2Ld995TexVocwAkJblcytQnOst8SisVDoo+yRFkdj2baM0pC9eSIFURtKH
j3C519Tyv3OKX95wvvDPDgnb1pIVhhAkRQnJQOjhnZH1zJXyBixje8h/vac6GvWG0ggd9qNPneVj
1zKuJmUWWvaevuLA4/TV08F/FzFFP4USfU1SSLtbESu7qwjwtZFfMICR1hbe2CZTTJcXdNXurcPJ
/dyvr2DAxzq+LVpN2DtorYhV+p9rnoLjime6dAZZE/xBt7iMR+aDNFwbT4LS3qViI+FzUVNNblDK
3eerCFmD/Bc0UV2ZeSjYNyYGu/ccLfl85icjO2m/oI51dTaWj3Rcn21gfOR7N7ZHp7gJ7SxCi1LE
3mky1rFOCOggom1Qq3AvSj0ShYa2FB/s48fXPNhCTEdvsOfLOhwgrJI4CBzkvPthIJXUTYCBNOET
jleJ5ya3e4d5mVD8LiKD0p6sHxHz6jgPXSDTWmIJu3Ne3/AoqNpkB8HXeeL2yCGQS9emAyjZytul
sPE8pJDlj5gbDAUXSQrv1i5OIwAl16w9GnMdWJkhzT6knCx84EPyPDyc6HeeBgT+nvRQ1HABFpOA
8uFjPZxqKLdN6aW1IJWXGsf/v+xdshFnDuRLhWfLkB+Krxz+PTOq2gOYxNspXFLJX6U1TMXz29c5
KsGnghs5VPS3eDZFSRiTjGNSWNtl9li1C4af9HtuDGmsX7TehW5+WkEF/SOMtOEC7FfQQ/UgMkK5
XCue/VR2IuiWNSByGrjFftLQneuwwa5YnWvv2n+1hLjoZf9SQcvcdP1X50OIORVpThoFPkacQCqJ
ljjzW6TtyA7fJaHVx9ztkxmz6KTTf3fpXiQOa+dDbeDh0bF1PRlJZzdDu0D1yXNOcIibfZWfna9R
rT5R/PR/8MZZCo3PLA3U5aLHrjkqB7AVoorRpNuo09ypNoJbBgbC9Uaewt+KBGACLh9AMATv6j/r
q5/w8EQVagNoWbQ6cJyp0GS+cWnhW1h/TK9AwFsxtoadaN95kPSORLMdqHqlRgZMWmE5AS7vHe+3
X0zLLpoHLhwWkt0X+0KBYnN/a7G8S3jlMovKpdeeQvuAu+dOkcRqLPJZJuYuYJeuFSpbXvryaDhb
O363pqNFGc3+FP5yIW2zIW/FI3Daggv9QC63xdyRJSTGKUAJxoUGyrJmPQdhduxizV2luzYmjaBr
tTrhfd4244wcVOsIKusS6h5ceveeiULdQ1EBB5sVZ8QcS1u9sweMwrvrFJIoDxsuDVi0FJ5NIAV0
wf/t77tBGjbAJtQJupwrV6G3657BRmD1kDsArSJ1TYCTkwVWmhne4QtL/7V7fe3bmp8tEpQHwJgX
1DUFROguLpJxpJbMtMHooEeFBN7YiZh+fvIk+T5B/MpUNb90fldS87UGgtghCMiV0+GARFxS4dBK
h+I7gIozoBxMSzd4GXGf3TNU1dhu8U1Ck6JywfEVak/RNT8fCXExhP0E+M05rfNTu5jEfGzLEfIo
asLDAVvv+a5kwddXy3fK0EICit8epoTaWhzZuvKfOsbm4oCXN1JP6jDnsboUmSmLnuUhpvbCJuPe
+4mkNFMvX+1Q7f8EhbusY6HEqNYNoZD4Ue9kSnj6Wjs6572jyMq2dtevAISbo+YHPh3BoQS+gGPi
HbkeBlVD01h715MpB3D0jCevyB3zC5/UnhzPCEZnC7EbnUMmQRhHPgL29OX+8qaeS+0k719H47+/
tLnbQtT+FIauCIxnHEgqHRdQRwmA/qd4QBAojtSUM0WmW1YPK2b7/oQGkuWVyLoVsxZzm1/CKkSf
aepXS4mP5CnkQtOrHn87tiTHuo3SuO8XlP0k1z+y0ncKBXvMFlOxsIUBmVPDlbmv+i09PxKIsYTC
340NaCs0AzK1vZ5l89N517+wC6Aa6Gmcnfje/0I9mufAmNe1GpEhLGFhRMhXQGxkVP5nAUcXmuW0
zkGlIRFGRRyZZlJPV2Jgxs/j9RHfczE5hyjjTX7eMQQfewfJj0LG7z4NwKQgOM54ePu47QfCwA7V
Ps1NN69JoemIGprKsIgyyTBDMx99jUNqyiVg5k++CpIjiMJXz6P8P4HgfRezUqLWe8hHSES1DQDX
CErtdlTDJ/mSQ4NqGzktChdDo1/CpwE0ambDYwsUrCtZPYC0Gx6gKbgGpEl7qXSho324ETf8nW4N
pqB+1ZaCSeHYR+XEVHxEu4UK6bmK67Rsr5yJDmu/RAOV8D4YGcTqwpG2MlZ16mRKvKwdN6rtWFxk
Kj1B1cK8XpGZ5NfGiLDpN4ru3Zkn3pUVVXbaWuEJPZb3BNlIBlpjvm1U73MQBqTCZWgW766LkBUs
4oKSthIQglTgvZKX8kgyR1rSpQHmrMC0Wc1CF4AARhI/QLihTTaqnttHVJwCzLWjs/IDiFTVlCHC
p6Fetd1t9tWHA3wgE0HS7JAPRazRowx7+EJNTw67D5ze3ujx5yRasarU4M7svHuzyWjjZOdF0KT/
1MXZPRMVhxUzDA5cIBBhK5lKzwHwGk/o/esnReIpQaCfKysr88Ag/wYk2C3hrr96DKAFKmnmzPnR
VJBOJ8/ukV6DCiQXTeitQb2TufpZyrzjTU41uAKW/wLTHa/J+PbHXPbTBm98lYqvYjx2CgTkJ/LT
SLiWaXKdo71Lauz3ubBQpN6M/UheXEupD8DMuaAXvJIbVzT+wWDCTOro+k+sWeP/fPG71hbRvFO+
BFWWcJyXo3cuiVXTbwr+eBSvFaLiWyNTK2N0kb5X6Uiaa/JpqNfofymPmJURGtnQuEbePRgDMwfa
xrFdpnag+b7ewlAwBtoIMBWNP+JXDH5FtHWMeoF364iG8nOP8RdNVNYwJhIVyc6fRmDjsavm09ED
vA8QUn1rpmYUVDRAvkNUusZW9ciPefXTjK/N02w0hYHwnPwnoWLGTkuPrKgMRlgXEBNBPDa5SzZc
qCFDz2YVfoINHDqJDvUY6rvTen4+WWN0DECrakxKLHKa0PI5NrIgpZGQnscDgMDQIsY/M2IURcux
7BW4konWOWI3KmW0mbkIuoM02HL3IdJIVDD8TgAXLCZqSND3bcgSWJwmynR0xY7Sg0XGw2PFlVPU
X7cZpMstjawxL48oIId75zj89sG7O28nULFEcBgjLVnhBJF9F36vkHZUDTmN8Zx9+unLMKt82q0Z
vHcZ2wv18SglBzIKJzpRyfTpwJp1UTg6J6jRpkyVXznQZ5XAGmpGM3+k76KCK6qRJmgjR6I3CXuH
9BQPw1kZE1yRBndw7qa6c6kU5neOlaUQo+V3Fz69Ko5b9wOYFyk6T7q6o6+c1NOH6zMaK7FSmgUx
hGvCc2fokrPJHiUIPN3eOctk9gJfkadKd6RUVwXAdyaKFDkHysePkve79CXZCwuGuYiCfX2wZiLl
TQcjf7aLl8kIrERnEFC0Fw8h8ChWd7/hi29Yuilc88vyW9+cxDjBSxRK/9qSKfsY/IRxVZ5YWpG0
0/bWNIzBRSJqTcqStVpLdH/h9nxLzXJSYUIYXLX9soE4daDulUhzTb0vVfyY/juhEp1DOGmMglXy
ElhL181wD9hWrCMHYWFfUrRQcJxppNJiiV0D/AABI0cwviffbK9+2hzdW469mP1oUQQy/3lrgjGg
Kary8fvJkHQAKBvBbkV1NkvNDLUd8zog+0IhvZrFHO8g3LAWwk4gIPJfSDFcATHbmsASrLdvSbST
ViJHPO8Pb7nT99Kv8B0DkdnyZ6JfSY25ipd/0ouIJsGAWYf7ugvKx0CaqywCP27ujzh69xqSggNw
IRptoqxBy8sz6E8coZT3NU73s1jwn14mGcRZCSzYLNvnbmPcr6nM5xfdmBfZ51o77frKwSHGVg05
MBaLafF2pr9LuDbH4gXyEUjOBW9iiu72wKoUKxVxbpBYLrTF3bn1D1DQv/zxXQzIWHjy+G01UMvj
ahDw8F4Xy8Cgjrvxsqxh2IznXquj3R2zJdCmnYrI8V41K9YUBYD78Yb52BeT/N67s/9FLaK97yAJ
1rg5443VIjHjZw5B0xCONW/PoKDXTXmtESTzwLY2+/yOyKj/Px1xHx6q26idWegGl9xRfA3PzQJp
1RTLWDweJ3hWgx6VV4PRygXOZu1q2EGP0oDEB7MKAhNdHTjqTlIozzRgFmQHCLGJ555FfDDYpj69
aeezZS4OIJs32DLlBDUqy5tuNzFz5wNKCq4xW3pztsN41CfdshgJvAodZiTEQSFDlF3XK1gl3mYn
GQuwGnKjQ+Iv/JhH04wTP9Fu95f7601FFn6Zxa19XNunYUfX6EqiljQHJVTUplQQxu7mKKo2AP1x
CtLJ+B63SK2NCwwXMGE6WNBlYKRo3K4qsvuCGPd4VGR3Auu14u2pY+55M5Vcd1FFWkpvBbqIW5eM
Udp1itHfpA/6KfDe2+s4WkA3TuBpOVMJtjbrDbaH8GdLdciNsZnE/PEAH/TPVWwq0SQYbYK5CG5N
oozUFT/4qzxB08dieIV+o8jInyprKxIyR2VfHVf8IT6JeXy5fkwlbVQ2da8cj8e7+FiuIxQsKYFx
60AjL2lJyQ1zPJOhhVMMTzELo7TT4E4YpcP3S9xzIqrjYlNLDrABxvIJqDphaF/kwg3hPJ7YavET
SzFRSvKibVGT2eY/1WWX2qAuYWksvSJlnSC6cXnim/afi9ETblj6vehHxfSy/Gi+GniXNCbZZtvB
+qlrsnOolYg+YrIaFm2ykmVnHcFVCRNBXj5og7eINCEUCHLdV5aiCPUYarnAmvsNg67Zvm1CuG8e
b+HGhl0adcXcH6CnpSrgA3S9BUoJ/WXa3ssWYXeVTfUj7RtVLS+vbfAmWX/FXZotRhkPgBBTxFLO
f8n1gNbfbo3wbEt20lp/UKt7ZFY1mamBIPyiprgi6YR6jltfR7d4pK+YKOe3vdSku891IftCKalb
N84mJE5fUlIXQCRb/StPT5gJYMhmCOLkKIjITiPJ4GILEk0A4hZbKLeXWJZJ5xc0dP1x+SSJWPRe
HLHETxYIbVBYpRd6KHe+XnG6+c7lflQGSfihHh3prNUPgzeNlV8jzxrNIR/kN8285lQfgu5FPTB7
btVD8P7v/QK8yHpG2NQkLNRKZsYo48EIiJEmOIXje5S2dOPat5E6zpDGYo1+kaJmbr3HkdRknOLl
DZUp4V7ipaK4meQAaoNvJlVXobKe5heqjR96lk6cDcqyXZXTFQnh6egiLXSaVRodcsIWAv8DLnqD
kpr5HbMgOLX6Fi17CHndLFxo/2iHsWXogmV+TWt9Ti6SzPneFSTFrhwnvEFN9EF5G8j1RznmR4c8
ovTxtw36DjWJPwI5pgqAi4gUKKsFyqk8VvpXC+NB7/IZhgb4n/kV8mW30ojBENhwsDVuPW2tQTS5
Y3JsdSY6OnZZBxaBgyYFvw4KPicw8sjzIdi3IBlLjmyUDpaGvbWivRWjnHSH/z9nim1oblRIERXA
zvozL6BfgmxrbK1dKPyOHgaYcNl6u7vnu3nrKo6sGW68n6EBVJt9SwzQxs+Ly6QdYkkC20BdAvkh
Ok4hdje+/rFmjax7FZrc8cbjPIoY0FnLBUgkX9a1OborYiW1xPxeFZUb1DRUg0t2p82BmTGLXFhF
SyUCvw2EvGuXmpnxg9rFtfgtkaJFNcinQiHUB60x7BSAvk8FBXPOwA16gy5mtly2tSWjaG1pj1q9
NcCX08QFdTKfbD86v/yAUVI6eLbAjN7A8oQwCikbfETBu3BWeTg3Azc+PNQsJ9nDugAdH1njmu8n
skAEk5q4XLrGIB9uw7pC+pSH8FYlEDG2Bxpg2lXZPo/kkN3LSOuLZANRKqMgES3EJd8CZ9nYO5lZ
cQ76QZ26a037TGDZi4np0sAzaXNbcBoP0+tSQBWVTd1O2O0ltrVmUWQQ2APBawAIlSqgDe2ySdQs
jhsM/YTTgZH6qXdxeppUKsyZcvvCfEopMa+IRVA+zBvDhIV1/V0Zwd0m0RJLcI5oJIjfmBE8+YDz
mRkB7m0NDDxizccwo2nchhpWOcSMmI1/L3FYx79/ReTOJS8/xav/fUYVR/W5ooKP89SDcjUs3raq
BFf8pGcJmqU5dDMSQL1EK65uiG31LeBPzGLr/8Yg4WzEeGO+F8PY2Tq56KqSn7yAnNg2f0MuX2Ux
jf2Vz9+N6vdp5H5ivUgYV89BA2RC6cHC2uSHDAUm3EMBHHuqfGFIb0SLVBxa8b1Xs1QmqkF5ydBb
/lPNEH4Ozx6e81zYY8NByHtJ0WM6hRUspq9tRDjaeuiY/R5oIvfnLoCfdB48NV7lz1KPhyN7vtSb
jA6FBJYHCle+SobBux7ivNBZzneoX9af+HPhTL3U7r01lj0O0Ba0J3TBEgvVm+EvAln3B/9CsY6V
4SnG7Z5xhGaXYAgP5SERrAmTnPiwGNyR8GBusCJ9J+ngs7Ij6R87V9/aymUWNaJM52PbstN/F/eZ
PNgZ/vQ623aZea4Cui7zSr/E6PxGMefSVW1PCywDC9zCmSni1UIRfpw1MJ/vwziZJ4wrA8kHFZVO
/aljqHTR6d97LC4CLJ6lkPQ774CUEQcKtpILo6I9ywXFkU/Qp7pT9VDPhbJNS3ABwVN4SCtb+4it
IJ36fDu+4Si4kThS87aXAlKpQeGzhQ4apkEgk+YGd7SaLqMh9LKmLGAwckJ3KKTWjGJ+9zRUVI8H
4CyGNPyv5fpLAoUs3ZyWZ4akfO2c95DTk0DELAiqaR0hchv94uwOBl1bx+f9tCbQ6k5esLvWqXpV
7/BYflv2EVWS9BMcPzWwQlubOFrMc0xaHFhUyGIpuhDvX+v9KsGpVKTR2M1yAFmXpvilp60K57Id
7yL2mwmdmu/1D233o3MzC3LLvgtjEZp+gO02+AMUQDiBry9zznKVI0Nk+gH4Bke2vXmfmkNeENfO
Yc+BlnHeVMVpFlOxT1b5MG04x3yiJoMRBAtNTO3t5QsW9VK4wTNbHeePfibFPeSDC/Bl7i+Z9Bsz
fQ8i3oDCOXcPbyJs9rVlVBvnVzIGdII7WaSDwW1CencImg/o6SQFMGBDeXpilmAQY4vDSraBX3d6
pr14c63dUgRZ1MW6DLLLxXVf5RUT3s2WLFH0KML1kjLEuW+2noAo+8AuW3HmEtuwnaX+lDmvcf76
nrMQRJSQCiVKFu56IhUVk5VGq8GxTYQzjAxzizPe0WmuET3AhgM9hbV/ChGp3lpiMvqGl7f6TQbN
7aM5RlADno9rEfH/GMsPHTKBd9iUvA/FX+qM2Zus9if8CVoFvphjH7+5MC78aBbV/oPxiiH417eE
yMtZyWGtxV1nvsb5V2FabIBNhpme/gHr5FPLNLzZ6ouMhrRIjzlT2A0MfZOVaLpo4umBy3aeaY9N
Es/d3k7OY2Kh8B4pY+53DK83C9P8NQr0SmwxSnpRAxIURau99kbo3/pOEQqtUC5A4vGcWEh8dEge
46uJQRAtNYEXjFTtpwXE6hbIT5Ou34BnR8nNZ+npDwdHMKLgehAqZVTo8NAWSrdTy0s/P75n4+fk
JHaihnwm0l5DkJaE0IpoZsGy9j6wKyqyAZ9fFcNd1Cja0WjJmrk7K332J1n10cr4G4e/ulbuGYiK
FTwWh1T5JH6UCYb4fUe3+pCrpQcxtgo4dxS9CDSa+g9D/hA3atZobWRNzME6raxYSYGwQ4TtzFkD
aa9i9fI1gk2fXKNqs5bGhACf1od9N/qqpvkLIJ5yorLjD91y3b/VJLoZTipBkDBXXWGQoKrxsaQ7
S4xvwJnM/VMXEcBOR51ASidvFiLb0xhKbdYGwyIfPL6I8v5j4O2M0qRMjj3sblE7dPLIMYKuDc27
oTZPRBev9eDLuZFxatn6IP+b8LJ+3/PUf6fF9mcp4eIB4Rx8K6DI8tfN5HQzc3BciE7YcQs0KXnp
RVpiX/eB/0FparKXmxdk/8TbsVbRVoq5GubhH7XXaEs+OhvOAxSeaXmfiYPuy2WLetWGO6zP6WMJ
zQ/MslIWic1rvk1bfMERtQ4gRApmTfKl6CCSMb2LlF37tM3Py1Ye0kU1+138aixrgzR+/qk6U3J0
FvorXfeMssuYd7CxIwd4xlvR2EUXYz64gALpdAIprDjRt1jPkSiFPaesJ0fmJ5JJbo3oUrxSkbJ9
e9a2M9RCc2eCJU5SdZOrBjvxEhJIJ553LFwQQ7SOMaBpM2H4l88Y88Wdq8DbqY2bCBHDj2INATVv
DAjX4UbYYNkOUkgF5k3fhLjf/34J/yygwHrvoaMSMqVLoWvFHrpIsEXUjWizpWZ43u/TcJ7V7nfd
XqIMW57GWrUDGXtlAAVdpGsm64lCQ/BiJGlSzTJlvbCE3tR6wjqG8Dl5EX9u3yMOIgNaxrIXMjj3
Mv3mU8tgDSp1N8r1L6rwSdZc25O614giFxAlGN3bqULq5Tsko67MPvs7zw0Kugd2fheIMHegI/sj
RnPKKB9bqqALvqgTZqOhYwJBYuKbQqB+yZele33EGkFpkA+lynJcgVH0abuxVZwazGv8PHOeDWLg
ziPFGoTqtMsdxOSBgDos9Ecn04csEKmZ4/AumyPt+qptS5JekHh4gHplP2eKoWu5QNvyJm3hFc4P
56K+clS8LsBmmblIqcLG4dNqfTnQlu4iSwxa75q370oavQEpXMdLuJ9zTJkQQL0V1uwlb6j1KWRF
oVGldBMw+FI7BTQzsitcCnlCZ+pGU/YwYEiTg88eK8TRDgW7/FgfHUl0XOui7sWA/iZ5Lye8GsrB
KdhhMk95lac1GHs2VxyNTbt83LrgRKCJEZ+/nc/BSeAomULksbIFH1bSA50mE3czqlb7+K05E6jv
KrWoCnASxJX4bmB1d3nRFjP0yPCyJyCUA8l2nnreSXC/SBAC9idPP81DyCscE75bol1D4dJ+jBdC
VqAjNAVuye6hFK3HPgmNxQ2MICTOIXcspccQFbAOjH5b/R8NEFb+svPAACgrbUax26PANQsCLCsu
jreFqugk+8XERdO8K4MOvKcxPM9beAmFEftoYuqjqMdVPZJU+MIaQSrtEvbQehEqCLHrMgJUGco9
GT22z8GDYAtoJJVDJvXfzH89u2DKHKrDN+BHfwbwYYRilJSE2wriU+P1qvUPlph/uV2c/S4X3BVe
mfnmxF+0s2MMjjraY1bJIriCSwXVoSgYTog8fcI6F96tqCgazp8vGSexy0jhvCBCrPj6bHZM1ZXP
ZVVnFbW8HXdP2mKBDwA+YvMJrmieiRqzytKlRpLGbLvVFfg9TXODApjyyytv89WV0jOOpJf798Ry
FnY7tgAwaY8cfsiM0ayEVdWC8x/VQ84z35yr/ptkF1pshteNv4rp6yw4TX7B/8F6dKpSwEAWwGor
Ee/YcmVABCk3NATOid4TC2gBjO5oCPopqSS4stIhSBxwAWrDjTIZbg361yzA0RUhqg76Kye7Qz0m
u+nTGjXnsiacd5Rz8bLzsWbpsUjU0pGvFk0AwxS2pjjRA5ccNnWNBgKoixBo13UkQQfnMJAmlVdP
7OoCFiFKyoHGPa9SsaMJwOyJNzLG59Y3mZW0EhNtBwSvtHYml6xzGapyKCFogUBY7ao4ehirX6Uh
f4LxiUBkDZA/wQkC6o2LaaVhGXYAsFVuBOib3TCnqS09i+8OsQO7XWdE0yt6YBN3YQJYrgI35KdH
FiNEMs0nSjr9A4V0pHufPI1wv+hyAQkgKoOtntpS+AixK9P4tJfu+IyVVe59QGHZTae6wz7WN8gI
ZV9q4z5eHpgHx/pIKku3RjKABxtjkIBu+lLFELUhPdhShZf1XQ8V/VxITMCADsaDbt1wY30fGH6P
o5gdjZv49hOmobgD2DReH4tISKtijEN5BVXSbaI5O5WXciwDC3Ub+sXG+6Va28a6fXg0LkoVjIBA
Kwlm/YVarZK74e82UK3lkkP782gSIsZOnOQaNdZ/zZBCh1yxaBVpAeHGocA6GuVXrBSv7gWn31sa
xYnYDvCkPl4i7ZWZKH7lppT8msGxoWNFukpN+Tw+l0tubDK1JcBwdobiriuwAK7klR1pd0FISy7R
qs/ZYX/gIGg4oWGG6S7bt/9Fv1d9ExiUxIclQR7wTYi0E3ukBr+x4niqWMReaiVvZ/YopL3oEyOC
wKCK5zo2lpivxK4fNOYO2K/bSLR4JXEWEEW4SZkMnCvPCvMCir1gtnu2kwih6j0jRVpNoQA55Qur
H274CrMTNuO5mC75W65hW7M2lcwKIJLwNIsRo/UrpQKCELn0F+g+hdN8wDoBkW4JDHuDoVUzNBqU
klcKju7obxVBsZ0HmCn2VOudMDJVeHt/AZfIlJKK4u+dRj1ly9LXumYpxTKeqgtHm+9cXbxK9cH0
lOo0Zhl3kSxFHcNOVQPdVuec1DMTCpbVDkhTxCudtSsisLM62pGSDb7Hn3jI3GyS8P6scbIgXZSG
5IAD2toITBZaBWddV0jTvtEx+gCA0ru5o3UKV+srjfNAp6CLjG8VVrDH4tHKceN2WTUrF3A31uRw
jkQbbJyrmGL4hY0JPObPRn+lHmddZZ/xPFpRyRx1T4LtOgXPhU6OZRyDGHukaKyc8D2O47jpSjwd
S+TuKDQAURmMm3+ngeYr5dvFDwn4of0YvJYmWyWJCc1GRM1XFtXbBmUXBn11UdOc4rvbCgWwEdpA
7myMqMbJEbYLn5qKXFnoHND+K42kwjlkbmtqiaP9wS4hDTC9y9wM0WuO7OqMZv7ezs++lJbpktEF
9kJ5rBQiPqzIt2piJpfhF7P/LUq91DOO7u2t7qUaj/QhWmpf6gT15DIbsbwRCRsqlAG6jNt+XB5A
e1IHKXgyRmNJQnvWiBwbhZ3J6cIx9bMYf6xyXy6jBaKKro8XYwhFv7wRAa6zulGXnUac74K5DMfv
n+YSsTrJcuKWARrPJa3F1ojwyrXkiJ0E1twXCCPPI0hFz0Gak0sYNIbRz7StCaDn1VTqPdlSzakJ
VYzrmvXlfEYhHkZ/PyqIwg4K9pNHFuyVOUbvIuaZMKWRCmXZTmRA5UkfYLrKDUzDGqbBVFA3wbLq
lwcpihX+gTkVg/QyFuQD743wwd/oz019jn2vtQppO/ZovLDE0ojPuv3VPxpHchKE/R4XmZbDHUfv
Hx3oZSwSo9ekqapZi0MR40ttkBrOgeEUoNlBfJMd0gDXENb1HHEA/YxZOGkl7Wj8nWR7LNSlfIH9
PZBMZCfLA7m06f+P21oeUnjn9IcPhg/zkQ2hjISLdcFqaIE6Z07IQP+IO7MQaxuK/ykEuD06P0E0
HvYk0pQBJsJjzzXbpqmGm4cMZhtKsDyrZxaxlte6kxf3VpNfXTbA60/mT+gSilCdE2NFEMR6miWn
LbLxy/71drddSPN67M+7KdEyyTkfklZmGQ+o3Bz3XIBMDUTE74MIFzZt1rgEUJWSsXIDxruJOpE+
LDivllGsMgNQ5CZ/Rk7h+oC/WaVTNb3CDvOaV2ugkg7Y+BZv7RQ7Vihr132/NfbOC/pn10H7CCvI
CNdVI9EBx6vuntT+EsFhMfbZYYoT/NekdLZ6SA6UDimv3ACv+pgbj65/tMIvbJgGosHaSnrRtLzN
utlSDUaDurBAsWbGpvR81PCgARF/JXaElKlcQH0weH4q1xkCLbxFKu2qyY8r5Zlgc7ARsj3WkURK
dwW3G+XSKZxGhJOSdIrj9/wkOGY+ZKtpOXcbv2KBCPfLZfNfZNKR9X+QZImBfIb+O8muI3DuQi/l
Zsa4uJQtGWj5ubUlO3Mf6QKxvAyurO0a8J/VZE/cWJ2ZLfvjAfm4v9/9EtcppT7cI6zNUkpk7KvE
hoFVY7lVBzSCc5S/cGbPqU9n4ZiwPQG4mtzZ/dRHmHeO63qrqUulaolp+dczF7dEW29vGv/Kn1n6
Fxaz9w9442Ygu5I71+MxNQwsLMxs78EB5bh8adKobyOc8TYi76vn0OC77cOI4NqKpgHYMjfMVvwO
lXI5ErsYSrXfnGaV53g5ed+9dpQkO6UbeBgj676FpU4t6h18TySOloRCQ/SGNz42ceCJXRfdjapn
ugzADTDg1VXzZUEQssPSP/pmeAdaQmCRNR4DeH72A1ufKOt8xxryE+WnwF3oz13bzHMlMGr+hYTZ
9WuSMBKiihm/bt3St/YO8zKQ2EZw1HGR2IEJN+plwFWtsUqFP3KVm0MmHLTMNIMN0xF/D+1itoph
kYgewV6mq8J6OBpiNbG9beBnJqdXAxZGBsbU/iNVveio2PvAFAEcuzFh/7s7/+9s/ruxfEERvMqw
a4oq56oRpoiYH2fkybHi3jrnexyBncUoE5saSn+rC3J4X2Qn4FY1gQADadcs3QuRwtfFBCBCD0p5
nNf4YbuHZvNqZDIAVzqbf2lQ8gQKaFnpkoo8pb/ajvckqjIb7tTDKLtrosjJNyrg35Vl+c2vJttV
0pa1g1lUODKO7uqhHFBt/yyL8kGFL1UHoD6wdwovdeDtIjDlirAW25GBxbJ1wGO78GLNGbajsxKT
TNNNvEqfu8L/G/ltIS9dg8l/PqUkhvCF6SFtS1HVDo35eniNJWDn29BOhNeW65IIZXjYETtSix6E
/MXT+1iyS5jATxYxLZeYl6Br+U8ZPLSTi6aVXdE6lHkWjt5Px5mz85KmMJL+Y2RYcridHazGrYO6
5QXy7y31NesPS/N4zbn0r/W/R87PuALfU+I/uz0bhW2s7d018AiE4n5vt/x7JpXaUhGn0JQzikdx
GQF6yCEoKR1SiWhGh/G/NHDydrxVGvWtF/4M6v8EI8RvXmmhtyEQhUph+jWpmNIHv5drVrD6vHHb
ypQHYuqko5Cj3AfZLWpNL421rjCmrzY6NOKDSm0S3y0XzNJncejNoFNF34Bis899G/pBauR8DUpm
CwFemEPpaJNt21g8037pE+nlDdn2f72+S0RDy+9tG3XwIGSbzWeKlKlPNzkWHHc3A2Ta3KYdQRpJ
DLS0MXO8k9NgJnQdubVd3Lm+2ZDIdWHzILdSrOjDDeJyAmH6iXKog9QFyDctnWPnpS4emJBJ6sJg
e4TtV9mUmN+HJT0I+5RN/Jc3SkTSndajXyaJDbc81zIevBtjhZ3XPSLWxdR3MNIGDW69Q1kxHsRj
SeZPH/Vk37Ld7G9iDgWKPapxgxp4GQM6el8eWNhEMqfWhR3jOghAIfce/ZYNRgTPNqUONPexUDgv
h1hk/Un0TuSpm1kEF3RVOo3GuglkWP0obWH0/DdewMdidUyy68EPgIuajJ/ntIOm2xuSe5WiIcBl
d91yrgu60xG7L8DPYfxv5pKty+5N9yEsEFgWl3+90S+/Er1Vo7kFlcmPmsvC8FBUvSLZugCkBpHA
84jhBzbzQBxGuzNQJWmzaAWyFiwZ12TEuc7ow4+28RiMSr+nA8bRxKmPW8CYGVdji+ke0mpqPwS8
2jsXTvMOljTLuFQKpRmtAWkT4xkOxYbe2z1RNaMEs4RZZJAyS67tZW/BJ9OimbeoC0+v/l/B7AwP
33FyMxYqLTqC73frG6iGBwcjvHGPf1uRuI1updUnocf7ML32hL+0K+9bB2Blo959Scx/kUzIHOax
1cZT9DIty3G1fugFCDbEJ4dvcL7oWCaFnQh3NRQebzrQh0Ccl5rGLzLlrNybpBzBCnIJW58YE/a9
WJcPhCvKj0aR0VGFxa0P4FZICEf9Iab1ARP0//PZFeEZA0sNm93x3M6IUFeQNAJ4O+U/LdLhqauC
bm6FYEjQlyVy2/FOeusdHh5fZnmnj53+7tGxq7VupcXwlB7Xtns0CHqBea6RQaq6X8cLHS067zrT
zQe5uGbPIZqAfzp3dRbcpl8sCCl9pXlnzMJj8vIR5QYJ+4NsoN+moauIfwg9KUI/vV8LB6o4nwLz
d3MSZHVn0Ws9LDzUks4/WV47vmR2EGT84wPp3CiY9zgvhkolWdO9u3mvr+ZNkRnGF/KFOeQ0nut/
JsnaT74Bep92GzURqsqad/sSqx28/drdiH6eSuPAtrsZhQK+ki5GDe6ac/PPYlwf80zNIaFtBOCf
PGArPyKQ7mHRG/RMjxfn1+Ak5a53cTWFwijVDjPcNlFVPVu6/6tGrkCJdpu4XHZZI+4VtYn0zTD4
zpRIf5FEW8ZRZ6SwfoWXsTBMUZmeLgixTP0srN254RZT7iH12lYgTskQ7PpXHpL+IITWDzkNf8WW
9XlqFHzMLBpWS7t0Ekb5GDaeKoH9vAdMOoYFKEQEQ8UIDHHoqpmtBXLGPkdx/9w5JH+401c3yznF
3uFCxHEZ+NbCiT5QGQa4J/p65mqxwGcZ/SnBGUGJqikaKTvhi9qV8LiVA+aMTDWPq+jSHZqxWgbP
Rcy0nGmMGRsVNIp3hTga4qC2G1PXpCuiIHAhcQr2Jdlb1OND9kH6rjhLljfnC9B7YcOlbxuLsNOL
nxGavwJSK28Fj+hwsAJ+pJXVitpZcclNc5YARcHy2FaQu+La1eMPa13LwAByC+InPG9P6EUIvokH
NNLhx2W0RZgY3lwuI/il3GEaw9J0OIWirCpZqYaW53qvgk/EcPYb+lkIQgS8H/s1u16/S9yYgsmy
SFTw0MrxdGJ7husjKFL4Oys2y5zcYTRyrk2UnflBpDhkJZv9yPUWmduT/zZ3horCwQaaDaRgJa5W
+zxvEf9IyUo60Vdr/H3J/OwaYGrHldzql2I9/xndLZBHSSH4p+g8nri/XjbrP30pQIkBdqSjlg6q
IPJrQ+OiHTsU0KRz2J0hGRsFLgsxLygpAnqHP8u+ToNgvtB+/7EJv14WoeLrYp2gz1aI1Q3R1vAr
ehcB67KVPF+UELz2noWxHBPFIz25pADiUJNPbfPF0d+qEV1/qFvGgMKvN+MM/aWHEHe7VNaQpA31
UTD4xocP44OXpIINnwAMnVZ+8rucqpWlRtUGuAm6Sn5QeVb0B/l2VfPjsxoGVjsX0/f9RX1BBx71
gehZYVgY24v+z7X3E+uW91qdSxCZQTMh56XQ/EQuga22cD+JXuGPtSptSOgqFKHQppgRV5i1aZg4
MuBWw6YXgSJCZU73JBKmRAwCoV81Ijup+smNxosw8IenMdMyVHsL1wfv5KMTBYFKtLu4myCJx2CC
1Iw7hbM8ycBIDPQlbhdtJMT2310tlEgvQgAuNNEXwkMaOGCDsu7dvueCOQi7drV5/lJL/2vPuL54
69NSjVArFXsS6Ugs8BtsJ4UyLr7zDFYA2MUrHVA6W1Nfr9fhXGIJ1NxwiMmZsmblx4y8aZVB9J9g
jCLEPPyLuCmaRhCZQiCPeKG74XwoStvqaOMdflQl6DY3Uv+nl8Slh8gxkZMjMSA3jfyxvv3rWgG6
VixCsKHg8+W/hDx3vN2vxK1805S8bXEaJ6wTl4VdraZv4SsHq9ednFN3Nni98g76q38N4ZseowSf
FWI73tjrOxowSVJOnUJixu0RcBCX875+Xt8ycFOsP9vAJ8XOtdIJDvlRkrPo524DmOWxSokq9jFi
3yrlD8kr5KXlJSnRQ3BHWst5c95dnbPOec2ltMraTnCQkjzXCYsr7/pC3+c4P3MA/VAjJRBUBzfg
8iE1uG/BwksoDzdkR30vsXSm3gZVURHAs07Xs3KKP+u02GjdPyM5BXnJ8ww5kW3LLeOjC+3Wl9cL
xMuFVi0SMSDxY1AM0/b6osfsmDFLPbE/ohJWyonb5n8WyrwfCRQCNhsgDQYe+N4pXjS0Dipa69Yn
rV5Zb0OVu0pM0Xr3o3fiCbNTywrfLcIb6b/ylWjDTFOXhru2CdjLDoaIOK4hlU0ERLAHdDsR6sYi
AK+/+Sa/YRALSnFLdH3SWSKq+OwAnJUXKHZuDGlbpq12FpnRZQvwP3UDL1JQMwHIKaV3vfAhJ2bI
v9Pe33A8RlxD4FCus7c5xUvrLEMqqw1IBsSV8tsDBz+W7zlCgeqDk8Ypy1FxFxF+e7RLi1Qzx6Tv
TqnyuLcWEFZq8VOk6cEjfTxiHzSsHpTOezkBjHFtJtOS/GCaWej/ryGzBbbiZxX2oT3UGlZV6B/1
aeKvyygz8GHnPVt6mQ+yMtSHLJAcaz/9P/zTVU0WW+o0wUie+MtYNQLuQkDHpF9DyQ7pDiiLbKDw
tgNe945CYaGTOZmBllCApbaMU171xGbWEMOC6RJ5zHDLvpUBctPo09vm0w/CZEt4xKMbs0WanrIj
YL5kkQCxnf/RFrayBX3hWbM2ht4+2n5n9FHEAf/FGh7XuRZtsD68DBfuM4wRkbRw0Gg+Kpzm5ffW
ZooRuvnS7FqsRmWh7tOs4Q0/VU6TtClNAX1neDI5laOuQ1ESUBJu17vPOhozR2FicRZJAOpSB5bU
qIaRg5WYbjyguy3/WZwGM+Q8HXK2Oxxdo8WCwNserJcDxvtQDP9M4sB822japiyKTEYrx11FtIpW
PhnINon8Y/5SYcF3SELXL+sh0kB/zSuNVLPSKPBP1PfoT+0xxCkB6JO58W3yMxzUtnigeCkhK5Hz
dHhaq+zLkkAq+8UAFnuOljo6DMb7CxV8YhY4akIEISvAD/LJ2NY6yJ0iF7CzIUkmMwUMUqTrsfcy
XnAdylOGz5LRjNmWQ56xK6LTJLnFqd32Q4Fg+dfR/0YBUVnrQBnk0WmD/Mqy6Xy9DkFqF0GXyU/6
z9b/NWSkTwByCNGvTVaONcLmvrmUOz9UJT3AS5Gg5tpsJp6NEmDA68hqaOSnj6JQ9bt6fecew8dO
9C6jg/qFmrNYn22kcJEzXy4/d1SmWWCStWf2HP0KWbCX8+nWvLek0+Wn49u9P97ySiLDI73+LNy1
Vg0gvyR3+N0R1PFq8AvinPUfgh+mMCXk1PD7Jbp+KyaUod/mwVt4cL0rySsl7C2BvsMEiNqkAjyE
cMJmLPNGwph3Xa1/hs/3NkS9IuWMCeUZfV5wtpcwsCe2ty42RrZ3xlk4DxhnU+UpGUbBiPTP6q+Q
8FUQVuhKkBpPs4f9trhtmh8OsP1uRiOLpQ30QnfufD+qwLornK7AIUQzUH8noPf8vGeF8tWCLSzF
6tTkw869tZ62awm1owWzcX9YsKPm70oWacBkkkv02ULB0vbglbkT97wDAL6D0DEhZHFEebmeb2dj
ebDYofFbOTESdGwrCLD5tcN2GSLUGRszvNvyQ/dVyOwV6aPGGsXmaIuu/HS8Y4kk651C9xHbhYAB
xCa2RXb5lyZ1Jy7245jvpeOT/7tRFO3YUjLi21wQMGO6FaWYUHtLJJfdtCEz2LuHIi/ZdVWN+777
P7QHzjTwQ8CqEyZ3EcLs6zvtuGQVkdE7RDN7EZXqbNRJQ3uAzjUVjT/emZh24ZdwSvurwekPRKvK
zdpDHhqIEtdF1axmSd9f64HKpfN3Fgvj4VcE20b8fSDXED0RbkGwI42/6B72/3BWXJfjGGrTYaNB
S3ExfBnOLd7XoJb4k2XwC3CrEeeXtOkkRZE7mYos2h3KcTeCT/OF8FAT9TbyNr6PX7JUXFn3IO5Z
uaemh4UhxV4O4z8GRUFnHTC2I4z2hyFfuZ7tX9iJ13nc6ux1vdB+DH7O064ApbjFXrmxnW7IdGBX
QYgYSrdUkpi4jUZ061jEew0hxQ0izhKkqKH/t0pCMW8gP0SlaO+rEIblewZZoOWzEawgGyfoFVDw
wIuziwxI3a8k9xSJsSrpG2D/FHsFacRj4n/7XyfMzZpIUOX4vxzht4CSNhZ3LiW6IC0c3UNSkdSI
/dazh2z8XqigA16iBYxZfV6xJnmyJDSGtSDMRbO/4YhqHd9W2Ss94LyC8Or3EDO34xtYVIN7fqlS
QvGmOTLiKOTnzW15VbTmztf9IeQKzD4XKrrIf3kvSiLNcVGBogAtlVJf2aLyQZjWqQg4LgCMh/KH
jOg8qCtQsY6AJrNVjTZedY+wqR3IWkT1UUe0Eq2K6XbP+JuzMxHRG5wG/1mm7DtBN2FVPcHHLX0P
qKoWws60jXFG1oTgecPjfVZhJ18NZ3FFkd2TwJqpeRiTpqCmc1pxPoKc9p0H0Aj9axMIh1pP/UWe
RrZtFDC5ZVHHe0PSl6LS5ESJntege8vWiTlGs5Y/SfaF/ntqe3aRxk1gO/j+TlDWFUysRiwGgE+8
chKxRPHR1eMs+9rlEa8aXVeyE89ZStya9TzgY0VDdbWYPVh0tgDbq8Gk9zO7ruegjzcHR1+jI8TG
jT/lnQsbx6m5s7jdku3kAD8aD3cVvPSr4l1Fd1aExvZHThNT56IJvwY07E9e0QqjVnLrTGgQuef7
6sxxbdEDboCxeASMsrRlTfZAHRRd+P9/tGgWwP8vDTAaZS/LqAHU/vbGBD0z+IxQQANkI9YNtIuo
dcuucuV/RzCsxvgxFrDs6pdQZ2SgnOIqHsdsDlOhUFIYrPkhZXcx0aTnzsLg9WminYARxi/hhEve
doO9zTYINQBs/NyX639HgL5X56vAVgff8JqWcbseqt99rufE0zDJVnPwd3o2qqAyifsXoi0mCrFF
X9ogBzXW22Kond6pokmrgZFxy2pmSTUqINthRfMzGObXS6Ze165eLPt9ehdCjALWG3NwzqjoCWz2
ZWXQtCBa2enofnuUN+BKW8w/cyaW9H5I3Ar66pAEM/zOpxVkmkwBJF+FL8U+tmb5MGbif2tXbb4v
rEIVU2nC8XSl4YyQYpt/XKJr+9dQven22MYTfrU7pAox75GxS1AaHEerZJBbuHJLPWfs1qm4TeyR
+XEk0zYkmIrPWppHf0oJe3yLQKt/nVNClOUbAzp5cPJ9buPIr6T6UsTDht6uITGOGbClQN8CLMd3
ozRBm4mp2+JUb+fNGFpxNWp1w+YWe0Bnkojeiq2LcoCvy399oWAwspaJpDk5NBo/7LtdXWNAha9S
jF/Vobjs47yC4mQt0kOY+gK+waV7ofPHy34jki9yzaKE0xIgszuNPmIqMccGWX7Q5fDPoWYuwFkh
8y7b+7zL/ilPs2SosyaTjuR3GqwvhEBS9WBpqyZ9f7KooBVnFswT4Trt9yjefKzWIvaNMaSvkSAw
PEm08bsksV5J2CscYPAk9rTpVcdIrSLfMSsywKYKXagxVaUnnWXf+BXqFqqpDcJysXQYLDqFbcFo
lDXYYdqYYW/mYX10fo5ErQNNf/1qOUkMuQ7yOfltkjF+rFJ9I2KUhkbV88dzCEyWjwPFHOcB0X+2
I6N6spte3x8VYTZWvLAIpwEtf+FCYO+CVZ/bmyF5RxuA+nv/01y2o3kyOQ7bECIRNdc8kxWwcBFR
ZnmTSsg2qt2do/n2gBJtqBh0GufrCo/gfOvsltX+SzH3/7G75tVRoTUsJql4M+K/TMzlqDbYz52i
qieLqVAuzteaix4uH3glj6pZh4tWhjl2167NWFlT3Xx2Jy6+uuD8o40rRFDIuZaFBqcAvc8X2NHu
iz/kF2b7nYrsuDgNahzrKS7Na1zFwZJFCrojOJHyw3eszJLZU/WyS3HYQV9e8iS2lt1ZI6vYHoWG
TVT/ADt+sAbcKKQagFrIl8223S+Igjgzy0WscmTGqjfR7NXHOzSolDp5B6hMGd9yXm5enHsvJhCU
WXqPmG3MXcrjb9tFXhV20rzkTQX8MDVld6g0R3VKXRwNLzZlquQAB/0PoBJ4vmHjAFEPMjE3cQSk
vWIjWM8R0KH6zrhVj1mYq9Xu8GYCbpdf5/JEwYZfDLmUfaOO87+ePED0Z0fGEabxxcwEGIoWglSn
1+TYk5y2nztwVJY+A5gA+4cqxmltFF4O1VfYhEYZx524Dn3v+ZcbT8p/ZRzaJEIHkJMBHdC73K9e
Fz53bs8WjPTU8tEh6AlyHxkIl2BOkny2GUtfI1bmC7sWitW02ynrKaGy1ethfsKhv0EqMsp9CK9W
RjZTMMWzw7oygY6yUKNWy1DiSl6ioYp6OEcqgsrQr2w04FcQjTnmNNlE0W6J6nPJoEXLcJCyVoAg
ZnpbYwhqXS7S2KvM7T49wYRVsW1Eo9hVRSOTeAxaCqeTUaR2fdJv/NzbcvokD7Qi/q/vDTixzSso
E4Ugs8a0Qv+bDs121zPLKn+qI52xz31S71iKYynYZfAvOnekMLlF43sIWD0fdiZeFB2u+X8jR5//
CjTzWzg4Urs4sKAokWEZXRWzpDClU9WTyshdF/M5Z5gyxtqTqTX7yqDexkkKpnWy/IcWCoHSEtUM
0M4Yl1OGYj3MYfv5vTvCdFm1/YAhTVfh7gtTDCfGnmdZtwC/ffShX9cMM7JmDv4qrXeB2GI4xzvn
PsAw+z+A5v5o+H725IyC8bDtYLCYxFQzDVmgvvk2E9DpO79XbA0r0VsFOuJphCRh8EeIWV0uAOwN
cB70jfyGUgPwsnfzhPByuBZOD0UQso+Rw+emmDpbrYOBs48kaE5hbzilqtOkAI/hAcZCc0eJrNXJ
4DcPbdIouph8jYecG/A/vKYj/ZLmEedMA4R8+DHhwHUWS7kVw7GZcPa12FjvW2puHc0Dz4OqOS1q
a6sjHT0KJZWjpx5KMi+q46HLX7n7B92fBnJnyz+XqIkBF/8zoXKLYBBnMA7LKqn6B4h7DOyuIQQk
BQVD68snfHHUSALtk/jPHBfDTwTHE+8WLFABLxBZS0GzlRqkwdlr5Fo1bUfflpHlUJDf77BU1e8n
bnUGqfFvubzP+IQ6rqss0gkuaJYeLmZoub6rGO+evVW1vA6g4x0QQ4jgj0+jiMjK/v4xiO+fcV56
HNsIP7I/+vLmavX/IET8Gbhnqtr4VV+dBPJ9TA5rwdgYKmbJwWHyFBcQB7ncSBdWFLOZn4evDhnH
iWoI93+pAQ6h9bShnwcC1pe5rSJiwLLcOXMhI2cjs7dulNpO3y4iEsZy3MXKgNzC4BkKZYn7MIjk
ZxaUnQHm5KWQCN0GvT4Vo9DPi4L7Xv9K6tcJS6ykHImEpz1pH3Mg5CicBAH3uRJV+ioFEnSh2UbM
E6detmevdBMyOxuBJqJgHKncNAAeWfteaNCTksOs3jkzUGhzSIUPCQQJaeizZJ7Z7h4mVpXQwMei
jy+tA8/UBw6AShooIdV5yv6MNqVy+3is3qur1JQk7g+MPL7jZFQJpwY+FGx5CYOPmff7zIaKimy5
inyvllPamVlwS4ka8sllE+H0a6jhpFS0eR68wWVCZ51JWI7/2PAcmYZLulVMjb42tm55VGL6IhpP
zTusvKF0DAKvdLbtufMRbK+Hp0rlpswL68C22+wqlwcuBzFNPu2NA8yXUyzOFIUSrNsCx/QDLW+L
Awf33TMIvIWSqzDgav1pE5s1uXNonVGacfc0yEleeDzZQIFaThRRt0UQUo10N4FhNW1AkiMZd7vD
/eYcA+pZL/OBIuOjOQwtKsVzmtE/Nnk0oziz/Lx76F7UrlIBkowCYRtsWohSZU/BktRU/RxY9yuR
tTS7S8iYFlbrcihCa/4ZgYQCiLn8yJWHDMJ5C0p5hXyq+B1P3QjRESX+uYqabxvWnqFFAEqirb/J
+BbvRxo1Wwoir9j/ENWSAni4LIVayRWxdUdicKjBAHyqJD+EWaAqrWkUnX/kyipu5Hj/fwR/8OzJ
zeboVoAzHR+Yib1ezupINRREUmSNfAxyNrz2LlI1/FwhZfoudRcu3DNElM62nnwwB/umidOPLF2T
Rl7NZ9F4BxK6YGPch9LxTVxnGCzVrzueBaBPA/hwvB9HEyuKKkuQyO/wmTPtnqY4BknwkjWuuGk8
Sn5uYG6WrFAaT33SVwxsFMLCbrUWTbQZlLk0OkOe6S2Rf0IE1cw7Z/otstMPPGBSMQUYeKqRu2Ek
P7DM7UKicP5eviufKPR9eer14s50aXj1yZ58AUMbQYAlFV+t+meLgRhZOyhd6VeRf4+IwSCeKmIm
pukC6EmyUDyqlHthnSmPzQQw4ltG4ePD4a9tAyi2GiG/Rm1jRzPIcOsdrKJBi17pCCOjHAvwlKyj
GXCeOg0e2FBEN+wIVkOUCd1D5H9EUcMKqpyFkNfIhcxQF0akp0cbI4uxMXIb0S+BXuPDUjJMBh/F
yz3kTgDjfGahd4pus+YtT5qt+We8t3KryL+deK1Gu7F2tGvPRhT86VvPM9dkoHNa7NCPhk8EV5g0
+REWCwFsgfVNqOuCm8cEMzAR7b6LTDld/aHRo09ZhjdZ9P5lXQc+dXmeCsvFW/pLyvqf/adq07Xw
EkJ3Z2x3KVEknGPJDdjtiuJHfuPd+ywGRSv0UMkJi23PBtkviaXtNXKIhp8DchMxSG3Atcx47ObY
LzbYVRbnPV5w08ESlKlaPw2UceBXowvXfv7mXu2+KZvB7fSbRZf5q1aIPJQ2FEq6FmKARTMOnxNZ
aqaSFMhldCbOmZZK0PLBwbhV6Hlv1YfcJdtWjEfUY2ulOEYot4Cm4wCS+sSNxng4PxUdnN4C52pb
dpB06fBXJgvslsAQe0beUw2x76kGyX+DiZ+WfDNW86hu5z1o7GxhwKtt4uovnuLZDDWFy1rntq72
WCtVDRG9f7ykySUyAmFOaci+CWHTS+JDbYMgtqf8Yui01jhxiN8pyZ0cZkVLa3Sxmcm+hhIyuxv1
2vdtKUTU/sG0DzgVmiynZGVAEGw+t9+4UlDQikd6RsHedm4U/zP8v4LiHSfCN+/+4DKSte20YKMZ
HaIaOrB3BkM2/zzVxORebRpn9zV2n65tKdkdSLriEIIdH24tjqdiHnp9ut5g1TYDUjCcxxfCbSS/
XFfLQKOHMWBNTMqk81RRt7LkrRQKfBx008rOmzUbMpftvUUIYGJBv8VgALPCOabNWW5Haplo9LqQ
CvtwEvj24XKk/JH6N4ourBWXACqYnnnlXb9DWwFWgc+z1bnxzxl7LTIpaFH8X8NlU3DSBEpnDG+1
JUEPFAAT1tMUtCJr8ZqVfs3hw19BDPyCfrx9W7jz4XezgclH3LqUIJ2uJucL+qFutn/IBLcZ6DlN
FxeZwxzUSfnTpqumKhMZXDRZ9gDgI4l2AsrFfSr3uKtKe+EIvddNVplG9jdF2V/skrTkuPKnY2Bs
6tPW4PUYVSvzZPqGPZ0HrcxlJfH/51eDqFCEyS6DBKrlkNn2UOSGL81VCVeo37QBuAxktCr3O7Ra
JsxxsZjx6BjUprMwfdp8pkY2TGCwE0o3dIYzPrxVvKMXOElq+4qc2SzSiVZqDG+79ZGJi0poWkkz
e8fZmMwowy7/LmTAEqem9WeIM3WGJd9Y77wcq1FtV8jA6wMp8P57FkewUL0fG21X6iIcfhjg795Y
kAwYt2g7DNGb3opu2Y0tDEHXW9DU/askspupr+2VPZoQNdbeXuCiOQSOZrdM53lVz1gEL4FkzfgF
uzaMZ1M9AwfjX4VSL+YK+kHnOCm5n16Bg9qllLUc1KVX14xRdukMIXgQKmCvn3AAV3PLu3HMYFA4
Mf1t9UK9RN4/O60P81aUqUXEAslIUGsOoYYXPeDFD7A5spzvjmdrn8XSy9Exo/+bRCW+YpJOiHY1
o/GOKramI25KlI8y15T4cKQvRBk5nLDWI5yTRK5NnN7zjmZh51mJKsBqMHwy0aizMS57FPuy8J/b
IZHOu7tc9/Gho6WbTL/HSVe5u6T1HOeHqnziqUfiFcTNNSW3rHle0syf55F3Nk4RV4/SqJkGftrU
7g+09EAAlvCQkoj1VYmMn+Fe2o3zCwlLPil4K6iD3Jr2+GWy/qZNXVmzreCtXQLPQJPK3I9WHpKB
8d7hhllEWVQqtd9XyAHErVfXfbQiaIJJil8LNGr68lh7jWLYys2KHPQDlBCmC2D3EBIkjAFRr1NR
f7Le118J75x5jUYUpWkSaMNlA80NK1gX6qk72jnzGBK5hr4AiHX5B2RsMG8Hdc9Un28nekJBlFDK
ICwFE7bKlIClF86eoSsUSkythYpMzlca/GpLkD55VlxtR8jekjJ0SEb14r0cIU1R7TXtpULAbppC
qKEyWB3vzt4YkcMR2CZesJUBBEyOnFHAEgfyM/Z8KfElohznVe/+NQdIJJNodcf2wVqWDF/3CLbI
4xR5eSgLxSOgqrjgDof3L6ha3a8oYteixYuWJucmT8fJEg1fU10REmqwifA2lmfmDubYvXWqBgRg
BBNkWmoI7lfcEiSF+09SV7lrs3dnqD3xzEAi+T0rTX4W3BCxs4wG99QsXf/cIyyvk1jYwwXVhgIk
NqyH4hrylrx8fBkd5MDKdhpH9TZ8K/RqoYDrEWzoGPJG02PcUJ9tTtWn/LEh0BzaZ//KhqS44s87
z0VOwZ2c53kkte4fInQ1oL4grzs1bYfmvvFJlFXADP7wnxawL/i4caMhPomMahrlNy2+s9XxDmkX
LyB9ITCzpUQ7uu5vUgMHih4mwe5NogYk+fvEUKl6PrHbZWvYeib6Gx8lJZuz7QIRwcvQCXjgP1xu
BEv69NgyqcnzUxD/pREkvkyQcHKIvF5gtCY+1rCaZs6WQCOVDfvwXsWw07dn+3mV5/FstsmYbdoP
DxZizHJ0mG3OKkRcoUy55M9PZqGsTc6MxGoY91knPS9AQqvtO4KJefg6OzMoXSdbADp6JpvODpnl
oyuUinQfIDBGU2T4+SldHFCKZomP8RyKIp1VM49roxo81nXwo1UlqGO1s6R+zOvavd88yZPyRnqC
pBgEd3fBHtLfI7NbOQLvHpQBEPK0EfCivd83zsrTtwZo/mCEtZCnoqRJ6k0rXl88XTeaMy9EOg5n
/UrKOZKJIZABgIrIW+sS6OdJNG95reu5d32kXI9SsuN55Oq4Z8R3dK+jeX5LCMIgoT67CNoeDXz+
O2gis0bwAFB2AU57WCIEBrVpzOSyil72XWa6DzkQIPz4vZbSsRTEgHM9iUX3H2U++YtDwKgmltdS
FSYi6xuBB1AgQAMIBYylFyoxvAihdrMl5bdYvHMj6EbNtD0k1HHi6n+ii/DU0OABafwLI4evdQfW
Z0EsyEbBHdaDLGLpQMxUmOJ3wpfhO6ilHbOJnI8CThojKUB3pK08bGMbW1H+9JR9UX5uqCBq10Jo
Wj+QdqI3eZ35UMWZZ9LDGVaSUFF7BcGuaaJwJz5rmuUskZT7iv52OI+93N+3GcYbqxeSi1OxYUIP
nMx8mLXR7xjnv3fzWKmb6NqnYbgWa+knlRZjVihskyBWuz8PP6QR6nSXtY3o9TrS10U4yWiDOcRm
w7v6HqhbXS5JHwhecAf1sGya3zcT5LMzDILB8rcsEmaqcj+0qj1lHfBzGAhXt69LOEnMhowNk2l6
aGEpEvWCt84etYoQbKmJJjCExUG6odb5TzsC99MCxvIXHclanoSpNGo1C7fiZ0fRxRiZz/GA22Kl
fF7AX4YUH2/l4FH8r8drNRrcVhQB/aZedJHh+EpU4yiECDw1Gel9ZtRCQcJI+FCL4hcWtuv6OV8U
0mQwxdymQzuu3RdMBDUT+bTqotIDzHl8/OLeqbxhSdRqCUM7Toevd2n5T5If6M2aDApTFm3/2VqU
aTzxD2xXa42nQkkiHqqyGa+CVEAKznGPsGxjNWgtPEkx2qG6MvBORJyNtHAEuh8a7/Oc4tUu1QKX
UCIgyrO9mBErO6jQAv367SnIIE2paPO6Zv42kvMgOP401JNN7nSNkGaKv79jgJnIlpVYpUmTMAPC
QmHqsWcAxAbaufj7KeJ+1WDDOyT3mcKjbZjxbTCU8e7eMxAeqYZ621D7zMbjqSzeSn0OyqXTIdra
TunvsGpFTKPIaMmcDVjqT12CDVWpnBguKFwPyyZkYvfwwvOVcDw3+2Hxs6rQNhfS34boOA1EGzk4
CaSCyCIR7xkKXOmkcdMc4sQOgVzPYD1UG+tw1J0P/8W5bf4pygo45ZIZe1MPBgaN/a546NnQBehV
ZOIsylUvpn38GcSOz7qHh/6/uGei/Fu97J3USQ1+hT9DnX3Mg7kkmBo4u06oeFYAA4kN/YDax0XT
aPsTwm0B1RZjpcFlxla7sACbZrcTI5w7UJ6AigsTrcRFEsCg0AXwvzMqLe/AnDhSvx1OJGsHlMgW
uxh/6vhu/wiOOn0mgmiulMB7Q8TC4rOhTRhA+oHxV+hSCZ93zE2kAafa4leTAbemFQFygz7e8ZLu
vJX+KNyKCczFdUvk8OSP8yzEaW1xV6VAiqhAOBHbvSJ6kjSwiOMwXDZpqMC2H2NPBZOPrl81uhp2
nc4Id9hCx+wut3jCpMpGpF3/+Cj0TsxW+ImAkWprXwTorWuts6gODgjmrUbQyLUMh3UZKxwDTJmU
Cf0oGBJPuX/lU7VZT7wNGPNEJFKBzqCHVaEPFDwLetqYKBnPte2Na2j+QquI2sLgu3Z9zouvL5pi
jyJOQyo5wmboGf2leRecu9BnApIYNN0C45eFrmbN52jLP+1oQtgP1VkQAIXhkmI1kaP2M6MgEw2m
a5kw6Z6foRhXA0rK7ZO5eeSlv0akIPoiPx68hAJucGv7b58thjsPsBpu5ajwUBYCu6fNF+12RamW
1OjypRlTXAazmpa57AX5BG2EAGQ1Hhy75YeP3Vq+IbPEGcotxdndD8t23l5vpHSXQ02TFBsVxKFY
3Ycpv9qxsA1jy2h5pJvUPqZARzj4rb54B2jcqjtwIAsoNcDhrDs5E6XDMTyKAzFfBOtIo65QUl2j
MPlDslI+1sQqBha0XLjz1PJ6Gtdvc79wzgB+JSTnldOXTZyxcgzp9DLD8GTHN6q8Ff+s9lAq1/xS
sLP/sm1TMxGeX4cbuKnGi3G1Hn9tRSDk6qTd4x6RpeUzRQ3xQzfFcWZp9D6eNKkqy3ndChLgQSOX
SheV1oOLaqCdwzRsOwa7gSsJtv4dQJfQyfY+lKVJLQHYmmxGxRuWxIak+XxdBpRPMTGjef6fHo/d
LagO0I60yjW9wuvynK5XaK5q8l5qEywEgSGOScVYcbUpAikcs3IaTU8UXa1gAJZAEjKxM5k+gqnH
y3W+ekW6Tky6razTj1WOt/K6hilTo2KaHH3Xe3pUHomn6pazcVXvUZncUICHgTDzwP3lQ/CBI3qw
kJMkJz2M671i9SEj5HZuM//84sSPRHiWevWpGA4s/NTM7GtHyOM0cTJMTSlCx1KrrrKiJOhIU1be
sYzWPJWPY26TurTWw7YPoFrcQY0eQnLClIDwIV/E21tCOfnyJ5w/SBUjKqyadBitMQG7gSye9yji
+wlY1NWRIFgsqU2Hd+J0fH7Q0lJbm6cXA62R9F/X/EBhcw7jE6CjJgA251cDQ+0Q2BD84JEHCJP2
8tn8Xah2ekkAU5szJ36Q3/6Kj8pwR9DxHH6q8QyG0qwG8N8nJL33k/aN1pwD2oO4dc/p3rYPsPRw
K4lh0j+ZBE6CMIPKIeqBM/jSik3Pf46F/ihaG9438ErNfJxtY/TlnQDotlHlHp9upDanhJoEfTJa
SHfgb2ErAGRX3ktL0S1YX9QT/SRUPc5Fhi9OEmVzK9xFFmzMLLa/t++72XTQNDZJZ2Cbw9wEQk+E
oXRctgB5JOLxm7u+6UnLjx9bdSj5xjTMzCgLasV8DjjM0PjrdYflECH7NJbbsRnmqIT7K21jizO7
G71vTi36FrXvbnLbXJeixb2UysAKkrGDB85ez1OZnNVBD1+hxC+LUBA+OsqSovb7wSLBeErDveEx
ieJa3cLb2fHsPHnyE4hJQNE39Z+oPmcDgxLZlG0tLqmAg4FhBOztKmHEr0+EUTePHBZP1czIaDgS
pEDA02QGfokobGcOYjTnFNhtkeqWwgBzBtwg4+aTCIY9xuajlt5ej07RzLQPWnj7Dg6xlo4/gprH
BJDOrnZvbfvV5wyvc+u7QlvbN3ny2+2Bbj94kiut0ZLKeOUkK2z41kEa/hH3+/JiDfMiqlXZNR6b
QaMZwi0IxOlcZvTATszYeICwDmURJ38rAPGChknCr/jQOZwGJlNBtPZQlcOb7tt+sLSdlTPShmCb
V08ubp9cyOHG1u/Rut3asGPHYqHCNGSpciYpfynskTrperQdrLQRskDcZvoppqZ8oCrapTazRt6G
Z7It0P8Bp5EsApKnGzlW57wHMlqdFhL2sBSK65wgSt6QShKIVkaEOx6syYIFOtiMVp5vXR6G+Vm9
oxE9BqzjD4eOFEt+VGAX9s2Rin3YBxlqYi8sLgCnfimg9CP6PMqervMQhEago6eIg+Z3eByiZRY4
i8on0/nEgSDriuKuEbeFHZUin9uWMVG7DXFRdIH+7X1hH9YuO2xvXSD9I844qQmX1BoXhqOlwWBK
AJ+ikBNQopwdGdRxOMZV8yazi8YrWsb61arAK5hwKNP9iQ56NCDl08uPjgKjI6NxkBqt3ipnB4DF
d8kPrw0rvLcmivGLz/MiG8GeVpca/Ei7jIf4AONq+W/4VIWAFTkhuLV92TB7RvzzIGF04ghIXWlG
y/j36feHQHZ+3Aq8yICY1XQbaNGuwQ8euOYoUrGX9cBWN1krm9wXd89kn6TzoFtXFpNikRdA0l47
CK6nr1u23l0U4aagCO2UL87RhU76cJwQFpobcOKxBfi+eNtLUonasH3ho0Bd/XjuvfvcW4UDjSSK
UZNRKQX1s1zQPINu13wsSKqoJwGZC5BdTux7l/5XRRlYxuUUj9Epe17Ek67C15YHlbiRNqErtMpi
2Y/KZfRMR4htGBOci8MMkDiSuUeeAlzSYGnuK0M0fuMj3CSKS7OMXaoJuIEztGU6yBuvPO26X4RI
QUoCNZEv8T91OjYxB9+IvSnDyL2w1pRJbLL9kq20Vqga+jx6pAiW6lU2Ghtq8zvTnnDJduYPIrqM
eM6JjGhrrFbV79viw4dpUQeh8Fb2abDzr55XetvZ1DxbAbxIX7naDXK8ndqJKtxWGTJ6QBAie9P8
4LTnQIzYV2vKFPzjh0d/abw+zs8cIpIwsNdbK/Wr8sQY0FMYEk2+vwsYySVbSrkEgmWQznC3WISp
o+qT/G3pW6aRnbp9i1bwHb44ikGsxbH0eUG36rVa63AqIY9cYDA8a2+jd4omuwkR7XD5mysQAYoe
oX+jqkp5Zo+hrMPpBDZKUplkScD0uq9iqJ1FiFokjelXQPmuh3mj+DIwb/4OtzvuYqwwUkNkj3u0
vnbYelAFpeO6DOC5HjxNb5dAgu/Apnm76ykDIu3oYaDE2Fj7i8Bi8VhR8uvxb5t1mRjWTU/ypOGW
uGGSTg62MBc9/+pYfQDoGq39sk4fSxuQzxIBQRnuJrn/xz3hKv1SmtfzAScNHy4Io9BCe/tFIkDs
PFfKyIKeeZvHRuuVfh1CpHzfnZXBDCENvsFNnzYvxZMVlEKKoAsu01h/AlbeqH+6vjZ3h97zxcEb
DYpftjOmOGpBXZgZyR98LfUgBsBm7WDp7EqtpkT6A9hjrexNs5A/S4iiLmaThoIqyJFGT9Z47HF3
HbK9WRP64PKDpZppzkn2XaiKl82pF6HXjbFZMxjtGtZf1prL/TdhlzO+3gQJBNtq6UZ3Y3Gewu5q
TWXfCQXwhZq6s0YAIhbwgafh8TtyTGXfT6xdL/OJEe0DvGlH2503YC3NEu0HC9vxD9Snu/L0NlpL
l4LgSktpQHO/rMu0Uqahc/+EbjFxbu0ieWMopgzgI8PgEoKLGGIvy0UuZDx0yC/v11h7gX9hxhOq
DQgNPgzXRXggY/7D+hNx3AaDlfiwp4GnecxpbfMDVsfkqLy/8aGdpUlEbCECqjgOcRVBPizY+lJS
PskL5KBo3eHSXW7xT7VZZmlJybOdjrITanauqBlY1D2GaQpPqJxOusb3gt/R2vMzXYjaP7jkJ7mw
Ct+d66v0EY6+D0pHlZnOOODHY0M6DAftWVROeQZBbrZkcRYrSljAKpWVFm+t7GL3ioq11AgoOErX
SHyMJYj3g/7AxNqP/a/NAnZ9GqCT6jkSb5Tb1XrUtAlFjbrNz32E5iHbH2rFZ7Qe+HQweeOoe5bc
f1KeenDomHvHEl6cEvpCbrdGhlcPOSQY203IBlWEscS7PIcD+Sptr4WAUBBPPrg4M9NmoBVRpKU6
Ma1Mya2to0amIfz4fB7vfE/uhFxCRjNtjpXosG78g6xTm3k/+zSl1U6Zwy99c+SDhvb8y+Y5VUhN
cQ6liZW0kxjMZaQn+UTL4qbPprKXZ1li58wrSsaCONk9lO5nNZAek1LJCk0SfcPJSCzvtIhsKfGm
79VLYdRgxkTC+iH6X5h1jb7hbh9UxseWCdHS1tP7L34zWL6m1z7AeKCU/UlxdZBIaSSBOTlSQbtO
qil6o+TsTXS0aL7ObBAWcpz6lsLO6tRh5Ez9y193ypCmFFYJb6eY6HZgqepPWTnAgIF3gLp0GTsG
wpzXY7riTRy8n6GT6IkwzGE6tdXbILfKvboAOKvTFE5DPHUeoDKsjyFxflNMsXmTjMzb/chy85fZ
hbS1F0z3gOeOlUSRRXyTRRQj9+LwyOmgrgsIxqF+pYiDZP07UsPHJWmklpE0fzoCZQ7VSrbZDKC2
fGuCZyUDCxgGufRaQ+NSUxV+TtoLAJbF1jds9iw4oO+9VCsGlkSlhhktE1x6NP48DgUYvX8nC9dJ
5MQquIODI3+KR/PMR2Jo0uv7lefkfJt1lmyf8iAwErHb9rP89CKBuk1W5ULD6pk1lQqVUGpobf3G
W9OLUZIkgBy4fy6fdvc0cCIQaz2Nqv6KBPEy7uw9LwxMwIMzhiJ9OI77JBOaOTucC903f83s6YGY
zV6jNlSkKvVwyLDmwX7ejO7sgu870/L+AzdRXc7lHoftHPgXPiY2EjkLhN96lcngkx14Qwm8HbXy
fmfor4DxXz1sh1RLWm/6xv0Pr4O8OoWeVOnmBKgZL79i9JSnSstZSzTQKNISg8+0X30YSr8D8p+C
0mdxLG7IESIEAU4W3rw8e09rHXCskVzI3YgIcHOljboXk9HPZaqaeCymN+GsCeJpb1KVh/UlsB/B
EdBKv4tdrKn3dBKgm2dal6OxqDtBYP/5fpK1c4ZUF7kJOdzuYpVUZasJXkirM2+owXzyi7x/1XYV
SPZTl7IqUBll8Nl7kIp5YBjEyXiB6hUgq3jVQts5N3oXWynW+rVrO+QiGvkxozGkXvu6NGEtGKpU
TSEtWdaDMhVg6OTyvQeMquW3ZwvmrW4e+p21LQYK6IBBcpEeSEfSA01PSWvbqwbOR+7tNw/2uwSd
Bo+iMrAGTJY23Je6wUmPzw25K0PmnJtN+2P3JY72jhwDDqJ9YMyO7691n5G+U1zL0uCRqj7N5TKR
o3O8hDdqF/uXaI48anaKcdrMIOBO0sr62Rxxz8aC+RnZFKx427F4cns/dNgMXTY0tPS4aRo119EQ
+q5FYBN6N35avAd63d+yxMVOE51KXW0uD56FovQ2evRfjcHaDKBgDw8Afs5hPjsPKloaEXZJke2q
c0i7STo3ST4ap1mnIEeWz5f+pqPu9ooW+fNjrp6qw7wV2eZfc+18Qf6OzeIqVvgYJk/aDFr4DO9/
LTqEQHmi9AF8TdZeto7M9gcurkiizhWU2M9BAMYz86WiJfScdA7M7lZvNYI4f9fZ7we9AAK+fCpJ
GxZjdf7pJCTV0Kojzeou+Hke6Xj8kd7zbheL+aB2kzNaATGDfe8jKhBbiszcn8dEur2FoqHblXMs
vmL6RpW9DV0JmdQ9BsBRk004SxG2R43o/fc2bM/rHbyrDYt2jCFrAfql0FL4wqXIOlJP5EKdi/1O
saaFQgUZ84PGeyrw8Woou1seGmbXBCam97fByj2e3nFHSgGKYY2If+Xb8CRDlsRhqHX01zTNBZwV
QcgUoNcZjvAQ6lJUMhhJL60BPNg1kQbkZkbLM3MNwnM4Ok4HYuJs7KcszSF0nXbLnmXYu79hluH+
TuL/8dIfhfOxJcnxTkEr+mceMfTpIqzo58NwxfhPvXnH6uLaiRm2dJd+QYxzfZcmHwmq8JDP2rSy
QeOhSG4cLrkf+t9127w4PHVBOSVcEspq0eMgqwT9G8zuXLU58WOxHZbmJsTzUArPrDa0wYFyqJDY
c2qvG7/ReDfnQobLIjdjFGtLmHDm1U95QS2xkibAL64HirhSwMNWLo8vijIyXwvGEX3DfBM6iHGH
55/iV2tFqe4vrKEEtkFDmODpv6ucUC/UyitpZisukfowbsXEaYKDo1W0Az5NgHqif2JRmywnUr8K
KGizWQqRRmHOpPMpziMOcToMAlWU9iYuOQTcoM6xhobxfo4NL8hiYKfnL3ul0uS2dwAtpVIF/AYS
QgxjUBX5K5PHkq8ZD5rRnWDoIT374PSfGENMatodzr1PELWTFphg/sHqNoawKq0xvuJlV0R7/P8B
gWHkkVUD6yT41dIfDCpUyv0bKJ7bm4we8NR01BYtfR0cCr2RLWBkwwKZ43hctLBzEAMKb1FrtGNY
2ix+vHS0kAmDp8IosHVEiALrAJN2cjsSDkY31g9L8tFHpQm4PhiA3GNZO9oygZYkvAgM0soYfE7h
9KRsQmIkT+lQMo51RcK7QHNDKBfaykM+sav5Xm6TYAoXsQ1IXzs5owxtwZj7vOKwSwRYFbj9Jsk3
wJv/tyoBuuhgRAEc7UXELp/jYGV1NY7EEHe9VzFIDhafLbkkIwF+WH7YpEP0CvJodezynH9Twnys
4+oVB1RsSVoS0fdkD7coiZBbnhsT+cU0IK9kqgASpKUsiLO/NA1t1tKo3Isq93KU/0KQUjkpr6ya
HP3F3C3cvct4AH8i2w1PJyYPxHb5Ev1845FUUmE3cXvb0cxtorzuZB9p6Q/ebHhrWp60htBhVmG1
4aBNtiXqQtXldyw+FEfd6WBX8HGTthFPrDQj+RFDuMJLEQ90L5O8i3tFod/kmOQypMyhLUAIYV5p
QZupCij2VYGZl0jrsJsIQLiGDE+e2cqcR941r2LBfJdBcXWvbhxFHfAeHl8LYlRMSYhAsaGdRreE
IJTjfUvLWrNQLm00MywPE5PTj1hgJ+/uR7qfdXNDM5bgNTamO77nOv4lRJOLFsoR3L9t/o7zCTd6
iP4uKRxNK2zbZ+DwC1lBd2ngsBO07sjzgVYSeT2dp/Eoc21Z5PVfeNFYWp8ql2nWeEwbkI/mhazX
HuyqLPiftAiigBYk+mWq/4XDFgaZ2XW53ejIlaX2BYymUuV7uleGRiZskoTGNPe813QFb+KYmpvI
riKes/cPhDyiOgzuTQpf62EpuAGQ7fMMTZjn/hPSuQck4VwQ4XGSy4nQhFVec7+AeUBcYCy+8Y0M
Af/c/d7qA0KWui4MLHxH8eb3a+nKHKIJF/x5H/EB4o4IUAtEsAvbXAeK/zWwGsaM/jPT/O8oV4GQ
yGluSZa94MMuk8lgjvkCv29auoexlgjA9/+ngKYD061yzAVy+e2M85/qt9K3LhwMmz0zHtDOs5t7
9gxmjx5wTGcsjhus9R55s7hEXeNvsvC0bc8GYbx+QxF6skh7EFqA1bd6iTIaZrNqh9ifaJ/gsyaN
CAjLT/HPz4k1n7PA4FPGUMcngw1L5qsJLnQbKKljWt8HPA2Gv9QYGRoIsvxqSQdow+sdvJ8Nxsb8
J9Gg/zsD72wWrVpMd+Zu+NOazhnkc1dGSATzNRTUAYI/VsB0o+r1lyqVjNVgqwao+AmdvkVEMADi
/UPOrmNVzpsHAHA/EaitdkCIcQx8bNow/YHXNnf2B4B3RtXYiJpgjgXit8ItMnyIK4jQvS36YEhb
kYaQpYVi4RZG6cs/rowYKLfCvLNeTuBeXb1+yKDl0t0YG/8/ItE3NUE0X7s+3T26iGZxr9YTYbtK
7s2WmqIcokT1hMaE6RSd6y9SneLC35FF7RH5vrmKbiBD4rKSJWHRezw9NnG6es8jd0dxktFVdTF6
mwA9FZPhMRciSLmtf4vh9YjEFmKYQ4ZjvjiNXAmbV/EJ9JnHyJKrVBcbEAbpBpc2tBOw412MxJjn
CFHYhQ7Ra+I6URsZnvTgu2WXE3MpYyijz9t1dZVKa6toYfKGjnvjPsDEQPNXnJSka+PLbKvPFw6E
RmLSRPbwssvVe4UImazq7+3u8XghryGf1MuXS2hulXBlJiPb5EKVMvRET0bAmiGlss9dHCADqGYs
3IYFnl6AJudsEpPa+Uf3gZ4vtfRp3wONEmVvtO9ESNIPSZCzMMX/LgosLTJumOU9Yaa2mmWExmsl
R58WFaRJzaVBMVlnbXstvkNHfLTmGlhtl0VKIN+yeCxiNSvjKt1DZvlV39Ev7ozOQ+9/RYwEG3su
YM/lIe+7TMdzzRMjrRijeZXO9gFrVqqLYchzouEUOgxz/Mfk+8k7YqUvS8NLgLw/RIw2xRj+6gV+
xwhE/IqViXFxcSIA74/ccQCbqnIt6hJgzxh/vM35tbhQapPVqmDST43TWhaW1QaTgNzgf323HbS8
1DjvPAJdgQD8zz5XQO2CnOebkh5sWxrW7ApvGnLhwdKJaY0YZEpaDok+isJhLV8ECrfN3uUwyD5v
cVgT5Jjh2dkan0Oh+rbZtT4KI0yTHIQTXhbW07G6Cl7HZWSRK9Syso27R+0CTjr1MeDNWrJF9nsO
qGcDIxiWNpWf/lmmbjyPD8SuG363XTAOT+Cpv8s2+mLCaCh2E7kAetJTIuDIPrSCxvsDmM44Dt/K
EUcAQp41zSe6VygMw70WNeGBiU0+OGs8A7bkOlrOhfPAxtrXXnT+7IaRJzLdq7HotqgTB+o8YNe/
yMCTxoKbNJo+j5G7ZFbzBkhMnsqd+ftcPul3DtK9G2r89UFoFddamX9d9JXCxZF5oFHQ1qcn34Bg
e887XhvznZDeKa7FT8KWYW6JZdCGsa82/FcURciOrJWKvAmZYHXuKnIC84weuQrzRiFTcT5ozqUf
mIMFlQZMSAn22ueEJtbJG6v+tQKdCv5DhM7+UtebwtSsNMzBG461GdlGRoWDDVZbqHfNjFYvT+g/
FRn0Nd7w1nAJpcGqSalYmJfr6d89+MYcwv14Pp9BQxohv6PhvboxMEvr9hk+vg8V0/1zM05YpLwE
nDqK+oI6+DHU/gxJRhKt/hJWjNch58fUAv35m+DrxzqGPm7hRtIOhf56OEkhTfa8HoXRl0EEWU8q
bKTSoOP4maFhbhfiCpcKirretDArGdY6xcpYmgxnfsVo6S/5vtZzvua8FRFLMZhVmQwSSftrFZ2u
kNeXAEmGyeugLgTItAAtqvIiLmqKEAzKxBLV14dLZpVupjB++JRRXfE2GtXdOPm2pnvTZEglDm0e
IHevHWMma6yn8O/+W/p4KbCpC4NR20+rIPQOcxZyxnXc5rqFDoPbTEWeDw41AfNk4Eoax1oSMxok
+XcF9zAxJejrYhwxJAyrpf7AbuaYmZmHIv3MAqPziEPPsaAJR2GG/2EQFwtjHHbmFRAes+MUtypd
8A7D1/R1I8Z5bE91qHej55oQR9kopbR/t8sbmj0DfdXECqll/DsO6aYtJ7naD4Gag3bWfWaX33dm
1EqDMIHU+MNqQxF7CdLuRpy+nJmL+SDBtp39+m0RxQp8lgmgZJPB0a6XhbNwyWPqXV6RepY7i9T9
m2asG7nobcgqJVkBlS0XFPJiZrKCGQZcjlU5kA6L5f/LLgP21EmegQeDaV5c5aiZy3x6hMq75W/d
rmXrPwk9UcHu66vFRAPnmH9lV5qWHxEqkkbkX+bz6G+GelaGq9ciI32r+IPYJND7UJDyJ1o7Xmm/
YR4zcgpXpXzuf+qxz8tHyLYKWaQD97xBl3iAUCPSNLw21cx2Jiolxg2Ng33aVPFEcew7zWoOctrX
HJYSqADIfbxrh89OB4/OoWlXFHzZMKk4zfm5mfCXbQxZiREqnERpBvusHGTzQidWqAUCXjBq5l6t
ADWOYvI95sp8uS/aoye8CLjoAR+iwWHzg0M+w7u0iZO5nxHOkoRd8XBeFlWyW7AcBnDQZBpW330Q
bUhxGxtjl/T9S50YM1ebJiE/AoE+gxs7EMiqRNZtt9++1RSnm3l/xncExH4EM4NsC4+vTPm7kigw
hSQyMsi5EFEnAMbaPEPNwlV1qL+mJIbfzqgX7cALXQD3OtaezTEUR/7Cjv2H+WN0QlGvkQ36HgRo
OR1at3JVMDK6oVARvSIfcBm5tfIB9Tf6FhKSBla7Mf55htkIizcS6AZVlzVXe2IgCVfYIxb4xieK
ddHS07qfbU+x5YpgXkmTcIlcycDUA4USVHN0Xysv/wjSoeJt76ktmE4Hc7ebAKQcx6A/Ja/Pf37B
ceijXgajRv14B9p7B8flBV59C39vuCPeP3P+XHPrClgAVsZLIRG30Ir/iMDjhzvLuSdubn4Z1rv0
E06jpFWJLnKyziUGqWIQtLElSDILqV+tLGGisDEyUJDSDr5qmKWsT/sUOHdpUFvrnFDvugq9Aczm
t/RHepP9dYx0BBKlT+vjyZnFIoGSmVK3A7H6g4+OeDH+f3o4C94pWvxR3KkphOHcYkJo6ye/C/RM
GkiBssas5Z6jDdvqEaPpyNS3PMNQIOT4fwdQbcqP0Gnmk59Gn8XYNPncqfYIjsxYMoiWPMVfYduc
MW7I4QmS7GRNVQ3V0BoMWtuQo6kRxQ77IjtsyImXQFpWxSMxZN/1dr/9XF2a4yIerS1a6chH7SA8
1WBKMeTTXsPyBwKYb/0CFaoRZWJ/ow5dDIt1GB544ppquTJPjZJ45ABvCTvONnxjsr0yfvruxP9Y
cBBHQEGCtieopjTdp/b5FwUG3OHFu0GyCHzxiEjqeMkN7Q6U3nq+7HMpu/LD6eKKZIOsxIZgtw/P
UIiMGVO6hPRxDEi314REn2DGi1PTd2k8hBFBnSyzQw56dGtqILsYix6N0hDf6ylv4xVIS4qH8hnC
v+jjHVhtJ3yiiSejnLiq6d4Qvl419ETmUcjIq5/nT2f/drh1jedfYNzApkn8Ga1Amp1QCWsP15uB
vL6BEFNqAj+ngUjGWkqFOztduqvGF//mr2hMv/19Qwhi96idUB8Y/0BJaHTGHjidMfyQHxg7U5ZY
spsQf8l/FwOHlt4tKs20QWdT5IZw00KWezKVMFrkOfDML/kYkxDuBsHC4fD8VmFXUyVjyc5Zhbor
gcL4ySN0B96ijCPNvvv5EHb3RulpJ5KFCCZe5AAt1plu6wEIryeSofiKyEZkFSM2P/IfyPx2mMBU
eI/rP5QlJ5sVRugGkrtDT3ikeZal/AO/Box2r4+EbdixV8C6IJO1mQqpYzMy590sNXyIpobSvfQx
vxpQVezCH/3pYyp/H2DIAFzVUtSrsXyhdpaqWpv3Bgaw8zLNdkd4yfe8mO4eORKg+6X9Dvwj+Eah
+LObVGHJAJWaN4+Md5FsunPGBoVhT3WAoSFN0cLj9R8mB0uuvUeTnpG9w85hHfkTCC9LB93OPvwJ
i7ThJbaTVRA2Ka4VBAL9WS3Lr5lWUcoFFSRHWJzHi53e7RUXR3MWSfZe194eMnCYegKvtsq2z3hB
WOMAGuEQY3HuD/9Ow+pY/CiHCLL+KNQ7Nsm3FY0sLnIBX1Kx4rX0sPvf3Xe+FcNm+0D6ykxSbmX8
sSQsA1sImu7gtzMmztFKDM5OSUzr3iHJVpDB4ZUH2Qlvq53vBVakAcKOvXhxlXkIBGjgr2Vzp8YC
FkETkwPbkXfFoeEXpdFRcsIM/txsf/8KjkC38MoWov14iBrX67UaZVJvMBUH4/eVLmsMbTbnY8gE
DghC3DI8ajaaiKOU3RPZjjx8SYaSS3RKIdrzRo7GUWKqqaTE94SwNXkL8Y6u7sNMOx0MD++girRi
l21hxTlfunL+UeDm3aXSBvDwlk+KxaRrb5toaoZvorECk5o3xO5CRm0I27gW4Jn34jHuqFoi2A34
IYhvyYz0DOPZgx6qnpEns5Q7xApFeDI37xZyH8sNkgBEUZGz1ku9QdzhJpXL/fGdEW6eAQ8pEPzy
eP2ZijS2qKu07UlcJTgmbsFVe8Acj0X7WvrVugqvdWlgceyXpSXslFdUzsopItbhNVDRi8mbdcht
vANCD8C+Y5zj4uHUAqo29OfuiEeHkOQOExmsHjojDKzoARa37tuVcYkgMH+KLoYb0e9aH14IxOQc
3UW74Z7qVKYipHgu1zzOy98oAUqT0OKxRV6tP5NC2ydwo5eJZrDScKxoRtyg0GR60oRrEjRMB1m+
hm7UzeVbbly1pMEMyCyl2OtBH5zL8fbHvc3vl0EiZVTaD9c+ntZ62sj9+Vg0dLrp8GCtTYI5IRWL
geJxzVr70BIb0GuiGoHmMtQ7R6kbLhQSxFtd/J4oOgSr6y0LX8fa2W5kLdJoLwgZsWZR6eEtga8U
Vram+4FMeSFhixer1hkdSI4HkCVxn8V6EUYGvWD9jpWnlwaWm/C+UychPsP/Unb6zS25aUdQsNU4
uoWAlZDRHfQWNtiRbfrMomWRn1Q4rPeCDkE9/mtxEYU1811Rdlm4h+tuDR+PL1WcrKKs9CMydNWI
BTpm21DB4lU5uDFXfeACzATK5KNHmcB2SfCCABQ2O0v/3+kPlZu0Xkv5mHZ2lUvW6Ncx0bYixyYH
nOVNR5QcuZDqYJ/idxok9WdxHdikydQF5PQHzRKr8YV1Xx6EdL3qyD9FQR3P6hVqC62DarRkGssB
4aFA0LmrBIZJ0cXE89cLP4rNhinvLlHA8Efbm7MjI2JMWDkXZB3ijRFMMUOzzc4PgbKtpmVaXmkm
bAMUCSmErLELb2OKMSNGI7rM38+VW6d1fBBfiYeeFlVAqq6M7ohGvwSFJpWzGY9iOUvaTcRKB5Lx
vBpWtimIHJTtDG9uHlh1+MFy4GZ9IADjcDZDa7GA7i2NIdHkKgA4Rv7r/PqyAzDAutHR4Fvevfuk
AboWAc/tAA1ICv3qpW49VM9pd6zJ8xYmsvk4nEoF0UD6iNynu8kd/WRbv0YoxYYLw9seWIRl/UT5
sgYoWSmvDEq2LxZJFWDw2vnVK2XgFCM9Innepx/GIa3T8YfHl/P+gHqNE1jCYXR6+yiZyEoEvAfz
irNv9ITgU07AlTlSvnP66QYog/OLVEjx6DQTBM5NAWmSaHsbEIcY4Vt8Nur5/lJumaXVq6kKEgJk
86FajnV3Yg7RSWS8AIO1ALKOnwOIeEYtkEJmRpELtrif35iMHvFyzhG2ZhYCWAc/WT5Xg8fZyP81
JSFwHKn19fDOqLA1wbmjj+9uHnbhBmpST9sKaT4KKswKuPJAm4C2QPejrsb46nXa0R1nC205ipuZ
OojKMrXoZqe4Z+x5pDWMoa72bWEwVZdG+KmP29XcaXGsfLUFuoPKkMUCe31qAm2RA77nTuBSuax9
Td1Rrg6gDb2fm4clV3WdrhLTTBrYM+fCboweP9JzRtB26BNICsX82Dd6ClKRmsTuhsfQGEAACOdK
uTEob/VLkodXSizJQQURpchtnxV4sZtbn2DicPK2hB6oGFhHOlmXlwG/Km1CTOHF2Yh758LH63DI
L1htn73KVjX13Eq6QOYeLQJJ+ZGJ1eDosOvDvODrCRM00oamXBlMHFbZLSovfpqR4N7hYz5y4ng/
9+CkY26bktvL25gxuQ7JYtnJbCHwzDTkcAPealsk1vwyG8NF6RmzcPAa8zYgFG0sCn5L+QTyxq2k
wxLY3/386/Yhr/pVBFH/swHMqOZDUM/7N07VjToguoUT5XtMaDXgxyOq6Qo1Oad8nPHAF8UVplQs
lwu37zpOcXdajItiGuXzbYvXTBaSVV118eyJ0V6qNKhL9V5SI093Oe+8avtscsmLXFjOBt/YmUJr
+fQddGvgi6HQvzRQD9qoAFVGk4rOgbpR91j86Sdai6WAM4ldP193Wo6sGvSEj/YoYBSt7wRnaukI
thWNmbMKD/IfkelOaUIA0zOEuxMUz/4XQb3CKEzP2PMR0fA3Muc+eZit7bf7Xf98MlYdb19STQoF
pz7Ym6qbJA+0NG+BexxSA9AdzurptzQt6DyiTInVfvuoRnrkj2t9pfiZOggnOCPo9Sw+TWF+3iGA
tY1fQ/hCcFuSqqcUEcQUmZh079ZcBmpWzgth3iHVhUQ6zGIZDw/ac1m4kL+iu1/CKz0xZnBopkul
TqTcjZ256Is+P612Vqg+MyTTYN+EwVW4qOPxVI/4YMxMMfgtzEgLmNXsHBv2Ig5N+nc7AykdsVk6
rHgVWkfvsmNwJKrhdqq8QtFmlqQPhVvWm14PgJ8OK9OpmdxgvVgSGpHZa3a5t9TJ73pJqiiqOFlW
GwsapSGqi0xF1bbdeXfuw77GhUlqlWO4TqLUX9i4HCG7xeVnfedrC1Cd+uD5JAJQZ4x8Aia19/Mv
mo5+CWpURZvIHsowvC8q6YUAsP9Vs9YL21nsZ2W0C90w1cWr2BQ+bfUfnoWS7ip7l74v7vs5VgDC
nnOjNwxycWnBpj4HFhE07nRX6JUZG7KInYuXnYKi6IxXnFKQ5usE/12KWYsa88EKKixWdsayCrR7
Nu/52aSK5n2kNdCCzPU8C+fI40ybRFjEdud9HAIXhcYv9oAkJD4SPAPPYWM4GXHQXFChVxZjTeW8
ANdKW9AddkzcbNvGiHGNoXHjtTyxaCSx01a90mjDhlqYjtqiZSZ79KGVzrFKWGNMhKACMh+3k1Sz
hajZSaAWdjjjo5CdmYOQyrbq+sgSDzPr3k9FCbboXTj7A4SUnuCsxEymQtpAqbuLqt1KpaXcBuFV
m0lvSWQNFrifUiGY1ss+SntlMGDuPXaAOw3Odi+qcZQnum5b2stOGEF/h2yMcLHwGP1EZgDs0E8Y
4s8ra02qCIjuVsEZaEdeuCxraP7xL2CKBKu/mYlEHsl624a2c9IbLnZBFRYYw1H0c+snIMgJWfhu
nhHDGLEXY7DAnEWl2J9MoT7BQgAoLZE1+EviZC7FhZM6n9Ruzwk9u38WHhjQm0oB8fk2ROvFe+tG
kiuhHrkrXoCE0uxPz3dpwdWNWzDvPyCPhSVXZPb3jGW/UgCfO/CpmDUO5adMaL5W4rJTiwd3kNPx
uJW2ApSaWp4EjU3qPMdNszgCryOSRvKAdve2iTxVHgPWXsKEXKR9O02RGh1V4ubMcQK/9AzvhLJr
YgJ4uyM3lE289wnj/mNBGroHbSh3kW2OJJGaZ5f9u3BHQt4jkbG4yF2m06uUdK0lym6SHgoassfy
INIxVqXlTAEtd0oyB9AcrkW2TyxFtETgURh3YjDqvGgzQBeRMwBIBsiC/aO3P602M+ZKt3CFLOEm
7H2iIloD2kMHOWHS7Rd++/zy7WNidYbc89ABzqelOoJ9NmKyWQUbCG87y6i23+/ZozN7VOdtfnWs
jO6stf1FHvjDL4BOYO3V/Vqxm72+olPQ88jVkqM5aiHl69XiPDRtA51Hj4U+WDYVg2mLLSeSPytZ
0+YHhxGsho3lR4SHTsSyjK/4ycMR7HPiw39eU8G+M6nOjhYzKU/0SFsd9LtQ0WLG5mOcUv5m7clJ
hIS4NzxbU9uNkM2d/Q/9rAfs4p5u09qZDU8eK4bkhE4h3kQlWXteFdHvEZ5996BXi18gyYAqxEsm
P8yPf98ibgAhsJKRitBXmsND4Kcs9PPdF9j6YyO6Rri6ejAvw1WfQioZXNFvWNGHC5H5IOgpk/5N
gv1tQxcwC1oGWa/chCFFmW4MSXp5qxCBpqjn8ijfi6i8h7Czi5dCziPhK5+zYCQO5Jsma4VgZ6D9
/HWDYGPblU/7RzfwIHXudEidL9fgZt3v7eXdsHoZboUWhPmv5rrf7JO66O1XZNmVMviPqTZO3sIK
fkxnMqunmhRTq5WQ74WRPrv2xWdrkkgxLfhL+uJg6KCbdrYK3fFKQogKYkWSkkWwIYipv0tj3aM4
0jv8Q7t085B3rFTGdDq8WaPjwFABX6LueWydkpZdxh71xCJ09taofRIaSHwmzaxkD+XOsiUy5yuP
4TczGClNvan2qIj3TDfwPb3LPwdC7WFQYUt5s4ayG1DLGWZi7QAh6Ez01kfk/s+u4fYmYv3DeTE2
ZzUsXWP47G7Uk0zT+6LLoIWVx9ztLNaZucUNCHzHoCalvBeuOlLfKIImGIZUq6z+tWfGZUiXe6ar
5dUzxdMKtpcWL491HXh3eCyxNc5S8JT/J1+8I3lnci5KZX9CxuGTnFuiL5BkbeXcynGDQIR1dJfU
wLeHgu5s7bqBmLYxyFlLvuNGBpN45bkIuzhm3VtZu9Aap6lvEXU+/zt0N5+9sz6AivGB4I+FU+A/
FrGV2SVsxHOTVhWN7w+zANLwHyoTR08TxQE8ay+PifohqvEqbPpxogrUylkEYgEdeCWmKG18drlR
87rO5+G95CPvefQavnIdnzXUHsIBeiPQtOl8gOTkHAJocc4lpEP3sR73jJZr48Tlb4b4tXsGW/89
7plAtVFTXpAqx1USA55MA6EH1iYyXJ5dWSc/5mcvin81CHlubvMpYBuxDrV0jx9EfvRVWlB6UcIu
iFZ6EdX7O+IkRA4WgYBRaP+1/3g+6GLKdvDqxanKJ6UIWOpIztaxQ99gUQN/py89eZ/0z8cLn/tP
4KItnYeJgV6E4REC/IQXQzakYGJvX4PI474bljO8briBf5eE5Ac6cToYeM4eYa3W5iqDnSIM1YqV
7ujsSsA0kRoL4rcrYRup+rKFC4e0PO+v8za/VwBj5v6bX7L0/lSx829h8K1S+21DZnKX7V+BtqLr
aZqeZxc8iK6uvOcbOTM6t9xXtOrXUY0h9YELg/ukZVUv3C830L2pISEQ5i73Wy/U3H73QHjigm3p
1m+OsyjU8ZA5FoXC+Xflh9Wil+zKGI8eIPjuG4Dkt+9zy9xOhQSxUrAmpAyg/sO6YlroB/nl3iqC
H8Z21meGT1bwd2Nr7Y5DW0yB3f/x9Raekw1Oh+yU4KTidzHZnUxBo9oNBXKOQKpHvGRvSdz70ofo
3Ws4ArMpGLW0TG7AxCJmqB15wt7+STltYIWNJiRuNIZufXguGhU2dqKQ1TkRmuTjARpOV14r2DNX
SaDiUcTNvZm3dc3H4vwkmTsF7co+iRVS9EwIFT1R5dg2OMv0VMNubo9ZKCDAKWLvrqa+vIeGlJpQ
akx4qsC/Gf1KCb0W0yWYJDszlsb1GzHnjxHEr4K6NyWHe1zIPst5lidNvYGIYEo10F/ofrMJIzht
MCoi6ULJ6BTetya7dujz70k0fJ0fURgoL/AGI1HDamJaqh/Iu7iZrWBGSyi3XkDKfmFmWCuM51iQ
qL2UOVl3SfUClD5vhPB0lJefysf2IJ0onF9jj26eZfk+eMsFbGTAr7wCKL/Xi7okLDFhLdizzZ3D
5DjzJJSlGPlfi4aHf1xC6bGV79pO2LRhkE6kr5bfmN+NfXyOytXnp5p/b5SckrQQOVkLyPVM4k+n
P8btEbi3QfS71Dzb1it/hBu7qUsMi6FlZPoCG+ThaYfK6GS/gaLmBeS6VFFhbmVibzDHSpZrbrx/
EBnlXxu6HnmtThAhq7YvJspW0N76X/fX8+0injYhx5hL6vyybD3X8Le0/tBt/2ZdIuj9DZpmpUVt
rPs2ti7kpkkGfFxCBw3l16vGNDKqc4Afk3DKfq4noxGWz7a5t39wtJSOtl3mzaDk/zBrwQkle9ia
cyis/+GtqlWFLdujM12KDTjjPmUxyneh2ggpcGzRb8/3n+GbAu96cQ0N2TxHYF9x1WMtb6toW1A1
/5zWP6D4AeGPl+o151auzbDxivDOJcsyjFukoayK7qecPX0Sl++/3xtB9Z+rG4MUjuAk6D0Zp9I9
PSd6sy1pP1r/fVhVZ+/heRvyL6/J8njs7QihC5uIW2xhvT00OD/hFyUi9TYzALJGFXOBs80OCdU/
txV8c635XWDG8qV9oEkLDQNwtVDDtL35l9XNP2nKApQ2X4Fgq2qLyUT/2sTV1vco1sWDov5vx7Q8
rE0b0foVelNRXXQSZedp1DRKZAKB0TLDDBcsoUVnmrQJpaUa4/x3tzEtTxdahpj/ck6ms0cPIbJw
CS08p396kEpLNp7UjaIYYbVOoIndh9N1eeH8SE0yODcBRtpQeH2rVp05IkFKytaRTQV2vyDlINQJ
aA2IATPwsB0w3OwlWNJDG6mD8en2psLBkIx9Og0aQzPw4AtIDZBC615N1WTDH+LB5A5CaxynQDw6
DjVrkc6wqUbG5f+OYrteYeChJJeac8whaSiFsCO4LHFWw4e0vOPP8UFiLY8eFjXWZHW2KxRcPZRu
1kACXNPA82aCO7K1cxmBYFJeY0ADqPmp/B02zJc5yKNBY7UAkwG3uIdr2Gc/mg2ayd15xYkJL8pZ
i8+JsgLRl3n3gBZdvY7MGnEUOez8OgrZsRsLNYyAV6bWlh6vHOU5TlpmVERFfA5F6LBpiHqPIA0s
jAhpAmRp/RUfAoX2ryzoStPhTNJ4qO3OUXd13+fJ511GLxPoki+nR6XHeyU8xJiFD3pMEDAcy+WZ
DXZH8WgQS6yOap30RkGYlqf/uhKo0MmrwC4jvfDPE3FcKLQGYfyAY9RRA4ZktL4dxpP1CogY/xBa
URstvZGXCVFfgPyh57WpAN1wQrvlqgN9Pn3J2Mnmo3ae9dFf894WmkluFcTK2tq0OWDnCUd6mPLd
6oK+0l12AnggtrR1+PEpMqOmxIrEQG6dqORYoqpRFQ39vguXFeckgNcF+wSbeQn0tH0zj3yA2uxc
1NKbu4gE2Iyz4Ncqb/3KE+1lIjAeivTcpmMoeNh34CdaBpSDKCDkmvrDFar6/NmluaNV3bZPjMSE
e/9mEvY9skM1zpyPatGoFV5IGYA/YwaBYeGBzyppEDqzDKBVSkuvwpz6tKoIhXOs89ZANC2mp/mt
Ammdshr9czqf9uwIgccQujlh2v0kAZYMwkrorw/Pu2ozMvCL5++Iv/Szofx85cDEO/8QTnXCr2Cf
/piUmMQGS4vCTp/WI6FWRgml7onmSOU5DDz+jphSYlV2X/tHITCGtJIqbnBTWPaq1D1Emb6zASay
/4c3TMl9dgKKLqBOZj1Pk5yq0MU+sSlQ9mgwbhkA0wXb37lbtGkvkAhRmjyd3W64e8uN9kJVcZHe
OOKw1S9gtiolkH3EYx+r2l2qbV8mrb4zJNvPW7XbBSI/qOQ+dIn7R8DCRVXwFANJh0BDzcCAL9FF
WAW/5qgI0SGpNUz7TxvO9aAbbqoSidzE/q8xO5A4dmp0d5ICBAk3AkXCJMszFAOn3rpBgtEzbzAq
Aq8XHcHopi4wmFqByHiKB5ovmFM0vEG0fa+YgPE5vqtO0ZlBEEU+xLve91WkxVcq87+gAM/vAKuS
iBUz2U8OtozK9Q4Z/mvGIA9Vcl0EMyHf0BvMBteT/Lj1mLVIb2vzfa6oguCeqaicllx/05hsUaBg
KmXUTGf/UjMAkhsfogAXNbfpgiTgpOZtXWQlxVIR4CSAOLcMk9rohPRqdgGTw8zQ4Xk9XAtJFx4G
uF9MpS/WGJTaW6jLlIycuFLlmAR7rnybNWHzNBG03Ku1Bm9U2Kl1kVROhPlzM2WDTWBYu99MlqLX
V9Xo6Jj/pcd/x8K3jNebdRlKV3Rdsr9QdqFxifab/2JarLyuLYe6/8LPj+QReUOALN6vD1eZT1M9
T+UrZlwhNaA02OhhUqSUc7D1cKVtM0GGRHn2Pr7s1EfJc3DfPpoLcYu4R1timV/XupAI4Xd5QzSp
iq4hVxVCBCrFMH8xrDiOVvFogmKm/EKVyU3+i+PwrUIFcSRx+75PPIQwo60zygugx22r2KeoO/mK
kV9Zcf4uONez8CJig071/pY2oSQh7PWLnnALG9UIjwg35Ux8Cy0R6Y9Vv8Ucvjf6GivMeM26EMZN
RWWVeNf37ioA9IQZyEFacwiOn7i4wy7TvEOBDsKxdLvDq+N2bsVws9HkJ8McWuWmXil0Qr/tQl/j
k1DTOJ+N0duQvUOtNe3oX8Rf5K05wNiE2lYEs3tEZYIEAFQWqXPH7sU3j/9ZlJILLjUl4f1R/0jd
jbl/02KGK+umW+gsSPP9yqhUOdn4+t1Khf+mvmi/KpenTq/qsojpP2reNsGCbFLW+BmyWg/fgUH7
hLZcPe+IdrquR2l8JIMY9LyfVWPiU4KmN2K7LATBrTWnUkvfk/yIndXVNKaGs+/kJX+HZZ43lgT5
QMkz53MLldlpG84xADZSqSpxXdLHOtXOakDju+HoGSVcvEzU7DGUaqpgjOs8p2zxEjS/f7RV3ct0
ZNz/QDRV/EFgsZWCk8fN8qD/V9GGA2jy2qID3wtWfwqwI1APcnA6BScKtRgTt5MGYB7F+l9+jyOK
lXkWPRXQX92JqD0a+Mr5Rux12o/HzrNilF3YcoA7vPAnzLhhfpvZ7/gJunyErL3jbxbg0IF5xvwV
Tq/kfzodxlYxG45YHSVkY9XbnIXPr+WqXylPnv4uLcnciDdzb5sFwNundGHosXZ8CwYoVioqDedd
sxYyLevTV1jiFZCGspqPcdjUdTzOgfKZARleIa/S26KrFbXRt9lMq5toIneLhQW8FRY75X/0lidd
d+JSB8E2L9IETZpzjbOG0fYNxBbVu756+1sRTyCF5eZ9bj7JlhoWSxeX7ZdlkrLujFKkSGk8JyqG
Bfhifyvpg6at6d7229CXCxK11o9OkHwnhUasAy4J9cwzgj4luKxsoc3mMi72hSWW2ni7XrJca22J
bCyVp3qkEbfn/cSrmixb2BE6pAnMPvZNRYp6QVNxHcQ9ZBXKeu9exN75kOs3rOMXYw7CLn1oD++b
8g6M62CseYPHK8icj62etPa3qyK5sKTtSvM/Oe0L7mFlIXELfSBz+45VR2PwpW0+ojBc+7X8i1Wt
7rUT3AgxzubvYVpUV9atAhm4Zd4L339xcnijWMqObLZ4Mo8dXCqO35rMgwLIIOau9Qpi7OInmDNS
/Dy3XV8zM94FHE4yn25aLF1fp+XiTDyqKgRz7SgV7pnKvjljEo3hEDYhfAgOJqjlAfJ6Njne5MnV
6aD/93ZT2zbmU8SIyDMIpEd39iFYdOOAeVfZr137YU2aF59hfDifOpNQl9D88wLY045wumznduAg
gZE5rEU/TfbRuqENrPqOOSrEyG06HofYZqDEFarwTFWpku2//nvv3/evbqOr/fdcLqpAc+hqndj0
Ot5XJHZqDDQn+GLcqYk1go4H3x2/qHVLwWhw0bIIama88JnD8WljJpV0kvm0peBUdcDRHv+0jJpm
7rYjssTvFZNXe0zdNpSAA6CKDjY8754HjObp0Y3tznO4LEf1r1T29QeNSGLmO5wC9P/ipyDZqFpm
McC8XfPvd2sNPL8aWe2jGzshbrNl3J/yCsMOmMLqVV4VB6yYVh7shJO+BVxh86HHzKfSh6inuYRE
xRieB6rDyxEHoUTCoWJRmgOmzdTArRvoPsf1aTtBhCkNnfaQ5yqnit918pxltte368tkB6Ysx4N/
OM9ZZL1Vivfww8nsEBV+tkKd1vvgCDMofW+m/9lh+XQ+ZT3TVXxMNB1sPDSilq40RsbgAEExvm7r
Zce5irgTNw6Qg6PYNjUmVxsf1kZE7IYtIThbz16YA+GaeeiIEMqXn2zQZOB0t7hJ2voV5c4KGVij
rqD2VTydWkjsF8t51dgGZP3lGbQXOj1JE7DLI1q6XbVY3izlvJe5vlK0DFlH+La8G6Tknq1gbs1T
p3j43hcdO1XyDS6gVLnsIQrkEb24YT501GZb+2ft3VOt2l3vNNWAjKWpyruF9J6XrKCDtJrVa7qP
wpup4Z2+ewW0ieeouxw+1e7n2gwnhhsdMS4MHZSfBK4M/guhKh1hsvljaWJ+eZMQNgU9S/CU/jKo
HXlP5LzAnhvj+IA0TgYVSeB+ERrJRXPiV5K56v4remZrPtKQF9h8PeDLlvZPYiId2SvDDNp+DbSb
isvxFw4Vd9mMt9fVO9OFNXPhyyZ3GdM9q56hDpXDMKRyNJgH89uSCkm01THhhxDNz8OPtt1ZtBac
ero15oWv4JvxyrkJTrL1D6mqL4wJX4iaXWDoQ+Uq15cmCUfEo+lt1iqGtqAQXc3qN+32drfEtVG/
f70SnzDKG4wzVGEhgDJ2WPL1BJmtGj5g0iy9xabKDz5STJ3ugVpdt35me+FDTBsr7klL607vHAwZ
CiZ9w+XXQf5nKgDGSyBPR/x7ZlYHhFXQk3Gneb50WiMt3zrxZxpYCy4Jn32ESl0S30kw9iGgf/5L
yGgQ6gtCSWGDAFlfexS8f6vxieKgvhO0msvEdqYHfR0OcuydP7JsvEgb3ZVoICcXXBItV3yQjHCC
pjcv45Hktwd8s0E38AZgJDQjEVzcFZccEsOWspNwEhCPZ20Z5gv/UIwMRlccfvQdsRoUU6MBbMSj
XBRBRNDX+NbU9B1fgTyZfkksIttzTiF0GMw6up4L/+kKfmZgU+t3s5yQBiuskMMzsH+vClCQ8AIi
KnRi8lFpaaVkI1Wb5sGzK9icdft8TyHDITNUsA0L/6MsGRz5P8IiKyS/EMlY6VuET4t/SGb3bciU
NdbwdqBQyZngDfA3lIY/kph6xFjFO4JqZScarOj3fI+NIEwElFNpmyP5bFBOw+esK/eHRNPpjgRV
AV3utCWS620J6CPNxdNEKJejm3iWrsW9H5B9JzzHNx+ooNApOuV3enCmuOgDZsgcIJeIe6g/1cEJ
P9M3Vc4Ujyw/CSOFmsS6BgPR3h4K2SCJCMwLvFOlsY6T4lfW4bTP4wodDvoMddtIQX8I5B0t2llD
AueP8eJmkuvNMp0AwU4DAyxs3ryQOkmPrxKfUByTg4QdFbHvjoazZwhkBBOyNDAnphndJuDG8mms
lyB5d9wBu13UpmwpEF1tcjLmOgzMNb37uRpa6ijOW/sc7DOW+dQpi8AiMtLSMGVVi/LwYpqV0evb
6/B/p2BpQUWSaod+05kUcKOVOzXMxW99iq3pEZlY/SLxrR122+OnXLQngvxh3POja28SEzJMlQ99
MX3GmbXUwxkMixewjrOddSDWyPIFMkc6KSbWC3Ai2SQChL8lBi+yc/akSPUHnhrlTnQk4VUaHtiX
nBXDKKs88/+56pOs4+sDyPcNbuJBk2eBPq3eELZ36GnR3j21U0MlrRJFOzNhh5kSP3fF9yf8/crj
L8NFGBF+Onjbj0Jrt1hvxz170dLCvwqrJem4M0/UEhBrmOxT7j0TPVAxflMjNJKRqyMxnMhNcLS4
ia2YSOkQE1msbS9S4Yy45IPcMQFjCZvHtx3LT/aNTu1DIQWtcHcypEqeRwr6F779zGieGTAzx7kL
GPtsrd91jJiOOg4tZ1NhSMFBNscld2GHfAma3ok/A0XDqKA2OYZ/zxiNAaa4sNdA0c0NYXEHdSRj
TyHifA8NQzox6Vx6Pd+q9LE64olPsYDrM6y+d0vNcV50FFAsWersAaF5cOylQ1e9YgxGw1EbmkHn
4ghbab2a5pGUZzKZQ/Li6Ukygbx6EnygOanO/MgvnVlLwvfuBKI9NKNTqR8KyoEgticpxFgnWXNm
qy/5eelRiREHnVkQHgci3fb1qkasxrec1OQ8Xzz5TQ23QZfWujnSgI37jUGiIU+KdJh99c3+J853
8b3o80YLB3O2y5RdnCBmXrUFMroR3Un/HBmUliIB78tcYz0Fc8HDPHCdcUe7rGqo4M/acSY87aH2
nqTHQzGgr9fywbfkugHu8P8nnsq4bFPYAwa5ZJuhiQpYjjWB77AIPxEFuRa4QXemruinhPwIU8y2
3iav0hNx1wPnfGpjDZHq+ac7FbbK+1p02den109p/oGQe5xdLDtR6Sqmu2UBxz6+U0+0TMFBARWR
IkYya4E/BNRizh7u+fp3nHaTGda3monVv0XgnIEFLpjrC/1FAuNXHzgKZDDEvq92IEzzX6yonbEr
vbQRe+NoaVK3yr9rHCNrGXHbhcM3Gi4KeuA9SBnNtBnag0tYJa8hUZW9Y7o7T36a29QeWLLgme2E
oX6OdfW39BfrD/0iVQkYVvrmfaghEQq2ItbefFNyWCnk6ImEwQeZxE4g6aHVAn+LF0vOsVBkwU3d
KhFPyHmSbpmgkl13td+NHpciwaVjLjnIrarKvVjE4CpTsG+VoZ2VP3nj4A2vjM6yewbFei5pte1T
qa6DOLftvJevxNinwJi7ncUECZ5M4tvRLdtllq0nxuPsfjB2YrxTiinKA8QJeiCv+XOSCf456eKx
ngMQfVJNKc1TN3Ly74nYsS/10AE+SBanlrqkAd0BHrzN2pnR30g7NEoKP0ck0q8jMSViHQQrS7uO
FHm/YySir3z6nSy4xhurxx7B5g2LVh1ISt2tN6WlKEaKiggk6tCiX/pTLmfDasKd7i4WMnJA308v
E9NI2IoPdJJ8aZzmHAjqmS/fl9TAVp/Dl/7IMPGd0ZqNtt4n3a7vT7gWYuiKDznl18fMk4myerEK
zKA26fYMsedc4jTiV2dEeEM0f+lYt5PozGZaNRdFeIDC42HqGWsgBDRiHkaUtFQQGG3wufaYI+vX
qmBHGYNTl/epHac3G/I3VWAq1VskVmzz3fLxI1YQhkrcpW4Irh3CItCNd6BOQ9HzBcze7G7jxcx1
h6Cqbgm313Cm2mvz0BHu4qxQs37FexFsFR1nlkiRUnOtpAmK6X1nZpU/Mbh/Ov5epA9kmi9STbVE
7L8gYnappISYFpKPWI2ML4hvYQshIWag/yi7jJeQqc97irQPxQuXfVF2tPZ09UaUnF0AoMg3Vl1J
bppmBGZD8+Ir7bIjetZyHzWx3dJsFP01d37bxaN1hiHOD4JCtI+oDDb2tbVME5eK59gLvGBeynxe
ZZpEGubErTFJCgHsKHMCeC9EULG3jJq1H4giTsG3yLOGnL6TcQ5jR8lI+3nAs1bsh/seVeRJa8Qr
Ob6nVn3IFA//lPCkdTA06/va3NNbQRFzWSDbnrtHIYt0QSqK2gXOgrUbwcW3uHEW3fSdfS60/E2x
kghVIbAcOtIMYiPsvchVEDd3i9WV3nll1gr1B4hRUUFx0c3hmckmAlEM40jnWSf0oY6gaC5+EwD5
E/VLi3wNYwAhv3bqi/aVqDrcmGpREFJU6xpzxKOyF8q+Flqt29zcTyoyTF+812e84lYkRxDrHB4p
F45dxXAULTtQHkCVPEhHjX0ZonaUiZjkLfTto3YmkSAYyZfDVddgBYzhTL+DwaljfstErOjwzRMf
nmifDZhDeRfPT74vorTs4Z1S9VkWGJXf1hxe77FkW1LE6//8KjS5jgBYHN1fYysGwmQN701/Y/Rs
aob8GvMdkudZ2bV9k0fSUeN1T/Lb+XBSoB7mxmeGzr52670+gxfLqOvCFemqankrAWsVxjaiQSbV
TVAB0t2zXI3JNUrUCDfRQXdK9krE3hb/1qwFM5ZSBVxXDq61i1oIYNoRLfxcTlU1ZNQ22FhUuclr
gZxqcY6AucXlj6EHvd5pAKeN3iAQjtwbm3+8dUJpNknKupSyjCLrXxVyc8NLTif5BBjAzDPrz+YO
mYCUcHrjMF74LwxASsPJvORc903VotWSwGdGGrSbAO8xlZondvtkXANB1Il8hXlcB+TVO516jiRq
M4o/r5fFvz681Q7CfpEsuPMrjU3U31Obuck7fYYpDAAZLhXg7Th1jZH1TsqGrIdc+2izI6F4L0An
wmBbaeAfh5uzCP5yn+2wFpmIdXOILJqx1etpZqDrd3VkKRyYmHPZXQF6jgzi6FIeV+3trdGEc1cF
+q2MNCFAZTJEtMp42BQXvLKM7ocAkuP3gqF9EsWH3U4vXQqKwrBy2Rz8NdvoRdaJRCydQmLMJB2e
29UdiuLMsSjFCplCL0PI8EGB6fReVRmXJ+TV54yd5NbytjBHLffarP6QN3ZOMNYLVnSC6y7BCP7E
KSLx1F8LoRNjwv8oZzKfK22/X9IQSJLPU4dnsLn5++3f2U2PablvaZ9sGZhto5sD8ATBhO3qmopc
R9bqB2yZZKmesySTHRcg/uFlg8uM8subctQvPcg13cggWEY+mY5BRbnjsgAdW9wq2UCuDlTtLBqg
hmbdCd0L3TjPUcGUue4KmcIU2ISFv+D0lSvexa1Imio9AdJDsL+WtoNoE3RCNFgOpSCVAoNMIhQ0
NAzDyslKUoCELzpibGICX1lEFaGApb0b+UD4oD/4QpygzA8XCA4nPbTcT4VGpEhDRqHN+bbw/J9n
AAHHTCYMfwKVfJTcZ30we0lrlcvyG3nsire9FHDWtvgAAMfMrfuADCUxLe/ZGhCiFJSv16B/IFvY
GKp9DiGW8LZfy4UvRw+RUgMvrKJ8or6w6xAKovlllKKbJgrSBnHtxjrHdBQosXYK6qJN69a/WraF
jSbZRggMEmjaBBsr5u2vK2TZmakK0G3MCRlo0zdQccdH+6noj8oxJHbMluJm5SlUxxEPKhi4bS6h
AQuwS9j8zhkNjzonBrEs5JRpqBb4Db1nnuiflJV6jbFwJnjN/oIb9+D8xcnxKr7w/00HbKiKfste
HhSH7tjggtn1vu1LGFhZmD2hQc5tUFs7XC8gxD3mbZFUA3eryZU2rBUn01XAp6muvvruf7VykrT5
iMhLuF4BRwhTg4UQnMJj2FBBShqxa3rrMUi+rqBbBBh8Evg6GW/kBIoqqURVeRTIdLPSG2IV4Z5d
yTNTbUU4tZPHQGgVWQJZv0AY2NkMoA6KdaBKqG4FnkcDDlH1Cri4SQmbRLA5Zl7uW50CM48A2BEr
GvDuVkMVjS4CxI/0cKeb3obo6o1LqBI5gIYBpiXVvhG9hKV5DquTqUveKeP0gfXx/x7bhGgYOoPw
Tt3LgGBfY9pRtkuG7PBp+k8SpCXG+zxId6fZOjhc5SQyieknDjnPrzTlMSC5Oksy6G5toob87xx/
+20iiYAUC01r4aVi76GHcPVdk+tqhkQurnxnfQUrdZX0bPhnyIdAdxdouEkS6A1sqd9vBQeZOu94
miQxD6rdV5N5A7HHRCJTHvYL06o8F7MtUdLpltZOTzK2gFW0QjMhkiSaDmv/WHUZZBp4s8CsQMhC
wAVLZjNxfJ851VvKp2VR74O8R+jsibbYJ2ULXtA+nlXWvGudVGMBUccrxyyEUw61lp9KoslwR7+3
6HMkSCWQHYS8pVyyWTBh+CtRiPVemS/OtB62FsXevD9Al9aa+8frd8LDSIIdiqc1dru2ZClNxxZV
o27M4nE3jLiPOr0xuF0+GJLbWNfkCwAEND3rnc4DmrgxaZwGXsshDRxTfjH8Lwiw/mw71FLxdOSt
tcF82Fgpd8t0jotAFwNuDtdllTlZPsMbwws/rBa63zSRFKAIclZWKQQzKOMWZ2sFVxUdoYpJ966A
rOZRnozkRVG9T39XDlPhIz/E6ZDsNusPShY3y2iYQUMZmmMyVoVztC4nR9HMxe3KAh2EiPZVAnSr
+c8T/JzgaNkaGtwnP7jGsVD7p+o/8y1I1yV8JrdjgOaOGDkCTDky8EZmAhALkO8ZGwSmx3TQhivt
vEX3mBqWX6USNvsjADH7NFCuhQFfd6csHvousZrVGe5mLuCSyNsxbOUKQzk3pFjQUgcfZKOnGkyu
ymdoWhDGPNNV6uRK+WPDNbqbc1n45jcL0gM18SzagAssyG1ZvgPQfGTTTC9hbR6yTlV/hzb9XkYS
VH4oql9yTfDa7gcOaY8atT4j5DcK/khy7E892lC+jVmtHUrVqU8FcSPGRxPuy6Q0lqfGXYVvZCQk
gf5KMwsKN6FUGjWol0QCGZOv9eK5OGLlneLmtFhrK+ho7GGt5bq/D5YCZk4a4zcVVGrfR4Che817
hbXWFK2ntuW6L/cu84skHfSPJTo9gMYGj+XWrvBUm+rU8Azq0B9TclLC/taR/+JNFAc0SUdxEdlQ
/iYtKswbMiPaRJhGpO1WjPC3Y6n3E34MEAO9QEs5w0PqSpXXyLKRko9Tx7h99+WCgK/Y2uOhjYgl
AQ7qN/68h+PowUr+HDKQ7wMAdXzsGRcqh72qSdPuj20dfnF72KFbZJDuJMnzwiZxmSHYRz/PafQL
36fmrjh2UP05HUs8Q8ue/Z8zRQOUJ/73xf5cWEYliqe37tqY1fvaBb2Nv/1V894nXlpC1yHCe2Pa
GrkBvOJ3Exw/hIMxByZ9+tFZIQ3EETqpXws9wo6k28KnCKJHTfHrthDHhmsKDnMvbVNKU/Qc4mmH
Zz1XlcDBkuLpKTwJrhlUZn7hRsgQKdQT7zT1XKY+T9xf6zDs9QI69eOiYuELS46pAxn3MjGTbCQ8
B2CkHCUgIPt9VZB7q3AuGCVFxDblLYH4BPl+0CQ4IixaNZN8FHk402w83G34KuuIsYolAJyZ24o3
e7yJkeuS+C8xF4VqRqEgOmzRG4D0SUyyO0GykKhb2g+uKxBru14Hz1M7N940h1jqnjqbupkbLELT
R4UyXsNXFAXiXrmNLEfX8PBZBjPebsV7ED8ZBYgeMK5SEuc3uUibKwLQoCSiBK8rhYmuSwdd86+x
/TKFWMaqOBPsb/Nv5KPbj7JBwCTvc9ilGOZepxpvF/nTcDiFuqPDHRigW6AKZMxk+ww8i9e2f74v
PbftzWHoFATpORrCVmyt7arykJx5hET7GE5cL6FfdbdhWBkHSUsu3xwSdbdtNz4h1CwisrXz88Nr
KtfyKAoabs2iCkYdU+3rvFsg66mbxDW4dExoEDzLDOOkSV6OHsfQbJcIBpxsmmRSaw2bofjICQuJ
S1kRetGMnCXr1leMCgrPpfPBEpnExxfNj2weAU++id7ADDldphcvV2huO0/hNwTJnVBijbarbFlX
xttOGpOPE5VxJP1gGXUkzPKDtyGqAqOE48QCX6FM8FQ7leo1Bh5ICnDYKzUKanBQq67C8sS3KTBL
kAPSb2kEvOPkosp3BaVrenSu+4oII72exJ6Vgmajp/DzUE55Ia34hd+WGj9G+R7ziaHwHNH9A0kL
V7NCBIU0WUrpQ7ANITFfH3Z4UscFrx+WnF99DaurMTmUBHdV7lEpQ2pEXzW67Cnjienl9eDwF7/6
9Ce6Vd9dOhtCsNb92+v/o/jiDTM8xWqX6RqzjJnSCRq5FsLnwoFhxo5MeespK5zhvPHuK2Fzj0V2
iwpAzlqadUQxTfgFQi8P1S2T3dVJa5nF5yqGH9WiWzKGeMyBHrml3HkJNZnoX5eVCUCBrLWayaki
2X+aAhfFVwMxCcYvqMFbr7MfXv//1SPCh0aQEokrCpbN4zx7Zk7qXEjKchTT6+SjyrYTtQLaAFcb
/gj48paZohJ3F95Ktxws4ZAzVqjQ5Wbzy46TyoQrDKIPCGV9QlsiRbiBiJR0R9eG6QmI3VZ/Mb2x
hpYDGgy0DTedT1f/e0hJmxs08X5NEv2fBSzTkaUZLdZpuC54vwoi+LeBjPr0zq8ADaDJzqxDoUkR
nTeYt/sJM/KTfA0MB2bhTQ7+rgn0pS1hDoO3abVgBC7roMmvhR6LajGw9rbUBvty7HG1tWcUYnRV
uxi2T2xAMMlis67bqnEcHPG40r31HLBsH7wGOfxBEmwHnBB/UtBfvJyRioPQn4TnGzKsLwD/Stb4
c9dqbHBXz8w4NvRGG2DKCFlngL3Tuo9cb08PUqURVmhBXq25SpME+7yZ900lfFxP+z+T9gC2jwgX
9KV6NR0xSlnvzBjsG6VAE1Nb7vrmNEdQ9zb6QA/EA/NG/uOQIvOiPw17xlYRRcMv7XVia0Qk0hu3
rNSFmzAqY/K0DxYOGAN4L4leB9kpUQQEq6F4cDnTmBvY2OEOOnzvAf5TX5I0HGqVb7sycMbsOkKE
JER0f7x50PEu+HbSRhnJ2BZv3MjD31J19nlWss5muLgtCEwn6NGuToBeGGDe7SelMRm+qgEVaOOF
2JWa/lWJVkpjupQPWUJby9oeCP43Ef8fY5qAEdOsXNzDbYlEww3ajV1E5U7GU9oHua7im9oplxPe
nYIZ1Q5BbrG5SbfiAJWaB/XtHM5ctUy2C1TlFJDX58ELCpi83WjSBM0A+OW/HROt1sAa25Ss4gNm
DeNJxNIsbuO0O1LgiWs9JHxwbDgsdrNYgawiyI07siBNJAO/CnOu34EakVMIIzVYr2ftiX7oKvJq
EzZMehd/ILwMXCl+mf4W1VBRt8pzAA53Ad9KVSql5fMQ9Wuu9adqeZYFPZbKo9fvsAN5lypVB9YF
+ovgI8J0bLHgcnGdDWLD+JChv9k1gdv5/Oeo8QUIIou/fnNdBYecpJNlt2HvrY9n5CAk+JzveK0N
9m8A5twyti6XBmB1G/KLf1davXCBrJIqnQ8YcYmu95iFfXbvp64REEvoCP2erXRkxm3Qk9s8gBIa
xUPsCxI8yYn8OzvSNiprRHp6EkybRnurAc0k+81GvKPm4C30tpVNuNBwhnN6BG4sW+Dv7SN+c0Ii
/09++zTTR7zFpvbbKdS6ODXKQZ1YxOW9FwN8H/Cuxee+yGiBoup1zS3jm78MFnzvRxw4I6A3+x9b
vil3abqadB2eKVLidGcfS0gT4nz3pm2ua4BL2OpvMWDG3jWHEH6si24r0rHe6CagubDiSZaqNdew
ljIq+2xsyJBo4j2CYAV6anBh+O59qGHDnYzvuZAiayzbuTI7PTh/3+Jgw9J9NL407TQXB7GhS5dY
Rb9uqE65fAP40wQxtB9hnHhTLUXn01ZUOldnLyMO9LwtY+2zgghxOjPf2hu1uciy+ZcBDaJehEP+
fzUOstuL25BPryG7CSrvuZUTBqo9XvAHV5U7k5pGMXoRGGc2pBkpiltv66IBRGQw5lhHuH17UAfh
0+ciAIlIIg24tPTcvIT9U2OSrwxHsORlgM+P15/qPcc1c8isTXSwYeCqScMQ7k2e1VvU1fE8lmnQ
6Lp4iUu+PnBYoDfijVvYGevz19LSLBIY0MettPHk2T0jgBX4CIA0UfHSu+YW1prtOvpyWpuae/A1
oTlPAoZs7uaEYvqssMuz4DAwxVbJ4KsS4EBqR/81HzrvmhhL0nZ9M4mQBGL0FiwebAvPxK+LYYEz
wimJ86inv9Y9Q/c5aosUmp5TlrzBbEl5t8HVDaZdaXgE0Y9OddLi1JyBn6iHUTFVHHkRJOoQ9VUZ
N5VewFOjPDydkmETC2Kgtw/NRi5+vt6SIN2eCEj4czlujR4nXD7or29e261SWTz6B/3T/gZm/v12
WV+yjz7G7Y6RSVzfDjfgbj5GmiE3sivZSdJ0HCCzhCsq/Dxjftw615zsMF4A//0FvB3RGRamaB9D
UYm2xQUMvrU5WMIYP+Hoq4uNJg/wrDr4ZLmepnlQQA5ctbfmZgZ7cFTm4FFHrIXhnopETMCouVby
Ef6hH6uSoc3uZc9tEN/YmpFM7hqF3iQr9CyLRpHx4LyKPkgERgXAczbBS+kIwn4l4fSHYlAV6q6d
oDqAOx+8erQfnV6nJ0aCgpJWPUyAJZG4QBkqr5lmndajIREdtrVPzl/5oQ94F20VlzKAwgS0Vjml
Kah4KWGpAsYca8Pys18+U/gLUZsq32DKXDOHszBkr+37tI/lFR23EW2EhmmMnExistlNb3KlnY3j
QLJ9y/g+JS7PhenSKkgluvqLRJt1jng7P4bX14KFd529Fb2va+NCOrsbfqN8inb7ephxsFEnpyER
pBxL2psD8A8moB+8oimYFLhHM3kMBasRQw9AU8CDhoJWLNGRfMGFw7sVieutpu7X1sB7+zxiMXJN
dEM8/ElIBPG5aX5/8d6mHFj1a51t4/gHyMvknajFhV+xzJsvAMFSWzzEnkIXi49MezUhvX5ASccD
iLYaUiWh6EbYVST7mxt5IFx0nSXHUx8MCSWthzTuJicW4uiWd/y92XTol66TzJAiNcqyw4SpPa3x
B6fT/M/jvghFP1vAF82yZHcdcGKXIWDJ2DnOMRgwq8zPpStUGpCqhy/LNN2fUYwtvHxtDrv0ovXc
PvHjbU2HQWhS+VcD4t+2QuquvAYWhnX96aftrl2LZtN/dCq2NtIc1ffXPerscZ79uPp+KhMRNLV9
KIuVtL0M878hM5umzPWiirArKabcXONNJrvpFKE0BgaifLFp5LPprxUXhOd4cs7JAnK3GzJFZASr
EcgLiXiNfIT19R1Vn9jq3FKTQIIEmJ/4dNqA3AFJ8R1oAFl8YvvL3hYXDl+/SMDtcf21fpIf4y1c
XBZaDdjazmzMSOmmGY8KgM61UPLI+Yoerbl7yoNLBxIv0zPadvlCnRpOlNE8RRLyyylE/sAn/b+/
R7gGQQZTDGYCmrV+4sp76R8z3CpC+l807R7L99PHmAzNqRXUdY18sZ3Zy/yTw6vvnk2Re5AdJttd
wj3jKjiKu5tgJwBV1lrlvCEJpgPKqGi6m/XRQTmOr2aTRf/0NqTWXrRRcvm5zCMUqTVBQxLpJDh0
LcKOZWF7dGLNlYeo/ZWfFkdK0MEBzHiBrfMndweNrnuk97q+W/P/KG2OEyroBR5GQbCw0M0AeD0t
c9JrjEx5dT/3dmlckpEKB8FocfCCT+pIb6i/16MKorim+iN5JYzdHkdFQOVSy1yTJYLH30/0NoOS
X+506zaG0zUVYzcr4ecAP5jPtW/mS2Tl162Q6bnXPEwX1w3NPbsnRYr7si1Wtk97spKQ7rf/z7Jm
G1pW2lllXeifKliMnjOpCG2p1f8GNHI/d/pwDraAwiO5NujVPxiYxK3owJnau7LUuK/1nPyE+u30
tQBLXpsCV9TfJFFLsR1LAvntdu0vKeac+QK2JYxnqmIPfFrQflCrO38WojLjMIUcDnibYsjr3hP5
vS/8mONtvQLHj886/S9wylFIv8zSHWnHItAsCJu56nHDV1eu7mfdQ7QbNpMzXCAfS255AMGX66Um
B2mUvYMCPh3yZF7ltUVsl9ZBPXp+zAGhJTdXRe3MIT1m7HDJPkw/ZnlmHQk5H4Y/Et9wquLO5N3R
BBEuPwMljEq55RaELO6iQgVunZuE2M+h9pYTwUxstUgn6w9NJa+Mp2IimHkumiMs2KpN+aScYaUm
AGnIH5llxLcb2WNCnDy0mFU+MicXgU/JKOn1nNUyttYV4mMZvFh/lNe5fg6nOzDlSMCMqWuLKT4p
QQIelW2C2eqr3lIATQgO+qsiSMznw8IVABd+JEX3QiZnFGGoABo5vlKGPtfrfW7hpBgATjO/ORcB
m0yhA9n/OEAqWRmx2kdQj/zBJGG0uZtVSype9b9nSOhuEyqzUIGH3mBWYEhJGCfqz/3dGFEIusa7
6Pq+ZSjQwNdSPd+uBmoYwhSewfslg2RULGlW6G8T43lr8D/1gCm9TFLM1toD0E7VBZvr7i1voqXe
lL7/BK+cwhn8FNnUIlG6TVW7lZXUpvWl6FmR9uKojHnEIihp4eh4UviGBIHhu2tvJeOviupy2e2H
z5CJReTrBRJ19o/o/PK4wh3Ot8hr26gQTOhdHnhUA+XuSj6EkdIyrQMThvusVU29GgK2yvH4OUZv
QHlfHaoAGn0CIv98SE2xOvXyzF/wdK6NGtW91pRxpyDG313NEoKWXL/kD/AF7Q2mcrasu40gXYkH
smZaJIK2OAa85KPpaWGY9dpDktnwNpzc/Vhrg/CoclfTdKbLdnjD05UbQlvZft314WOx3MkCBYGX
Q0YfRpWfYC0IpFcO3Fn7LBTktfOKqLiqb9m5mqWS0BKM+6h2gBK0t4Lb0HEyANPvgeJ6fmITKbpI
JTSv3GwhSVfmUxSWJSbltkD6or+oZGqke1SWwODgHc3W5vh8X6DGxF415NX5Jwg3QKiOjILnDQQ2
HQOQh6Njg6yt50I6noPRvpzf9NkpWkxbHzADYmyZLtxyw/Ip/n/hE/fpT9OIIqLFs7T/zoMcrozM
RXyTeeFLFzvYk5jYGSsuO/wju1F1SkL+XJk7GK7lzEx261yk74YidNFfN5EdsIHHsO6Vq7Ka8XOS
puyn2hRZndvPn9/iDiqSzqcI7VTW3/vIqrIHfUu+5AtN/+tjS9rKGgDtYj2qaDrELCSyF6v5nFYE
XMUNMwj3VCp92eXPV+RZyFF4RGtYeuZLNtBguyXQglY/bu0v9wBmWHub+4N04Gh8cNKExCZqVbc+
IuK54frSbyUp9CPIPJs3a34wmFuubAWCZapwaADBx6Zb/k6CmblumNUfSlZYa3D9IoeIFsVlNxrw
zrSDKH4r+wrfFj/HVPjA7d9vCcOj8NHQBUA7k9mMBvtVPViRH+FkrSepz0CG0a370NUbQE3O4yJ8
n44ttspz+jv3tNA+LDgdB2pLH5qzAiQ7XQU2Q11byPsIifd81NCoHeh06GhqFigakYSpGWULefRl
xPI5/de7sdE/kmqn1qBl1nHmnkZc3EiyENEwSS2EQu7FiEJ2o3zi0NQvsW5ByfSGM7dOP8xr2xmj
TyKu/m1oTwksiJBrxyTMlbSHUu7MrGkaGYjcEaLhf6nB+usPrwiw5XLVNAfmsORVsjRbQuGaJ2Q8
lwB4WxI6eNIrc3IYIvSG1j2ZzYk5CkNjXZ4Bcu9MzZpbG7oQ/RfsZJ2JfLokWPH/XEMbhm2F3lHj
p4qkAg/IkH9Tpvlyr7Lu2/a/EW0l5IUeqj098YpyUwAkS59cEORxvZwkCyCCqBmuEKB8pYsHmGqD
gMhgZ+ZE7cJR0Hh8kzNr5KxpJ41vw2qN3L3k/JGAfSHJVLkpF11ZJoXXlO15oNkzLIdqfz2mytO7
NWCyXsmVfpvBlcQXzY9DEDh5+D5aL5VcAKFcEJF677/3NVc/jNrBJjWxq1cy2OM0hMZJ4ATHUtMJ
VtobXeQLtWEUVjdLfb9KR9C+rdLKHitCkOUQBV1+JJSYH1k6GWPw2recKQ/5aLXZqHkOjw4VxpAz
yTe+JRCcv/a2zxmdqgbTwX+uPaCCosS/FeYgOW4XrEfiWdZNem/RJhXs82FR6qB+F58Jg0fucFBQ
Sh8xJ9q5y39zit8dgd6/wY01Hwi07oobpQ1NqYJCnjiRCvJaG9bdCcp87Mu4nn0TOaznFU+X98os
DrdGcoJZuQMowiM9ZV/+tvrzrScBmrXdE+HovW6oV1ib1HL6ZwBl2565JyxEWCr6sFvK9g7ipRS4
UZMXYHE3gpkfasCVX9QoN4CT1BA7nud/FAlwnVIJ/0HySER4nqG0C+i06QFarvZmWvRwUVyN1Yig
PpTRqAEzVEIDyb0yP4wIT0oenWsPXRANpMQW/H9y87KXL/FmNhBABgiGlA1gN4TwPEdBnHhkbAZY
MOQ2ABzXkuWE5i0IKsnFFj1tbABTRRoVI44S0JPzn97Gzwqv/v6qMo/JiLzG9FfqN9+QPUwro9EV
W431uPwKtlWHRu90ef/aUyemLmy+KarAB7fPo1rFc63Fu8KrJo8Txae23nr0rkWe0KWbkl3n2RA7
5B8xx4VsRVKEuGFeMWfr5TIj6EsZ6LiuL1QflqCk2cRBy/Tl3E02t3gMAKwBaO9YRGt5UiUow6j7
ItO3fzm7bhqydGMxwIMNo3WZaShJEQAhtxUI2gY1fOX08oNVYbQLMEj9mLLUA80KmZXsBS49pMng
/pbTusxhR0ZJ39rJOLE6L267ksqT17icrp96U7KVPu9+ZVGdlZlZC64dD9p/nz+esR84Dqsereqk
8jzocdvvzqW0Yk9w2NdvY4qV4r8glk9gv9M5BOvJfHX5AWaOU1+5wb4bRQgRrO+ojJDkq4r5ibXG
W9OJWwP0tASeAini77h9Sx3BdJ6EIhozaYM2NMAlN8j91u4k4wa2LlfDe9RGzmnE4ja6qNdBwy5Z
kz9qX2ZUI2iUA5j/wZ0qyF86oD2d13AutYToPVbyG4ZFBEEmE0DCNvc3PJuBDk0KbpHs1gq8LQhM
aaIxGKmpEaqW/gYZdPhGU+3rOJjQL8Nzah+cJ1nsCMvM09ByrEUYZyRZgoQtTmZfKQ3UR/tYpJ2d
0vATiHZgZ0StwDXvTUJtrePXDwEz5uvbJXKM9x6gxxZyY/ME7pqbThKoogmy0HNtZHKnYchL/iuA
ADrgGGW5ScOzmHCPmeWTVDp4a3JTGN8lJqz/cCkgTdHccScXEiFws9eVtLSsifbMDThg7pOovgLJ
exs58QdmeuyQF/ssmNembqv+Oes/EtDNZVhBT5GhwUPLqNmzdB9+qmD1OKc5iVcupL3/2nIknwRE
g1CDaFTtrt6WuE7ql1A1vyKKyLkkkNdCI5GhVOs31uapSFaxg+U11UhDnHZQ1453qkgf80kpbc6v
aTJTlxFWhqdfI2k3XwzzsJyL2IhAr9Ijtg2GUZaV+ewfBZVsf3gVbJj/tiBC6JQuxBSeyuAuV101
xh+dU+/JbumEPCapuCAsO0WJvi1k4CQPcA5SPrUKll2T7jwW0zjMQ07iyf6/FwKk+55uv2yv9uVN
a9dzz89T9Kulj711Lw1rZ/IvLYGiwqVB1gmK5h1cLSfyG0eA5Zy8S49lLW87Y/L+s+kFHZgF7ROD
uHM3NLG1zU/aZPONWjn9XcTfIrtc9F92/+Oozq3bIQoZxnZ5Zu1H7hMWsAb9PDWCsuMksUk3fVnP
VmccG9D0mNiaWNRrAX8sNGgu9Q2QMwqprq8UZY8UaU4gdvYeSCPXFOsQlgfxZXRdLS2NEkv1CyRE
+DCGB1Wiqu7VZvPkVRpPlG68FJJHSJLdk0Wdprw4vWvwD7j3lC/B21Cyy7JxPm5hpc4ysXYBzVmN
iBSuXud/GqnuqWVrzt73hjW3chM+fvXPVlc7DEpaMeC21h63/zE7njOC1/WECRrydOPsa9e2rAn3
97hRgUeG/0wFAMKlwwPnn18qmBaSOEaH/YgXMrrXAl/WQ9Q82CZwqeLpAZTodzjveNT1S6A0ppx5
ZAVpdU6cfwXO9lilTu3hXrh87IyqgeI83sJCG2jSTEY4FuCaV4n8D/p+DTQdi0O0L/qutdwasnAX
iwRS0fETO3Q1k8S0N2S11Pg0+9yNcur0POth7nk+kVcb2YcVq3gZzCE+VrcwAN+w9Pzlp/+Gjc9Q
MPe/31vmY7ITTX4Z0ZsbMpPk6nziYFpgHA50LdlbUYsskU4VyM/IoepkKIKA3N2niIeliSr/JsX+
vuUT3DQ8k5eZGVAxcm/rPwuJ9J1Fr1Rzhw/kzOC1404sc07eFGgSrsHlhXAGSn6fAgV9pHEVQk4H
HSnXumf6i3G3szglgJqGjGFE8sQLDCHQaHQaAb7Q91XNZyhoobU9gC3db5hpT5jZA3pE2O1oQON+
omefQqvNaa6+DpzJEIbksNBMfksA6xjd2hnGsWvFllyoEAtK/4R+Bp4mO9855NcSxxXRaHx2oz3j
ne8yYP+O7DbPgxcD+BQlr+Qw+522nJBemeC2iFHYgfaJ7FKKh4/BuzR11PC7hek5o5lY6l9DZCeV
5H1bqwwQ7MAcR414iWLdUJ8OHkuZS2qr0awPkiND6DMmRhkTmEQdWkSWg29NoBXNxbYg6j53cfcr
vxhgEaZ9KDa1lt6rwiQBycLurQcgu5+DH4NM4Sz1F2WPweVV+j87FRMV/zCXTGp/+0Gpdvz5aaOX
muGeXWWjpzzLAmABnJ/oaooDS5Ed2NNjmF6na50WEcvHgyzPxLP91pI4Eiy9v8S4Tb2H/WUJ5UaS
8mWXIUE/IlcZ0xBZhULE3INIvGQvPzNeeeIxsdO3q8X7FuA8w9jkZiG6kM0DbCqL8r+JMyGZkm/d
I6o+7pj8sCmxv64ErdGpSP0As8eldC15fdsVn1BFKYIhh42RdE5Q6Iuv2YKegptrkfY1t9CNDG1B
mdxIh3shRjGbpgikRQcO2eU6MjIIdBulu976qh9h50vP58/CtqeiGL3t+43BoPIwmzUFw4oHIzKP
lCNWwd0LUJ5NiHSosQxF9cR8SRGB88VP7IEt2FuOiSEqevhKxvQG1s/MiuOHcflWQI2lEMqCfm/1
yY7h7dTxuM3uVgi0wfrkOTH014i+/+rOzRRFcuEGOLFTxrZ49+zmeag4Up9ofgWRaML4BK9WBcJu
0PuXa6wXVdb2JAv1+6fL+e+f4KZnwS3sl+9GJ9XNhOO2tNCk9ExVZvWQmbX4miSQrB7RUwDNT2oE
w6dDZoY6b/ErUdzTwnXi78IffndSXsrbQtkT+zpUpQW51hpyNHk7TmhE5aMKlAIBGIGI6M2qmSbZ
1wjXPkfgNlayY4XmQawn0z5aZCSzgJLkZFbD+rZwEVg4X/SUky7IjJv8hnyWH4qixB0eAWBm3ZnX
tKKEbVBj+lq6G2faQ8VmgvfwBDOssmX5gbHaO8bzExjjFVhaqSnVLQlEZIJAjZYRIFYv1kBVKOBm
fJWxMmYrqIzrAU1CEX8OdN7nOY3YoZBpWVIKg86Ydn8hzEf+Ux9ewwLmx709jf2VFZZ6UX/q4gL5
26bPseb/jheG/JJ2IMccK3kJrwVzxzWVfxJdFO8jyF1/l2Jm0TY9XO5z9cFIf9S5d+rNGNs8OGJ6
bMb32SkPUAmLMM9g2wQDMGbmX2VXcclUdOrNUPP/NT71+Hr5nHVPwftp2LRmt6nPDq7l8VBTYDec
gNkPhSoxJ2+FyYnvXZXd6oFekk/T7AarmzzAyP5U3rJ2uZg4ZRde40gT69CgKAxld+mG0t7RxW6v
QKg0C0p3Jmap9Q71ddWxP6smfIdD2FGGVAuCj2llM0XBIVRoPL31xiNEinqVxlAIhmADTbUVe9Tg
gvg9cSp3u6eNmsQ8bY2PVNXK2B5ub2uSCS65AA7wCoqVW1Le/PAv53PweK238c70qCedR6KEAsFK
qf6CrJgtY3c1EVuU7BEp2+cw+VszwyBXW02RDRiO0CKbcYVhEDuCB+50twse1rpja1QVHC4pj0f9
phdd7ne5YuYor8kxxuHxlbTdNnd/09e6OoskYORXgtTGnS63DeloqbEKi4YXRXHd0PruRClUVjn4
3ML7/biEnYWDDhol8wUrIWjELec5ylxvYRVKvilutlfXiwDCfAng7WAnTHXUp0TVyb9bOA0tCs96
Xbzqk1T75fFgnaMUp3tYrIVmZDus3Y+JsJ9eehDyfQitSAfJfEOcAqr5gqaerMwz06ICWZS8RxO4
n9ET9LH+USygLhxFXwLYs5o8lCADOjjBa6QmOXIjlgVZql80LJFQ2SZuOHC8YqICIL57ZDaM7axs
xgZbRTTAJEyWUvIXfse2aQ6ZsLzZ2tZwD0LtRrp/YNYS49niN9BhDbWDtsoxukd1gXRTa3+k/YPH
JHA65hQUIFyd5CPWHGe4XxDmWshibJjrF1KJa249CWF/S5QtBCMauwocIRHaG7zU4rZHGT5Fz7Y9
+Kq5Z9y3heg/sZqp+WzL3ZxeL7FfO0VktZ7QSUBgiYdKko/wHTF+lHgzdqGLIeEvDUHXBfiNDMCV
hohf5gHnl/LJDm0UfpcCkhgYZwpUX75sdFCfjOuxYOU/ABflZfOCewVIbRqellhoioWsIaZ+lF7w
MJf5qXO4evbZAq0CklegP9H0ii+x6V0vrDJEprRIRIcy0xIMNG9C1KTrC+KIbxFrsjkgGZDxewU3
vFC0J1PJ/06e4/Gvs8q2oby+xkcT5b0H6J6sQaaEb65Cm6HBIpx4mwg7+EFpKRZdfW46cFV2Ti3k
194a/shmMYoR2aLaXd3iIqibdxnbOP7xPGmNTMY5Bhaopczg33+Xx8H7K6hSAXsA8uWzTrNYAbo7
G9q80C6m/uSSJzOxLQ/IpNINGYC9IBYxw46Tb/06WZMYPcP8OqetvtqOfpetwto/1/GMnQicd9OR
hLXglzWjI4d5KIqKWDMnr3AAJ4W12n+Gc3q5KbqDu077ycugiioRwYDAuwfGGgE3U5pfyVAy1kTf
2hlVR4v4sLew30MY29acrtdRE7ciAwY8yZpgYznD+E2fXMHB0iK2OY9Aawk5DLKgXgBpwZBW+Or0
brC7F36p+rqZDQ981fk0QB8avZMUrcPtGEdjqS3Kth1Epu2R+CSMfaudX1qrqFgI1TJ3Ina0ChnX
VnXUO9jQ/9Sv/RfETqocrXIGU2Wsl4F6FppdD9WKareeWG//1x6nUCL+2fQ+InQHDW7yzMWsqRAc
OgiQyzJdbRNZh64RuxzMJ75w/jVb4S55d3dgowA7AETq2NqmBZcYgdvgramQ+eERcSkdNLCce+IW
3/1yqAa4jfe0FwCaBz7wZ5Hll0v4O/oD9ck9Kjk5w8We/UT+lsGO20KQw8+/1wB6teey3dmc9Elo
yZ/fMNUy8Zg2oYq+mTQ9s7pDElhykhhV8+DWqCa6duccueJv0vQD63PG40S7wp0+sh31Z5GG1x8E
IQupPymtbLhZYpY4WCwMluwKqJjVwf7PV7siau3L+quQ73E73SstV1iQ1TkgL6ZELK4VQS/WFk6c
DwZHS2/04amCk2oC3C8/upBz8pnaoPzEKK8huO56pvw9mi+JAU2FFKQIpqWfts5JB+KHnlzcr92X
JDGitIM8AUiKBFtHIRDcBmpKhGJ9NgkjEURNbyXJPyNuVn4Y18sy8H2yBNCHjKoszlnJSKGn4Wui
PktFVXv+Zx6HA6m58uuKZzqsTtvyX4zZQ+pWcOaxKHP6yJIZnaVLg1TnLOSrTK8P+IoZD62WgEL1
QYLtAOGvX0HYJiTx7iHC8WKLFz/6POY/kfzVTEOydOqZ1xXpXtp6UDbtGh9QBDsOubdNTJ2ZADV2
Bo7fQV0pS6hNOLeHTzwma/kUEU279Sy9Nti8OktfjxZEc7y9TZV45GQ0jNTsnZ7EEssbL3QJmwX4
30VdzBEkiTLJXbGLvqR+WpncqP1tMru5gcxPK8F7ieYaNM0KFyrV6LcsNdknJ2I/qWP6TAYdS/D1
oycws7uLzn28HqzC0hSOG6FdV1Wgh/1F4vXTnvvTV9CmJyvK9YoWTkgw7gO41ds8DikbDbbGqVUy
hRLc7al36Fg8k0rRxG7Dm7csQGBV01Z+l4vN66Vaw/TYBMsqR1A5IxOBO/q94cR/dUuQS77/NmeI
ob0Yy9/4B7uJiq2R1D3ozS2jxeCf6bxpSZADzITtXIU6ZcxDov1D3VJY7gmRFMt93p8NZq49Kixz
100uvFJvsZfChWw7LkuF++04gbqEcUa5QC1LT1ssNuVXBIPhc/eh3X9z/a74bmHz3ueXOGk4MmCi
QCsgj46zMv/V/9o7xLv3GKyacRNC2yZmyoGnWSm7AG1bAyEIgLHdsdi8b+bEX773VMNpciIa4DAv
wa9LnJYEZjagj1De/39L1ZeKA/EhgeGYkO1sckFfMs/mW58hoOXTlwh8uqKQSCcMg0BGJWiHgmpk
LqFnAYIetwKzODDyVWTNEYUG5qmLJII8Igk8p4BqESXjiYj96mMXAr+kIRMdUCO0RvLYP8NG8my6
Bs8jIm1a7VvtPJD3T0cJ1Un++ksjv3e62muzk+PdgR4SQMOBnAALFmFpChznIpmuQsx17211kXGB
cMjAxuJHGzEk5aPGAhdMt1xxmM2QkL4tTLXplklXo7VF8ff+2VA9U8oeRQl5Ty3Nzjja60lugiMK
qK1kD/ZabgwWmIT/3txI0oRrvC3RKCB2qt4/4vs5DpUpPGYoCvUsBxEvu1HkTysdJZnXef+HDK4I
RnQvnCl4uuVJ3OC7Ws+k+/LrwLLPa2Pccizl85qt17nowfd4zcLvveenzUQrEmctSfNWaltPKSBK
prJ9a62MlTRy9pszZQ+3WGWaZ0RjvL2KEM+OUfXmAzEbZI99RpXIE488sAhkd26NEdU8RRBdiyHa
oQQb7kjTZVlKs0rp2mJ2B6cc4odMSp42dx0ZOCSTZhNlePRJ8dOWYAdr9EuFYufzdxU4RG0J+XYl
pInfR+7Thv68q+2FiVaEflueB7jo+0rCJGfciDFIuQ+6FMi5lEDI51q0otfsMUrcnKNJ3W7V2PZ+
X/eKMsaNS0EvUgadcakULQXyX2v1xk2Jjk6sWUgDeypbMpCBkOxCiHfBdPWi+wH6tpfYUY4ymkOY
OhqLvqoYYiOx1ESeDyUt82vR1dHQMiAe8VHhioHa6FcKd0yobwVzLcfjahGgqqDMJZCpCZMYD9i8
sD4l/Xd5PEVXe8CxH81f1in56blV89Tq131roRaoYuLgY4UEj749IqVHBNU54IggcuSCDhM4we83
Ni4s9Buel6bl/0ehIRtA2YgsICB61YJHHl0anzOkS/u2B1XksvBL/owAhsQpPH7qPSj4IRjqYOLv
b45/3FCllYn9DTiBqNXIRgqgogFKhT4JRivXVmZFnK0baNuGrufx48hfOy+t3Msa2QM1n1FWAV1h
+NzU28fhxQaoPKE9a1199Bp7Qm1/V/W1RXVNfRQkmHTx296WrfGuAFZzr4KLecEOIhH3y906qqzn
V7OjZZGf5N0g0cX9rpD28iCxqBAuzYaeTaMisnk0tEv/G58r3gzDVNDsvjbw0sSUgwjNiveGTOnP
DODGbFap3H3Iadjz66IeExxXEMcGgQ8vhuaxDcTBPwyg8v70gF3egafrP0bo03ybcLfSy1rnYXFv
+mXECAt/b2d3W33Q4Pdx6xCM0cAvzGnT+6B3VjFAHcekEmt86/6ozxkt1TLLLKgb4c+2UAtjcXij
RJDOkqxNrMiexQKE8XBfnz+ntFJnNweQWLqx5HtokNeHcN6ukCD3UPCEUckAWFr/vzrHXLhfdFOR
yakqZNhAdD06Cu5n0pbpsSZ61EFUv6Ty5dFQIVZsff2vbGr1GhSPzfofW5GqtsrqHn+6ccJO7Xrm
YFcQ6TcF4h+O+ELktas322nQHX1I1FQGmVjt7+xTlGMNcfCV6FhcjsoBHm1NSQLTENmo4OzkbD1Q
Y097Sr1JLNKgoq0Huigf3hfPz4ws4kY4eAbN1tejq/Zn7n9+jSvRgHzu3dxM7ziX6yL6gj9S6NCb
z3UI4NLpeHwHgYujeT3G2mp0HoWsJ6u++aXAHMwB8kxoun5H1SdkDXkWZ1jEJJvHRkIyLBWRZkNz
/0jySr/di5XMw4rzVpLgLgIbVJdWjke1I4SAN6UkCfIT61gqrUTz3ct1zIWwYmrV9Xu2FHcAcJFV
ArRyduN6ZjMzwAXy9myqDQF0frE22V8lrYkC2jAiSSkf3Zay5CbPMYGvkeA3byPkO1+PrbkJ10Zg
A5a9LDScADocieQDbFhb4nbdu2zE78N/qFI8ADUKCU5L0INS9UyplH3PVCPUyCtbnbB21QcijayY
POmff7B11e4e009l+lMbZi7dr2GN970753QBIkrJeJo+bgxR68WGVUQLnlLLZncSC0sdsxetOjU5
OMN+Tr/Olguf5ZfVY9sh+hbA6aBQ6pQyjcDUp/0hUCnJFz0xB1g66cozuNqco1pgm4RMiy1/1QTq
bnwIZZXWuemHKKpj6KreRZh0J07U1yMzV423JlBCZbknwLVncvaR1+B8Qvz1pvK3ed6IinKkjywq
E18anJ/sFw8rSxgirSIun2alDAV5FBFNwn5xSMk9kFH4uHa+KwZ2XyHhqGhm1JLKB1BAHkA/3xq4
tmPqciOoe0xf7MBJaOdpc7giQmkSrCnAatHKS6SQEVSeNItQsiEWW8jbZIsm5hJcfKqa8r7raqmX
6z6Hm5+wtyBquASsex7Wl+ty76P9BWyRIsizzFFAC71TFlB0j601N3Us5LVCtQed1povRWVm8ejR
Npt54fOfosRPQZsqBbHOWc5Fv97XkakWhp/9ksYx3+xt4fZND93exBaLKY6LPOrpl0Hp3jiqeC6j
Gu1EoSxivckH7e0VEGpW4R7KelzR9x9zls3a2ZECyz4zZh5boyp+XzOtGKYMsh9rJTB8YmXVbptx
W3BgadFkr10jXveh0O9Yhpv+EVaYhk0b3v1VKZi+wr7+d/qTePhsPfbsqkr2xRRr7NaNvIiWKmb2
/pG/7/aVq8WYCRfJzPg+5aRdLc55j3jzbnPuVUJb1Cw3nRbe4FsBIRV2/jHZSnHjxXj8fBsiJr3h
m+Osi3VCzS6+qvE9de2UtL+ccceRizcV/qMb64SlzcbaNDoeSJfApqZnE+ldEwj3cvFJGYdYFnsO
OzTJXLqNkbH2QYLYUYaDhugEkirG8NBnvOu5Udi4SuSTWyUvlkV8qZxvi35SRKx7xcZBEyFCZ8uv
pkYuVDPehZQFxm9r/gGiCvjWR5n/LK6M4KV3K8d6XhLIJutouQhlTuIUMiw1IgMxxMGRaikg8BGW
T+7sARTnBIXNondPA/Z0eE5Zr2c4QbLrwTMeMgbTu1XWuMIaZKRkaZ/p2MYrzxRtfy05sAYM6U0k
tXWnIPSYBLws7EfKVGnWxGpv82+IZbcCdPHc4UgNIHWtvhgbmVQipxQdJ8GCPbHIW9We8VtPz6xJ
zxMJtziNoV0dy0QGi7rKDID/nGj85tsKfFYNcLzcX/NZ9hWja3DKSQkL3xa1ImkRHi5Nne5d7WEY
nOzGGCsSgJKFQBCel3rZdnGf2dhNgYvOL22IJ6db5bA/qg+WMmmflpcf5MwZ0k5MBqCTvMgzzPTD
FGUq1YeE69+Xy+7jJA2C8GxQCrHW++6/cd1FqFh1P7pgagXZlRtTNU5hCEPZ/CPsdjctOju75BrF
Xmb1MO2NRA9zdsrpjy/aIjuqwK1MSwlFuh5Q68ANX8A8Rn/XyOgt66Zut0sDZIkwAmZqMic439SP
Hi/j/C0k9XWAZKJs17TYH7xWerCabSpih/oicYWxLnFmcK40+VGoSj4MxE/GLhNUQhCMBao8kDcX
5GRRc8cdTqsJibmsw31CprhOQInHk8DyhAsxSgKXNGxzdT2hsG6Bw9vGDdYKHcGTOjGqqWr3JRWL
zjqbHHUEEe8hj7mAACqA8+RXzb1+qLUfKwCRZElISh7KCv5hN+4BFYcVhVp6Cxfe0EFTXwO/vI8D
gIulNmhDV6IRdP69i4kSrdwgHQWEPmBEcl3VbmwO9x9wkqMZuE+20VlD8u1QF07VuuSumDAjshyg
I8hNlgtqh7X5q6HCWZ3ekZWE5u8SHp3J96cAay1mIwd7eHuFgpPQn+gIb29CQjKrywcaoxLzumq8
NPNy0//7OGK3MG069gk47XCG8OP7orabc3PzT3Meug9aybw8tUta/2UadmF6RMmi2BWmKcgj5PcY
1dZWx9TKRS+WyzE2SSjz9nVRrtagpTSuaA7d2pUgZaQyhWGf1tMJpnySkmsF4NNZpig6erGlQyPQ
Vkz+UpS0XKo548CgGruyuOf7BeyXSbGqjp9/ur7tYpg+PfQ4gqPpMDnIZUAT9Ew5wE0rKj6pOVyO
izSPpVk0QP0f0hUotnqI9dWKcjWzGJS6g+uY3RPF2kSjx9vReBhPWMLkizsf831erK5gZedl6MKW
goOjNw+OV/Z23ALB9XDYFXlNmeC43lFOBFeKKRh/jbtaLZa8rAS4b/lOHeQmpcO2KI3ZO/HkRJML
Xf01ZUnG8vzRoCMVxI53G4BTO96iRpB+6E99DbBtKPcyScjnd3S7i3E3ji3wwnEFesff3u8UBEAH
D/bIeVfhkSNZ5MlCfh7aZMI23S5tIvnmhIA3fgeu1aTgP7BvDSCD90SizJou6VaVdkXUpZvAcbIp
ulH1nq+sqaK8UQj43GJvuEJ5JD4xHixXCeOY0CFHl5bT5uQAnc47mx6Lf4LnHZot5mSXE/wUZfFs
f6iJY60//WslodnTGUGmiQYYlBG5zMX0X67H26XbBLm/z1AUA/havm/9774kRaO68S5yBmAD5Gz7
CJMTgIN/GuIGISw7KussYKFnwAiSPT+tt6Su5aDWfBnysJ+Q5M7fzr7PHAW2bS9PDU8oZ12rvlgS
k+/wh7AcI5bdbxYBtLm6BgrYy0s/9BApVSHpymEiy8oELmFGandDpHrZYBwgTGU2rCmTVdcffj0Z
MDMOJVwLPxbAANRvV3M6bCoW+5Dpk8udIo/FgmJAeKK1RjN98V89POdkvzMURPa2p3hxB4QUq24p
v3wLAJ+/3oJbgQKFlELnM6nyf/e6IU2b5emyFvJRGNMSwz8F0/7BNGmszGBy7nYRqexuj3foAwIh
mNpOXMIjdb7dacOmHE6Ya+NZOuLVnX5qbmF7CSTBH8+9e+6MTrRBj1CYu8KFA6c+mh+ca1l3ietU
zpbNWrl9wFLztQsQogaavcQkQ2be9aFovHHGxWm5Oz1+n8RvhV354XmUgqp2rEPkLTshl47LJ9xS
rZGp2Wj68FNT8UKSh5gAFqGkd/xJjcvg0xQ/vp9NzKZ80pmu49anYct9PAnmp94wtQ2h4hUECps6
S0hPKpIvCutisEjfui4PQlL/xkTR9J7K+lsObg2xBi7L2ll8ShYm5WTNNNF7AvBsOYR2Fdvy0Su5
EX5OZ382GUWmDdagegLTEu/dC/jhrYqfur/IVHdfIn6/X/rv/8m8WlNtemuBS85b6WSmq7/6rgSs
zaP92sy+gwFzBfVy8M7q0E2LaV1OX1uevoMGtZXI46l6Fl1DuHTZ6OG6uRdTRw6wHaRfUC4PsElC
uzquqj89w2t9kpzVPy5OpC+6/gQIw52TnQ6DbDsa2Ws1aEgwXwxPiU5+AL8LAgPrkZMSB4PMBtDx
4xjKk+nrm9HHPhJWN8FXT/3/G8xDB/QY0Tob3YC+GJ68K1kSv42xV/DOcHLeBx3zO+IAxgFNLr6/
we2C9+2beGD0fpRylZlbWjx6sPJ5MGeNZNJBOwMf6qQIeNThq6H0vfZraE7K1M3dIls6G1t0fSVf
z5agaOvscaspej84p/z3IKysrnuxa2EoEeTDxTHR3hbce6FfQCdm23cLSoHSt0ncYljozOL2Lntd
nKISDKNbm4yGPuW7CCCm9nPObNNu6Ytuj0lgheHO5NHyPjFdRVLjzTKsUA9lC7pgMjlh5MR3uL3I
kxCQGY/PriGYP67xTn46EgETNrgvAWkKYPg20xo6pegxVHOItBGB5c1NvWTrozRUQf1e+2vZZ48L
JI5uGOE7aEk9QYP6D6mYN5eWPvAebIn1rf8K+yp/QNScKgU4ux8s3SqjypJJYfzqbZ5wl4PzBdTE
ZNkHfR1kUlUZ+09ci4kzXgZKetUiH56ItZNDfdcoq74bR6vNZ9Q8sbBx5pb/rlF1odL1iKuFLVj+
OZri5dVZ76139VnYyzrlkOemwpeTgq2aO0PWZGcxNn0LLX2GhP3mksiY6XALfkNk4qb8jilsfLc3
TInL6YT2rDq/oNPTMg6FI9xT7HkMZMP62EyqdV2FJct2ReGN8zrutFZw7C3EM1ykJ6rNscc4euFL
3Ri7wgQh4IW2YZYVHJbQWb+j0iDmX6yTs0L3Ifnc9+1sBlmDE3plI/LX/kCta7AjCXBDsNc1YzkK
2uKdUzpa9+fU/TTBsN2Q+LOV25Y0zbFg7dS0yOCrEtCOwqpeJddQjgF2jYkr4QxzUTeEXNPcT9Zb
dhLrudpUIJ9Dkttzbm/mfew9pMm7tE/ROH0g80et/mUpJw2IvzpD1Di6XmQYpRkZKLjO+//CPXDE
hiBzXgSRFoF6YvW6uK53bRE0gT5BPGaeyTVWCJaiKpUPE4KkODc16nzHnx19eknaeMIqpwWEmo+T
CKcJXKmIfiVHhbewxJMszkJcHgsKLpO04OXeFdJfeQIqiaeM8LVj75P0sNfBspGV2jdV3892GoS2
ywClP8LdbIl6gCTmtsDBc6BQeTBzBBgC6djGyUkbYDORyT8m5i9LvkY7+WfXSE8v49sqbdZkrftR
8abh64fanMKCf4JjAfbRXNzT2QoZvMG2LH5bZpT2DyqeEzti1SecBWvg0KRDkx8EWXSkX8uxVvPF
xJJr8xqktN+9SFhLqDjlIXAklod5JeIXxB1XlY8KdnZdlXZbz43FHtrwLzCLT6v92n1lAd2GgCxx
q//kyBt1nCObu1tpQDfvEbKVHwXBVzPyDd3pFppuffJsPreuTxxoDdrtzOEtNcT1LK9oyVBSHbjY
1Ji9goy2ACegRde3bUsjbMVDIChQcj3Sjv3cCpTkJ3odkLLxkGpMxO7L4PC1srnHzzZrEdjJNoX9
wBSrixYcLmKgmuZIEg8xUoj/N6seE+2/3Bf6qy0DoFrn4hDyY/SNSEkaZD3VyGBWN/7rmGJ13meB
kZrCj3zJMDK1jLud6UodLGJcUfoBEMP93yiSRMYZj8e7ZGKbyeIMeRwx5lXUrq216u06SRIgvmra
1k2FyY4OzfKyfcu1509rboWHLnpKl0RaNRxGNxAWG543BvGJqtvBmooAYUOuzJwn3weS7H5hTKWZ
1DAaaVJiRDvtfUDwY4XxRwuLo89dUNaCjM96Q4DT7Iy+AXA/xFkMVb1I12TEkd8HAvxtsuZccfXp
Vs3kejMAA0OW5G8m4AU6I9iXB96T74RVkyIkC0AG16O10X/GalM7Iad9fQtLvAjm1kRKm+sRanX2
r20d7LTlXL8DEhKf/qwxUpTX2YDcuCmrQIu9iDdCCXQ9+L1qNRAufJI4GrS22dmGM7Lg8x/HTQS0
hQ+n5P0O9R0pYOg16u8bpT8Hm4JKNocRjVRuwwOjVRU3n8o7XY29EnZeN9BhTJ/sq96Uwndu7kTi
vdycRmz9sQWyQmm0sRrgsQizI7iBeS1RUmk5PYS040mEVJBW+rgxPQhug2ii4SPH7zaqN5NMikuW
Ob8dniWXWv6hy9oDYAWoMjtWGEN6lo/apRLNkuVgsR3e8+BLJyUS7OceyN4W3ZhrcTO0yT8YuEiu
OQxJFiJyzOf1M/i+4h1UXc12yxtmTCPDSZKoR9yscfFfA/PaV5vps4zwOSc5imdbWvvy+Bfx0N+G
2rBi9Nkl1tCY/6I/bcpRUs/czcYVSTKbeQWK+DjWnoY6IMqx2Ll3NNNaL+IXZa8pUycpvzoLNLL5
G7Bmfk/MTL1heEBk2eLyaT8OHnpeLJn89S7mnkK34prYMDVm74sTY7aAyVjkzyJ51tYNpxcoqkjU
pfX9I1CDoCFX8qvaQzOPbiZAQ3+eA5rQIwSO8irj8EqRvkp+bEveMismqsGEXU0QumngpSm75vT/
TUlTUSGyCaaZ6X1ieal1hlLUY+i0kmSq576fDvWFQQhAkEmknKLVV6oP7JLdSb88Z1Vsw97jprBB
vxCBIyZN9NQGObUWpi8SxUGcMOdmIGbb1uOa6RmHdZPVJdyPvqkUTcvAsjkHQQW8j14fi/y/8uJd
DfissotBmeO9xCroBH2azFLSEt62I6cb6wAX1lqJsZOjI+U12cohbBNo7xxejyI+SmzA7fU4CazD
TwczV3pjZpF+4EQSdaW9L20Aqerk0qNZwDg3q817zNpuNSOrjT6aH5q3kSIrae9TlvtQtGdnauFP
TMK3NYAbO3WRfRHcS7lk5Hf5j81WwnyDICY5BK8m+BgVcN+ZMknWZqCenhzkuZYXg2+lihLYhzOn
P6sZWKS03BnB16y4EAOLeFJTiQWPlVmN/ggTcYwZC+HGZo5wk0TkdYqjZlSjngy3/UYHscf9WN6o
NHtGlJGEZ6U0Cvvn2REn9Vmd0O3YGT/YLzBR9P//klkbGaWyTLggPvtERGR790tI5EhEHLUMASZl
+zGFdiAL7z7NATchrdXebJcBEIl2EvlSe0496ZbVT5gtHC88+CvOgugS6f4DzZBgUgP3m7iNa9Y/
QBk6t1QSlFUKtnHN/LOwzK9sWJKOqnH1P8IzsXNXaxK2eTFQiHI9wSJVDJEkxvBiiOtDoCEwOjlV
kd465ggQLylQji0ASrIEfI1LBPMfNiO5AK4tuXQ0NTX+4rmjiwLat9kok/otbczKvLsPsbaKaI89
mIwxXTZ86lyniMKGyLdhM8ezRVeq2gUM9t+iB60D4P6ZapNjkC3sgPWxuBhdQzQoDfCy+RrIDXkr
x6HCczPEHhcX5l0s1FlywvbDYudu+p8N8XuC1mXWBnJjH7f5tW3bHgTaAR06pMeY7ojeQ+Lr29tD
bQoLxpsAZbhEWOxfT/UrOiwTdU5hi4jCQYmY7ykIzMy54GzfR9C++i3IiEE8RFJ7Mg2m+q8EkhEP
tEvap+Wg71dOubA8r6lJJ5IXLxOUpxqYpOn0HzYrnzpBTGL/CtCVORW5C+FG1Df6LhcZHN7yzUv1
xGVcGxWQbQ71d6CMjIWr2WcSYj0buQLvonzuRjoPL4HSxRRQGWsMZ8UctnDs8ujKJiDXmn66cLCy
5z/c6bzhQu25gS/HY/d4xdq4qbwyBaoe0D+6y4jUfWIaC8eNW9kFK0PWZmoH3cmvTZSSeoFYNfpD
H8wuxOnWzNmJjeXc1B8Dtfh2T5gDMTA5Oor3/7SvXNarDjrTZ501/uHy6fuaC6C2iz/zH4+dJJ4x
7vG11w4h5+R2LBEYgTbwdtTsrmMEL8ZXuWayIJd3ynOH2ZgRpel9nKfqgSX6ApWtLnpvif5MP9IR
xdZd2llOVV80+f+YJRJzLVQO3jgqQZVHLssI5UXv0KkMrUzPQIcT4aBWiHW/0n+8+bQb8xNxga4U
eBtYMG+ZMU3XlUAgWsB+IqyyUKV/4YuMCWQSZxIMKgy4+CyYUWMrE98lGSRbUT+JoLWkQ3QcUtZ+
Kk+vZeHSmJdApr7o9dOOHO7Ap3g8c6WMuoKWsv3Zf1uKHWiYWK5QqDsX/nfXWdEBb0l9whdUw2Ai
EiTSMNUWEzm7v2ja/8F4sM2qX+qr5FCjedTGgDe8O7tEUURuKaqOVP4w/wH9K8wliBNRaHHmhFHx
UMR2ywj28MbNFO9mN+M/vgT3BBlgGLWDnpXsQuPVxwLukCbrr9XUPXGcAh4xuDMI1NwSYhMuhwGm
GsH6CtaQlZvguHIMFZYYbey8UDqGg2qRzn+yDG7qzlc1EwLki0cTP+GPQi9ZUkHF9SOej3IH8IQs
C2CKi23GaCO4Ls2cUWRwUWD0QV7Bs7oa5r97LfGJym/AGB/XSptIOj9WrFNfwRLLyTlIJvWV1NRE
O3c5O7euuDt3vh22AKdozfPcs4OkoiEZ7bbCCnpnktipBI9qOJQw8b/EL2xqpujjz+cfQEWVIhmz
z69wbnoyPn1EU/XyKz9+y+4yKhflFw+S8aqqoTghKoZaYx/5v4v0OonMg++mxJXVlsI50xzbKU52
jxJM0IsweX+6DKm1nV5UupWDRRe7Qe/fOAk92tDVvbMJLfzFV31pDc+1gwK2WQdYd0YifZio0ZC4
fHJ8ABw7wsPgTh84mmPJ5Kezs+0p7MiA+B06cBfwJwLsMZs+7YS2Cmx1tKHbKeZTmjwgojiaU4Xv
e9q8HeWQAXaPfHqrnbBRwDrrvehYj3LpPeIS7NZVz4h8S3cx3YluTQOQPDO3d3ve5q8+ScAEITOD
+rKwqoLo7G8a8P9TqwI903WUSzk2LBKG9L/b39FC4iFQIL5LJU5oYVPWI4cj4LSBBS1bXivOuRNP
BG3UNxiRKNqm3tWDzERXsmFaoxZONaIpU5hvNWP5EYxCB+aGaSRyoBB1DWb/qcEB2CWGx8HVTqQS
Na6aepVLrBgxyHrrJdO5L1JG7+ld/ZUFWkVPVAiymObk/gWLBmxZzlsUKd83NBGlBho+MPjHkeJR
ZiajHMfrN+84vL2uM1gFZaaCqZ+sO1NWQo6EFjvxzWd0pzUiF6Iput6QiumDbnPoTw++I0xNbI90
bTRvX9EXaNbZW4rLauWrtrSt6mMY44rREYZ1sgjhyV0PNc8PRi0AZ+4+ssk+Zzijd/v2r2QMMV5D
p810fnT+jV9FQFE05HqISwD9/0w0Z5xjVVe+ioeDgVOPn1gVWt2joHSpVnaRvug9bbb/7BN4+rtL
wPO7fDag6kCxKxPFKDBc8E1s3KXU8bVwq+FpKI8Ut0o3TVi1at09Wd4t14gGQx8GAxfWxBgE1sNE
xNHD7VNLwyr/95ugv5n6P6pRzIeL3L8wwf1BumqGc/I/r2QaG2LqaXtCARqlgWVwfFHOqW38vDSs
mYzuWmYM1AG5nVxvjQoKx858bn96/3EzcSt/Z/OETZaq+eWGMHKhSthUzqIUsVglpys5vIHQuonh
B+fqxPZSxKeRb9wVMvcacUKSkjIxTE56rP1+ZYZWQ+UIq48QE8GfJcjGx6iIJkHycXvAN+SWQZVN
Fbe+iQkBYxRjjb3fLvLR6Cc6SvnxxEAkeLZtGh4zEicdOqBPrfwTcFvg+YBFF7C9Ao7zOIZwixa7
OH9uaunBGQz4Cx2/w++HcuL+2YGc1u4c5A5EyIWy3EhLdvJY1gK8bHQaTDV66UqflauOX2Lh80Uu
AQTYefkd2g7tZG2Vo1pQRCk505zAnCaeGNtQ+hiX46xAhnlBCLK5mH8cNKeHYvf5hM9SGFl8xPaP
RjdwAEphax9lOeyI6oCR0NEA3BA0TRZQqBfSc03PnmflP0qcR+Gj7QC4HKpFdoEdtpjUhFJGngyH
lvlMOJJQTp4cCZnCnPuYuDkwrPLa4YIdNGaLT9y7Lz45EnDaRMmWxdI/djMbrvEPEwdbCmPhZMUA
M4LQy//016aFRhf6jLVxvQy2UCYZkqOMceUx2SbeSmPlKMi7JFhbQK7vWHV0hNby7DDItgCYR3iv
YGOsCTZUQ+dDkNrwOxuNWNDJkRofUI5wEJSuhU6K81wu6Cy4XFJXvvnicEZdyVHTzgbGSqT6NTpx
uVQ++Qz1ezqbAUE/fui71uCqQTGUpO71VmVCLTCz0RwWQFdQRluO/8xLBvB91MfsBFt6+ApkWMVt
NZwCbRt3Db80K5a4BMLjOJg37Xv9KhEevgE8+VipDjWORG1tTgkgiU48TOPTaI49DYtD2XlCrE7j
b9Rk/979xhT0ksD2r9O33YDMx+cvHu2rtjPYOnG3DJ7ENs4YHEiOAdpJclKsF4A/USGTCG/SmDbW
Lhz/dx2fV2aOp9L01SQRIUKChUCqavB1qMsF/64r2YteWyW9ACVHbIrwWDDm8/mKx7NENMK9apsR
23MU1Mvjxyggbus81FFu8kaEr+UT8mEGsV10+rvziiN9uW7Zpepgd/UHdOX8ilMUogg9IzSobfSn
S1wskBSqECOLX7l5WMCaLPYRZejWu5dxE/AifREonYmxUghn2vXm6uaC2VS8A0/QOUoqF3K+Ue8/
vvyzyD0hkcBVcUPRy5ju4Qg54APj2dhLqg0giZqW9vRjEbfOaIGj/Oc9lHDTGyJNh0H1jvwNRMHT
kf7q8Vg0u+1Jn+Ol1IGxZ86LxHda3+zxRB2bn41HysE2Zm7k2bZMVR+8/zfLx+IjrknwLjwkKeCe
ZJ9MNgMJPhy6N/JWiX7ZeGtidMb7+EyBaul8isxbwNWHFhzAd9DcMj5sDFZF2K6pBV3P2puDjMNU
NGGppZKK+71ITOjkbryZN9eI/CTN+W3vT0svnUwxJoo5fCOJQvJ4TYwFrPlL0abMtoHQHrjqvJSx
IF442qjs0thoZK/XxkHYL35d9Ti74JHfGIopEUA98RN78qWEFMm5eb78wwTX29eUo//QfZkS3TE+
dAXHjd4+7K/5SlBK1zhpaILJu3eBKnHbdE+jj799J9UfDAzHFJPL1u87HisjqD9r0WTLa0Z4MWCX
wnNmVIwqbaP/jYYChQQzjxNBtK5rrQ3KTLPNEPLG6GD3Lmy8McTIcie6a/ZKQHJu3VnWTjy6oI9V
vnCWpYIkE/73UlHc9TL7MYQgIEHwQZNs2BX3ZY7JTTftB9pZmzv553OmGZP5JPyEgB5zKT+d8cOm
4YYIwNy1MTeaUJymZViAftZJp9OW/ElGJHXz9SdwAdEEihQf8frDTHub+SeGUcRFw48LkZJvGQaU
V7ngQK1H/Ym3vJEQ+NmUVK3vsOphVAxTteMOzmzfnc+ZNBk2kJ7xdWrlHNCE7mz12fi9cDn2TpjP
FRPBCUplk2TUy4+6O8RVn4tpA19zp/Eqov1qV4WzC1pBo3APhReIfAgNP/BJmXrHM7TP/hCpIBUr
yip0abiBDELSY4slkz6ZTuBPF6pZgyvyuKOQDIYJ168SNqrR2g2szsqk/2rK2UjK1HGq1Gfk6Vam
f4f/jTGjDq87A7Lf2RJYuE0OsN9cjRNod95jCnuhBSVFjSd6Ulu67X2BA1DRqpasjj7KvGfHLN1x
E1sOAwoo8GPjIF/UtbeZ07MgDuKeGALFW5lNV1VW9xV3DKZwJxtNoocs5rTALNvNUqVrfTdTAhwA
T1qKlC+ge3fRjJ+GJdBCCQ3qG7LxAylfJqCMy4HPF8nPNsk8dzHJydBHGi6hkIai1a9AIzVZl2R2
7oQ/o46kzs3jIU1aTwSFe8pjZViRoujEKPjSY24PkIDRsnEjFVQaATmqLpQTXmVzATHXvKrLmV5O
wNmucygKKUE2XHnSAhMeOmsUd13NYPC2hLvr05iiV5T3gEanVUaMQIo8bqMXUXm1GlFWSoNz1ipH
eU+5Zh0SSqAEDc7mmjyOE5kv9W0okfiL7Z4WPW/MiOYoog+xcUeQf+6y2gWkwRC8G1Q4HBhmize/
rBJgFAKFFm8Ri+ud5I0Cyuhr86uj1KXFcF/W9mDsQoqxI77PWpzuwh3Q6RfJYtRh0Ly0pYmA4fg2
kDUFo0dcrDWKedfOjix6wMbZ6VCrN6jKmddcfCwVYYsHW3vVVTlzxL6QLcYBJWLDPmG8qxLKmAtY
9CQX8x/3wxhNmpY0LQUxsGNBxbRRwJLQ7CTrgVQ5NONeTStwys4S4X605JbE2zoJcrZ5wVtAWAQD
j8sYhZW/9LVXugV//G5Y+rUguMcWCfe52VNFZWO7LSlieb1VYnpuXd4Hz+AFveQX1XYeIxvqJaCj
zPwx2EqQugO5fsRhikPxy5GtjI60PeoRQpZAplrs9cFlwwhHVDhb/HDnmPcwMGSYqx82OAcVbUTX
Gjsclmiw9YR1pFrO2x43xc7a7k+J48S5FD3RptNQLyzsFDKVorRKqVxYrK3zrgS/ZFP/3Nd5gDCt
L7e8nRUIn2PepEmL2bySuGnWi3CoYblqfqReH8crMZejZHDxGGOcLIWpvn57vAucvXDM2DLCEuEy
HDmUGrHXYWeyiZHNQYazPKw2/JHsmjzd9UZ6dJvLcFI5X0aww397Tx/bxo4yDXsdAR/jLkGnBSsk
TrSUNq6fW312AM0XiId77GEcTqhfr7n7vfP46Au9b0VyBcupyWuAtjzrWrOtA5APQmANom4hKjeh
3PSDAMisiSQOGfren8Lt+lxfrWSfF8/Lu8u7HnFLDzusGAfKxgMY58N8K7kGcQ1bQQL9NLN9vHzZ
wvAtYoLptbNcJ4gQo49Si52mqIpiU9RrROzUVMAbz7+8/R/nydXl90l51iHKuVXM1fJAm/TLUIid
APLCkZBfuBDLXY9aSBtjNYmTaYjh76j8DLCLQmOiBrnOLVfRBpSYhiI/D08wsBXlw3cUA7ZsDZm4
69hyXTerCtq+Z/E5AIjVfkWDCk+gzGSivtxPDhv/wS49M6UxBq4p51teOVr54ADAQSk/9yXoAnof
KbwfmK9LU4uFQZb3PfFaYu+IDXEKoXCN6ABXJCaamhHrEnYDSfsBwY9UT7s3pEev3XDxx8JowOaI
iUnJR6YRUAO2qSraBZKi1pBASziOJoJBu961tJX2rjgxRT54udAiU1UW0kQ7WEaXxkIqu84+YSWH
Y9pxvdBJ0DpQymSZy2iR2SgMwaWg4qlprtdQ+YYWz4j9cGRE568juT/Sz6tS8CNsFa3KLcSRrraj
eNaZ67aocWum9Cejjvnm0YUpp3tHkxWNbOimh80INP0bMuI152NobU+dxwCAENb1XPwL/hD3xiz1
UM7HXgl1m4kcJl1JuzYV34zle6i3EkHQmp1e4XMLTTh+PLp47nkKlQiV5KL++U02/7gV2qK3l6rO
n+fGGRwth63slgCYnE/AdVZIwE81sm9XAzAS50ByGWTFlEhoeum2JqAwztwsKNIG5pQZ3jhQQItI
l5cqmYnn/buA8Od3fkSEcGDGa2eIc/T1xDIjd+84rhPtlZ88NmsEsJbcTSEK/C6iyn43Ks6Dluac
/KRTNc1IxIKg8yzlMTt4GXcvzxhtjUEuxaFMU4BlEB+PWufo3xGZ8tfAMc07q7hX1wfPYwVft2Dl
bYOVVgaCopEr5Eq0fGmICiTBuDKUzOSOLkU771wYlck88gaadwkZJCD0Rq+apK95WfELMSnBesVm
ZL9VwJcSE+/F9UmMzVykP+iwF3kow7dph6cWZ7ZHJ9aB2uF5I4p1tZjq6Ztp98Lg7PSjnywLpmDb
WSuDeWUguhy3iVXkmNrJHITAymqaClpo+ctrOQPu+TvElzaoTm06hH7pfYIFryWfjmekB2xwKvsd
2zhKIYTEQr3JThekSxr1v8aulrVl6+Mo7IAWXQoa26XLprIR/ROuB4iEPvpMRs2Ap1+CrFWPI0dZ
lNhZjDXEQpvLLnojcudlwkh0MYqWG9wafaRyB3FZ9Qfi4AcMdZVdSOipIIWcO1xxaUKxetuPi1Kx
F8P+epOjB0VpzHFxHRt/sOsjgBMK+16Ma1Nf05BtZhf6rYu2gr5gt1Rh/pxG3YdT3mpTm4jMFb7n
dVu+euK8ZgLYG3axxif4PJFuTgGk11siPVathprl2HiXl3oRBOjF5mYMw8qz91e9Tjp7eAS5YEmn
i4PP+h8wGhzPzJrh1TCkgW/o1htm6vBASmnsz0p99QyyBVPxhvjaKdeEPY8p7PJ00930mJ4ZwKF+
XhEo0bYkC0a55/OMHA6TeNWMf847Kv9nH2a/hgafm/jUQb+NN/pZbrtVjMTtu1wxrJ4orwkkI2pc
XaebxIhtLG2yC3aTQyOEloz995NmSTh+Pdk/f4C3mUsWHTAo3TAKz2OA+fDzygEVTC4N4COLtov5
Qm/JMC2SsssLrPrxiJi8KpYnBqbaJnSghk8Q4KSX/Wc/iGoMFGxl4HCM5wETNmHhFy5dUIpSXHHu
RC0zmxknF92d7UHRckrMfOkIoHmVYTVkQSKfkM+5TREuN9Vbkwy41LAVj1LijJC0tOYk3rlU6obr
ubot0eHgzgxsQcMWM9zg1wXaL7fx6q1IhUSeyjg/xgJuYL/LUSn95Z7SdBRBe/13piNzwUxtXHrP
Hdf00GE0/xPu3i7qr/iQ1HAzlQ1H1XNIZmEfXULhGabvWSS2WeqCTDnZZAASDUiA3DgimInBQsvx
RYSzX8HKfuBZn8kx8Q0a3p0Mkleq/R209ofTxd7ExMr50BL1QSl0XR1EVHLLmM8Rqz0a+L36URB2
izEa/rHGyDCCfwI+hEPDOBOBDGZ2C6/BN67AWmcBOGcVrXZ9tbVGqFhwhtDal7gX1yoSBSlBPxAV
KZ5P+VXfbnei5l/26fFSOYDyROvg2+nttLyw4C99CN2IQW731c6eqbyvCl/Fc94GLgrmutbTPpd6
x/XhQG7PSpPjIWvnMX/wkiBzBYWTb/CeLyE1nB8CSbNYvWXAnOH7NRoJKS9aFA2VtOcOMr5bRp47
Ekf+cVI5/4ZIvU8p3+sEaI4BZA7hYzoIzovVMjPX6w+RCMOtqQzyEJil8vBWL9Y/aTL7A59Fn2FU
/hdAyH6Pbovb3wtNNmfe9xljjDlvS3ERC9I4qPUiuOmsu6hDmaH0pDMKVGuHmVWE7wv30KOMG+fa
JzDq3u0sWifoWWX6AtIqAuPyaaX6t+xMw3IKk5W7tiNUjL/JWhmCazM8Oizjph81Tu1t9n08CdV5
me0FqDTO0qeDocwQPmkLji4ysgLjJYlGTFlQ7423y82hZGJvrjNSA72DYgNiNTnAtEu/qRpn5YCx
LTQ7QjTTK1HX62sdmpw2qiZPxFwQBLpssl6vIvPkanm5mOQkI5w4hZAolI/W1ZnUzQ+4A0CGwMdf
ipLNeuFJGMMCrzcEv2PD4CYT2GptSlRhvFYJvVNjcKUeP4rc90JWJNjsul3/I6FbhdJ/XmOW+v0V
sm2hw6kdygO7zH9jmut0D/FnLahLoHxFRjsMlQ0RF1LQROpwoJGe7gqAGc+eeJO+H3c+GjHodEbw
WRBjpBmr7rKoXEH34BbsEB7D+J5rRs27gMSLKzkVjln3i/yke6UZjOEsxthqW3d/a20X/yA624Dr
Uzskv4V+3DoQpVl3U6phLs1dGyMqSI+ohDPMY/Mn0i1ppnqzg/LkD3+d4smLIPzLuhLyP8E8GvoS
2nhhUS0/N7TMA+aNJ8FFNd5vt+/adkhb7UtDJTTNW9aa8WRgULxAw+I7n3mUInLVx/KL+6ejXV60
nm4li1gIsItEUIzQ4DCiEvLMSRPoKAI6YT3xpyqC0NVU7lxVI0k36Cxi+j0OCzv+9/0BY1tomhzZ
pXxU4F2U679dhBuYsogF7a5eJxOXCpLjIn1qdDJZpWDBw9tDlcNAWGM76WMiSdyHHMImBqGimc+K
ESVpgs3THjKX67tOrWpcSSNSm8vt/OZ9SQwIW8Gfwo6dOffUil/1Z86zjNhiyRNu2ww+A44Uqe+X
jkS5gb6H3Zf+ih9d1WlDTM5GMEYElSu66SDcUYunMVZuRNyLk+kXJWOzg+aQUPLOYqHZXjIae5nN
5iXHc++kdxg2yxyT7Bf0pZQU9jfilXZmKwK4P04hP0O9na7GfrpAgoTMMSpbrkAHe32XD4nxkwVs
/21HDAAc/KeeupAII/tTzTWvl1LPfPqvGGa2A+KdkiNUY/OMRJxmtg2eVAxX0jC5JgfdFQOQMZiD
iFIE4UCenOfIJ9xih+oJ6GcjtxJF3Z9U9oPsmDk/BvwKfGr0EvLtjYOIU/1gG+H0SVqx4pyTYSao
yJfSFnMdSh+gdxDm7jyBuXfj1zzZ6/g8eFjnn4bblJezfunMwuHKwRPDIQRf3/VLErfyiparaWRP
mejZtV5gUraK+NPSAsK211FHlHAlPWf3d7p1lYyHSuHfSWQ7ijxj3mUXmY68hZc9CcU2UpmVOBvi
5Na48V+fhpDmd5o8Lp34Jzirb0ODDxMoJbTWDznZcpY2VrQCiXsjaq0KeiYqoAiNkLEQs4QfySDv
dzaXe7/kw4p3/7qtgZnLMnn38F3A9asAEYDP1dz5f6zOzojA95TNYVi/qvdXjMHCp8ASdhOX4Kr6
5NyMrzh2LzyvLGsC2Io1v4tmUarzKJSmxjTaeZXUpYfe9pFsw8edCGeBNb3TyTCreYlpgmPJeoc5
V0NkOhwA3VOi/EbFj90wvcPKFQnSId5a46jvO3xBU28lfMq2t5KdjxIEuVWb5jg6GLz4z8Ns7J8S
SONlxa8rBP0+BjsVdtIQhXi/v+p+vNyoMGrnt81XXTqcXDri3Dw7DiVJ8wF7wjar8uAovLxYymFi
+SbbyVrztyJElWnJupYkJR3SmzdTPq8WPXREuBgFNd7zi49vn2ufwLt5GQpF0RiS2Kt8IJwp5Xxf
7nURIT37buimJj0MidMAYzL94geCSIbuXKoIrgOCqhMj9CB4OE2ZFMRn/mIgnB2EnHbHswTkoyoa
03iq8voAeSvlp2kOdE5Yt9BvYS44okc7T9Tcl8HT48/XSmJ01eqehhfp0ptZ/20lHd/9BTXe+tqU
Pxy77CI7JSE4a9CtAIsFbsWE0nDAshA9WMoY1FxWiCj1wC/JeREtCbjPx6p05VuUDwye1hviyQfr
KlNACIDPkS9DoOKSAF+2EkbqTnm0iL+Bj6mooDj6PDGn/CyLIfvybr+PYVh31zpNRyfyHw3WStfC
ax4z938cHpIYrX+l4CXjkeePqsYXFC11g+P6e340OhfhcJH59IIKVqZfoEOEnxmIHEn3leemb8gT
e4AVn9JNXVHEtJzNG/Wx/+ANSvpqQQ3dWWNv+Xdha3iM9+obUMPyFLmf/vY0dhX0IcDjvl5CPkf8
61GiCmAqd21WDm7Xp5D7qVVpemtYI7ofWhG5s11c/TofYqiyxcufjzqG+hzzgBSGJQY9ILyLDUzZ
fI1lAV7HOujsIV4iqEJscvmuvlgy3pFB9SXjvrSX/ch5jZpsWejT98i7LGZqCY0X+1JHvUU743qo
vqFVoDBtQrvF7DsTAc8V+DiLXsc6Eh6p+DfWgbHaoIZvTNkDK2AGITF/hliqWcZsbyNblAY5x0WX
ZGAiEdvTehtQtqoIq2Cu/O8D5F4lUV7goTPjAPaGs1Sk0/8eMk6GFWsE5sXIZ9cISb5jcaBowrIC
39EhZBr5ELc9W7L05O9phnehdCe0GocdDRoJS5pL2Uoy4JR6cFMmU5Q61ClaTC84sOvSjk+kBUgu
wZ4CI/D94oRtpt8L65KKhzl1lQoxKjmI34EGcUg7JyT3GFYJHWbUXkK+1UfT1qcR/ItQaxPgJ04W
xt1zDpiOazm559qunI4PXsjKhzCwNEXLwftSd8sEhBPbvelEl3NWIV2fLp2U+Ej8KyR8CQTVZ3uU
tAca5SyHnYvLfbYiFPd8dJ8nF+5IPpA9iaJeze3RnbTIpKPXVBx0pDDemWOAY8ZxnbJy3A+u3yvP
Bf9Rlw5LpRwW+GkkTh9Jo0Xf0638DZGwUWWTLQP49ZAXb9yM885t4mhxEjZ2OnN2QdN3GgRzEiiC
bw/tO8ko06lIGWVSq2nyYnj2ngpBl2poDwMbErdshelJd6oS9HFL5PH+8vbCeVFX+gqofrdbhuyu
Tq4zaWBboK4NY3vOori1aEvdPowuiopvpp2VXDVmsIrL/icgZ08juw5USmsIWTul8WHJl/FDs6Rj
+NUzIKbSwpIhgc+61gB/75w6M73TZHxMjdMzTN5TOok/6NLIMkmNLAI5+vImB/NKHRr+5acGjC3P
seUmwHOxP+alyb4tD8RCrW4HtzGB6WOB/JLB6201gOUFT49LXNeF/I7Q0DWQlfkC38XRc9ajxCZO
WVF/MWY1D2nxlzkl6Ta8NEG7wBvdzw6zWAnMCvIttKKLSVwKl1WiVDCeyXmcPCFyjbGRL7zGlg9G
h8C0cMJOsNqVePvH8pcO/97ek5hBrYNjBLxSuGZQRZVFffcKmNsPbKOXNx74jsm7/O4QL3Xppcrj
wJ2Yl5wkniqMoOOXaC1AmQZe/mlDtq8Uq8oG5XujqFRg5kwPLEaZrk1lvu+wYI7cCDwaLSRkINsY
UPCITFZlvDYnkHQejewuROTAwKhUxJZXKkwsEppbJqC4fr1XKYb63nGEF9Fy9VEt3QR4PNW+MX6C
2bwTfflyY4cl6Q6ShSGd6taidqKwEzomeRDZ+fNvdumX2FzFDnYc1cTh9ViC1cg8iqlimX4IP5Hs
8KqvvLP1m05BJqMZmuKkr42yYMRVk8gB1KDBD6jBTXYAY8nFV6WMpGKAytQo8cGqYxNHWD9u3eAv
S88zN7kc+2QehrRtWyBGzI/yLXDX3lak+9Ae3DrrV7ADuuk17isQgdlfseARQeKJB1XRgAWjBcf9
nzf85mIxxZySaoY/F5tun0a6FQR7ntHNakomU/v8RqIxf6YJ1wMefa3i/A+KHdeoTL+JP5Ty2lf2
5ALhO6QzCw2TABPWITun2+0j9F14tBqtc2woCLnZVZbmZ15gdGgqkGMpFi5Wy4gUzMwjqfvwFE7L
PybHUGmajM4zN1lI+lCLQq7vfKQyN8o3UpHeRzmJI8T4OV2ZPAmqo0nN2hQKeCSYBz5+kOgQQS3E
kfCXqZBI9yJ8KX0hSOUmtBvLii6j/hYa/5oEf/k/qRzB6a7GmD1vO0RnzkIrXDbKpBRI7ziJBez+
oNqBYXD0a/P2fOhEJCig8yOOPPUBWPW2Zb/0ITIdW+PMDBChXk3nPX6PpMZmQwUgWmSfMDPS15SN
wCfCp0DO6BZ1yKCV7fhSNPdQyN3FCWYaClH70zHNr8h1i5cjzxUxkd4FvpIgKv0NPwgAI+tP5g3Y
cbhQc22776Nv437ov+uYHEb7RQHuttmu5kITYhzcA6hYl2C/Nf3Ujuw1mnwl+/b//UeVABJYLRrd
+XyY1C0eB5WS/36sL2dB5e1uixA4M6hvJc1jxj+sICac+7dJ/pYvvegKnXN8JYjiYTn9tArlnrZ0
X3myxAjaWAuT4WMDzBdUeaRA6gfqFAn7qxUxqH077gNy8zIgQjX5BWfMKfDNfYSqWLnE7kgwG6iv
Sfv7ZogR3uAejofYqoguUDRmpxELxmW5liYvo1jJZZGkkcKlr2/W44kPHcondQnHl1PlF0b8nEYT
vLe4AHHoNZ0JkRudP0YkWhjBK40IpJn2MAhmALAgTmGTGGXlvGKXMPXGB50qWaajTN2xj3so7XKt
7x4pmdTwvZ6djQz34Nmaz6YpM+NNTwrh0O8VxtK8cwsZgZETZYiWcFXPggVSEtT6HerVQtwjRXo9
UAajoujKSos3jgrYCUkykGJVnu6XbD8Y9t1x3pA8c1oFZVi6HPoK1I3qa7/U8D1BEq50pMEJLrn7
eUsliw3EOLtcGtqDY4uoiPQFuSXlY8/c0HErN+2dvEI+FwJDAWIYYyzjkFJLB+P/HesCYIVUwrz+
HIZVPnOFYpFoeWyRwElP2HURUhTa0b71zmsjHpl1ZlkVM0VKQRymfy4K6+56Jeb7Yjdy9oVxhXi8
P1w6+zRnpnjCBHDWytpLxNmu5SXaoBujGNQKjKWgXSvRjeBEyt03RaRV1UTZ3KzlwT85s5VjdTE2
ZC5AXKmz87ohP8x5sPs/9lOlt9rlC2mYQ24iof3qwH9g0rTl9j9QyvLBQulmdmOopAuOHWaNkPRq
8ZZBwzZeabl1c1CPGBPjY89MiS1nb+UvCfCkMVvZulXGwM09Qe9K9QvCoAf2PZJL1TAUq+WqU+Ad
8K7CtywuySEVKllq8m/rb3O2JwfSraKnQRc3GRt2WeM97GQce2kn2Mse7QvZqMUdKqCyKPboI8pu
BasXrrroXUdxB4jxT/29WPjzfenvXGgs5ocmHEBi4qV9CJ1vAS1GiDXDSlhbgVbPcA/NclOdDcCx
tYQh8WHlOBpgcMTzZL5nEsc5wz2t4CyaBsDjccCgLqxtpgJrK35MgEWZFb4A8KW0sCCHe95Vb5b4
Nr1MuHlNI/DyC9jXXAUjEj3bDrmQnx6IGhYLiU2K0rykSkqkuPVu+mozB3U0OJu2sn1yFFLrhQAC
KIu0e0eV+dKONTpBL+yuMwccMnTMRGe69v3scwWe/EivOS9cH6JX9wc0F7U9U290hgFzKxvnEjFh
14buk0WiOUOyLgCa1HbnXsu0kJ8KSZbMK4findQtqdk1riuqrq5UDjqd5nz/izmhQltHYA5w/wDY
C09rWU14puxygMeiMDPQK35UJsQ8sEpRET1JAw6j25t3q+JeJ5BtoT/t4J43vgcGf5uQg3g/6mPt
RrO2uSF6tcjcTGnx7ET5fXR6FSvF5teJDyHundzlBRZI9NwqKuUKrIXQ+Zda6vBsa8OtBJr6FjaW
7vZ0T/o0sxy5lbjPiObOFrnwYF+5pZO0YZC6NwTncbf8s33uBG6eZScxyu8PQ9h7p7bv2sryjlUX
3vrO0g3LGUM3+wDZ7zGX65NVJD1x5zCnLckqb/mPO8pbe8iTWJ7UUOldK1CiIOWzdxaVx0S8rhUL
j7ijE8eyD1lQsesxgj1cWRU1O3oW2v2vm7JS5AlKSLXzv6XkS+hpiX27M7xx3B7kAypm16fNRH1p
NjJI8vPHf+FIE0va7r7eFRxsd3AOQ7cP6Tyo90ajvGcOFUA1BZ9n91jkqudZ8lTgA04JoiMsgQLO
tfqqTTYTYxkjGDH1OXhheJOrJBUquasipDVUnuZSxpsbiTNfXhDHgIxv9qS3TMHvozqlCYZrbweK
4eI8ovEfo/iNK8KOWXnuDMjQun54nrZbSpmwYv/x+A73OitiuKVKNagflOETjNjAOZhn+4rVB/CE
Vi+q5vhbyKsakuVhXB3heyiD1P8SUdcPGdra8EKT3jgQxUX8Ii8yeDMjn1mrleygKC+K3TTeiqW7
S0xvVQVUR97xZG6Ef679RwJyhcPZYiaeCiuvx4/eP0IRgG8JEUpSaeTKcwhnFRu/ZH5CpApScEd1
3n+7U4rUYdn8LXRYUSgKsNtiJ7wU3zgRsw+r/Bzz2oIaXu5fbiybVr7CqFvunm0oTibsDx/zSVMM
OBaVw4Um3VLtm3/wn7E65xKu2ZnwqWXGYd3bcycrcIMLo4OfNlXhZkfDO+aAuBzBSVitN9DY1JA/
bs/2zVOYOEdfY1Ir3TpXb45HfGzWnSiyJzbtaIQBTQ4TU7uIZ0JswsncjMUL6X6kQqbaKTDYoh0A
UNKMUQaIr+dG/ysoqo65xmKNh+dfGBdD72AExHiL2BwyNJmxc8SWwqDrx9i88Mdt2Dxxd3vQY6Dh
UD/B7U0PBQLy7ALPaVDqDeRQstcYEjUcVGnsgw5HfD2uIjtNUv8o4ff0Ne2MELoqIPa9rLMGrg7g
TUbRxf8LANCs3mLO0ZgWQwrFheMbEa+AoQPaDbFO/fxvAg0eQZltJhSCC+LRFo7tmoBf7JGpGvsD
TXsBg0iJj5yppjl+LUDKfr4IhM6t8vDmILd02ylclQlpRknKYKgZb0yEGM7yI5wd+Ylz9hboEfE1
cb/u+MhfQnwkTfIRhJkHdRKegba038khq2R7ndkXWPkxzWYbwkmKjkV6cUH+JRHajPThl8IMfTSm
n+Qd8dpU+LGo4PUGHAgu5SKjBkbq+WCeWKnVIgeCVm2UlLOFMCmWBPQCGT8g2lPp4xHWm0u7paDA
Wz99delj/tNHHxYJWdz+hufzMgzgyUaF9fDUC0hlyovbf5pZVo05TYJfXklrlkrK5IiJwcyz3pNO
2Vc0bBTqhUaAfAhvZS7Mb9NH7CmNIFIi2ORLcgS3hqnJDafi3mzn981jlX73AjXSG+YxHzk8hJrV
N4W23jvFeWcWbPORmM/kMHxqgtF4M+P+R1zB9HSS1TkVoVhv71tF/20yOKINWi3EXUdVSltkLKkO
MztZYQfOA915v4jqiTYRYebuui5vUmwXnKq1JU64jBPpquhdSjcV2CjzeVymD1AqHPdzBwa7doqB
wFtBPdO0Rz24N70hFNI4l15Ng4tlTSFmbKFZgLeav2l7tcAgZGPF9moXyTrpmKBX6UY5H3M7gxlU
sG5s54gExfe45P2QN+Nlf3OKAfNVDEB6nQJz1DD6h7FN/jwICVuDwOpWikn7mZOK3ku0bdJH1Fvn
1sX0Tku4O3kOTkNK7iPITpHfs1jyS+Q5cNo//fXD5OnLH7yIujhR7cng9WGxdRKMj8KADKsmmkJn
T+h3YX7/liKca5qVg7M3aLkUBYNDH+vDBrkoFVnP5BmQOhUkKFH6J1rHB2chAWreO0oSX9RDUTBV
K9l4dC++4hxvYnkKlown+6GGme0D5G/y/nsUfYK+GQ2sMt62o1XAk92lS+PArteQJt25I5oshb9T
2BLXiN9RDRsTwWk/9mPbNcAXQ0vu9SVdxscXiy6dDBumBXMqYGVbAsWN+WF54w8eqo9jdjJcQQPF
vJKm3kxi5TnJoGCbikWFbamBr32zuSf2BInqZ0SAmhFV4lPE5Q/CgDiJlyBy4Lep8LPdMZ8/yPem
n8OrUvAai6vO91vYb9TI9HrL1fbJ5mUkeXy9RLFm7yfXSZZiiFTgh+4Df5IXFcMJesaa1hu24cUH
APGMnsfdmycDbByskfptiZOe6SIQES7lzSzIjlHkXuepi9ztP/5SY1h/89DfXE66VQ/xDAQ2osrh
Fav/2GIwtnivTSQD+Js91hMp3Tr6dkkCVEKHmXpcDoSBQ3NCYfmT6dpT9lkJB8iCRljE1maCHKe7
L1fHCKgVPRzxKKOhjwXEmfVTK82LcgwVr0mGEIFAtPai4YB+PpPM7gctJ+F+olfv/EhxEwzYzrrV
WMKRqKwlGno/L9/ser5o/NTKv1/mzMn1Bp3oQD7hRp0/0DBYoUTjU7xjCgsHT043YfRPNU9B7OwB
fbk9nlha6q4fozuZ+ZLbBletPYsDPsmGY1ksj6EE+tTWUiBItFULcF9Dh+1wNHq85TQ2yDOAAkAo
zuIIO3RwS25m9R385gKEd525+R+JAZE6CoE2BYP9Y7cZTo4swwPpRQay6cDFj33Ks/RNYuvx5fW/
VAaK6Xqb4VtK2pBuohS4TOe1WfqnsQ2UPvqjBfkbLJonPHIfTpKJIWILB7/yr7vj5BHw5JT5ue3E
AOkINC8NHo1HRYCh4gjWcfCDJpvdrL4uvg0zX1E1NkTKtGcnStTKgff6niO2hDRwK03ES6911wQg
TDgtUCgHJMU31R6WGZBEICmjJAagUrt9ydVPdP0cAA6YM1M8eaCGfgY/rzjjqxk6ud3QUEF9aRPn
6QuoMbig5t9kBgc4wuAlF4BbBEqKpiS+lsSMzuDk1eisb+EeTNYGDavoO/P3DXDxGhq858F9vITc
t2cjRcD8hu2KGf+MDiVmJ6VokuGXOKW+dY/7lMa/KpB8yi3DFBrP8E+nI4QusFmO31fYJbDxSb+u
22pGRlWjBhYjI754r0ZmZx5FL2vWmMIWmr/rUYKXHvRkAA2gCuGiMCDoOUE9PQaEfX33uXSZLT2h
1AGAl5My0cozcEfLdYFrgpAmZQNtn2Hwb2w5qdVJ8NEoVnjshPl2ijOzNjfkTPRb9Q3sW5vG/+CJ
Fl2nOLVL9nmE4v88yEY8EP/PEjQaO5qM4VpSIsXcofk+BEbrC2VtJl8TEfOnS4I4R0gEZbpyv3/I
Y/4YtfJvuby0FjNX8VVkueN4qtne0F3KbD2y1r0WMR9ylQ6WonDDu4GsOYDyO+WKpI3gwGhMDOeF
jLK4dTXBNBn+azQ/SX6uRzqhsiM3S3cNeG6f0FgESGmCqvfg2LsO9cXShXOHu/t9fUEX9h+59UWu
99RWmWxH1SFGMySVh7ntdtXq989S6hS/mkZkU8CzuRUltniJXb6PDGncPDGUuDxfb2q2JsQYNfeO
sLOUhpsDaTQZT2gTr5MM5JoQrWR2inbwDWoTRF/2HlUBRrXq8K/Zxe45EQL4PRXj7I7vPjVDys8n
7eL6JqiZ1o4N13e6oCEt1BfeHxXXuvDlVp/9aULOHDBp0GbRnPtSH1Dy44zA2ZY+sxQ1M93zk56A
rmo+ePz73NwYXyUndLipA2cpbRdVV8axrwIwLBZuJiF369YAadzfmRD6Dg62BQM6IofJhkCkLa56
IRi4eL+/IlNngjusYW28SZnE1dZhM72oTFF5iO7B3jdB5J3OLMJTrbqzCC+Q3UJCjOC6kumwEugX
D7icgUHTH0iM6ejFpM93mDc1Gclkl3OGt1U3QvLQxJjWz/kfkCIgVwu02UdVOsrC39a5ucwcYusc
KrbHCdi21KQMqvOmhLJZDTh5CRVYVT8yPdMANFWvWI5eTqQW6aVpR/1PadoV9CI81YKsq1bmY6TF
sdCG6id4OHec8QeePNnKCt/TgvOrFvY0PHElr86cECOusKDzHMWAg3Z1vW/1Qwgz0E0iZvgj14XJ
lHv8ZAR8qkzh1ZI1NX5y6lekMeV/Yb4jij/izELWCExGduhrOtA8uXXNGURhm4n4jTcxA27fgPqt
wdoE7CGBELiXi7g3ZZ8UzZtr75CuKA5D6B+DKKbEk0wblkZ8HfJIi4YpesyD67WNu5d/N+h2VMJM
teZmJxjHbAlrd56sFmrGCiVFLPMH1V7qHpmfqbvpGOx3AFk5o7D48uW/VPxy9yXunCb/B8uXkTj+
wi8F3wU5nRstPgZi7UozR33lxOF7GaDcb5e4McCyouYmsig1lskfUxi3d9kE7KE+aAxIF1p1uUv2
4u1l8RJCzkUtM26z9sgTUuvjr0BoyBuTZYExua2zSPTGi06R4bVGgY8qlsB8rnPJF0mHCLaWW/Ue
Y4ilgEioctUG25pDdliVbusApBCOjT/OcZBr2WNsEupfpdUtYzVNdEmehi9Ya2ChImid5TfwWffv
ZIjTlaz2/CiCub/lUOC8gbK9y+r5QutuSyil8RyWwRSXfJLbztcbbefsNkbwtXcpJsKl+8r+jjPR
Xoy1km8K9gMzVYZkenW+euS6owSmdyUl96UbTOiFF9RbBZ4gCGsCpelcYWg8zZJkJ4aPgbpA1YHu
4Lmpkt/5+2bl/Iy5qsyKA4F1/QkUdNbK2JiM85tbATTvz1JkZChBT30su5om0b5wert5ZsMcbh0V
5f/Fw36JHW050NBCpAuVfFqeuPh456ir5Fc8oN4UO0ZU+acyxh5o6HaVkIqpuRTEyKM6DTFQvb4l
auiQBszdoL+j1swmFyIGn1gaXX4PDJhaOC+SAbu275Kt4bi043aSSzeQxcR6bshyEXO67WGlYRx6
UKM5j5Y36Rr5C2fYAtDoGysDQ6OIEyyF4p66k/3WTm4cyWdF7oGRG9JyyJvMHIz8xOhfwsdOpkCz
cuXzNGdh9eSDmhC3vBpRwqOjGc/iSjEZazk5lKz1MuhzexWbYL6Rtf6aXtG7CEntersyHzj4ESZb
cKU5T+O/LSSk/PIVnL2wmnWEOO+rviHY4Oj3Psw5K68vnHUba5CunuJvirQhVM7RFVEgooxfB1yQ
VUmpfFk/UxHcnPdP0s0N3tcR9gC6Km6CjvIhbjzJ7rqrkLDXziRmQYHSdk0lWtJOiB4XEZnYoEvh
e6UnLlxOdh4+gPQgW56HOecOJlGdq+cblZArtAKICW2hSueyaoau2wew8jomQQxLlid75IrZjTZf
fBXQR6u2vvtc0H9CUQW/Cn+ebv7saziElLd1QA1SYXjhvGNMsxFZUj2lg66/Ni4U7JDhAvn3ZEZz
e5xbAU0b58IlvEebvCAAMFBWNpZyZkYtm1PDrNe347Br8prrHHP782WGalsd6wEWaGtomUMUhUYH
hgXyPaCXrK3iOTt+wIj9Pa0AFpXMdnibxcBAHmY9YfPH1cSJhdzcZqnesLlVoT+XhWCUFTWDLc9b
I3n/85bturPkkMWBrJ/0+xmBVycRItnY2Zg0HGxul8dRRMQNQl5EPcG5AcFQj77SKX3oG202qClS
7KK8r59GnYtv3DwxmUXaeszm3AVNATlWxQApOEYggAK9NafymF9HCefXeTnKNQNZEf4QKyTiZkIF
TEONGyNJxfj36/PTCPqRrbRSg9PrQV+n/OI83YOSrsqQ0ixZJh1bAUjcfpw8sl343Cu8U1a2+b5L
1aGFJqEGKgJEJIuK2Bd+PvAXa9AbojKO+WQrNpkknSHx1kUKbJij/FX/JWhODzLs64+IdRn7axzk
r4AZNlBPaRPIvKZ3d7lMQYFI1Pj8W/2eg/YUY5zVmIIH9dyV+n/CFao7VJflBhGWoP24P9KQoXvq
cmybfxUvlp00BSEkGmX5EcJ1XgZTnlLEoVg7qka8me5gENLLepogqgfP3vS8vEBJh0Aki/68Xoxr
NoXsVi08NaS5xSEYx/7LP2t3IJZh//HqjE7lqK6h9VHn87HlpjkKTZkdsBrp4OwroJiEG2MgGbBx
+GMfdp8smHjXDqYGr2r6H3wjua5lOTHyk62tJ4ocNEkAKZKkMNpxqyhNavtwkpn0Q46bJJ2oVO/t
ekV/ZNSD9KHdLLXIz0Sf/sCcQArF99IuJoSfKBCXDML4dd+6muSjOcW/cq8wGhPsLFCg2+8BkxMR
hCZYfC6GZHde4+2n8bgn6X77xokLWYTSl5+KywUEorwpQrl1ic/0YGrcLL51883R4JpGnXGOLT09
KShfiutQAww4IJNrEJsMBjW8eIuZUHwI3yMzA2iwWnYPpHD9wMky9c736nMEYMsN3aiJxI7GRWb4
HgZJD0t+yNDO7XRSb8lZWmLHVt3v65f3AZfh6u/1XHJLK6RzxxGOsfbMSBlcrOY7mT5RL4bOFPSY
jJWPkoTCeaCDDjp5VJxzBBjZtJKcWfOYTD+TzB1f+y06avJpsQD3Ejs1neAVZ0XwsfpoOvj2W5nt
w1Icz3VbUOiNUPQVfNo5A9w5I2CqkWyIFGljLqBoMEyelqKvF0zGF+DRI+Wl5DDmWU0CQ38SXDFn
J2+y7eQPAOyvQP4BEWj+/K1nzbNBqEANq30J9RMkfoLlVR6VVZiq10KhkwDUNHLqcTFyKmZHAn2t
9JoQyLIQaT5z8LHlgFb5sbJXiR32RiuA25hY0fiOOhzg6rcKk8RquIkw4HpxdwYsiG19llV3MbGv
A/k80N8L+c+1ScBNSTU/g+zae+YaAleaekRs1q1Kn83DXOb8drRv3twv7DdfxhzTPwL5bCWunJwj
Sz48RsEUIALIPf0r0rz2AoMiZxcgyIDzsSxlkBw/z3dMzhw63MHy6glTPaDWu6BDz/OUU60sE/SC
ino0vsLnNRhcF+fPre4myDYdfM7YyqWpl4PMT6oDA4hqDmA3LteFlzNV9E/ugLxC8w187b/Nj+1E
TixAjonuXgkagVvl3TlszS+PGwwHBoZnTHIutkCpM1H2hTU9lpvbkLw+49gfqFB+75LTGU+GCbPG
319rgnilzlkuSWH9cb8d0nqH9oXPSWzQ1S5w28pN421asbzmt6fTVqeMUfMi1XmSEYixXppp9x9a
XROsnR0sZLPwFD9ms9Xvg402DDjCUWsO9shqwgn4UKO+k4WR/dS+HXdd3c6FPj/aWVDPqi5syMVQ
BewRP0aQbjhWO5hHrJ6CFsjGbv3CDozAr64/OfJr0hfsidLS8K8ygaPXGagH9KWxO2ho/7uRoDVi
AF5dyIC5BzvbHFZtTbWmEc4T/mcCZvnCHQ3bY1TTiPUsoPnayvv6FlWW/ndIdVeTU09n0E2YLFrv
0Z5r/AQ25hRCXt3OkaPgcImjngZkIXLb1s6uh4vpokxY4gHWeQn4LAjcnEIMbq+ncCj7lDYukZCN
jwUUcZAVTH2JRXRYk/c5Xg6PIJz9Ki3DF5kZ1QptaQV0AjiD6jgAa5A3H+6anipPO1PeHGYnpYVA
wP8T00pADv4edTVpF0YgxUkTjJE5LWgI4nrOSK3vCV2NUFp/huA6X5GYL3by+zTee47lIjFdufTb
YYNYaAnsxr8aexlbCQhUE2pG6FW/bK9rSwEfI7n99cCq7bzzhnHRdUstHxjMz+0ah3wWyKX2Yyz5
mhPcNu6hXsUKMRNvT+1djD3x76vj9dUCRWQuwfbHNSDjdJDZSGuurLfB7uWnPEaS9EZOENVbqN7G
LA93bLyGtAIXHxYo1HscP4dNNn+01i5hww1/AJPrsZv5+xmLsWU7EboBnOwHLjYowTh29cC/Qq7i
3u+mZV8m6fi885gl0XNZtb6lSpgz8BYbf+jV8vD+dTwpqha2dngzNaOfmI69zlsntsqXo10kzvpX
+YCDefE8xv+GQBAZXjZRaYTp6xiy0ZPd8AJpAyz2orFIPuIbGwrcRKZvkjMzi4VavvO7drgieBwE
ktg1BloP5IN4ZQM59FhpIJrc0Sg3jvnlY8rFIpF2CwcZaAZFzoy3rCQHZNXIIDbMdUUR98dA8EE8
Gv2ioz7yiaBJF7z1ilocBA3lpFS3qVRAAwx6iCsCXncsw7UEVP+sfoMfECwIbERS1I0xME723Owx
uV+xhA3dFZG3VdlEHl8+0WHWycozk23YmWg1rADhW+CRfollRvCsiPpOZCHg8+1q4LzgvFsXYEb5
j4ZNqh+hM5MdGgJN1DgSefYBLtro3mRH82ALymdJ31g66aBmbFYUqxY6kI4B1bsPT4gATbDmn7i5
T0H/FK+kxMMbgb0yNFYWJanzggGocraZhqBDw7e3BQVb75sl2ZhEUvw/1Ev4nDNbAMhprO7dqlV7
lpQvrq2dCPuz9z2g0HO/JLYR9Ia4q5GlJoyNxu8BqEytlfYaAiBgNDMLtlbfvUQePg2OhBFu0xHh
ulpn60O3GMPFc1FrJWVYI/uOTT0uwSjJqsgRbB0jR1UUSdzBysHODXBdYTHLTbLst98Br21aMBUM
rndtPfNvYg9lVvp6WWtT6mQMWA8KOwdEj8tKlHcGTr1I5JoItoGsWpYP8F1OC+D/Dc9WzwX9augr
5Mnwjy/sOCqibv4jIEPh+lkzvwNDikQqlEDA4LTbarruA8gbyzFLxJthvCqmDhEurUWAY6K6Jf8u
j17NZeapCO2qw+4Mp8qkbE8z8hNcjDvaI0LrgiFxYM9oD2iD6CCUNYQZJ2cDCnsoPda6Nrvf2Pot
TX0ITykBxl17wPC+ce4NSod7/XZkcCf1XUt/FIqhoN1/sW4pH963AtvHnPckf2HNdk6CF2Wt2Scw
U3RGlh1ppm2+8TF/pAA+aRlXKATX7mNFjZQrgXI8bqlH2uWRjNEofvMWZQSou34iKE4ZzoVJfctQ
8QMBV4tO8lwKo/B4fWKYVEhaim6PcxgYjyvIh81PFgXFYu3DpZd76VBm7Q+jVWq1ap9uQ8NY4hFX
7Ji2IUpZ/Z0wBZLVJnkid+eWY/kplmvmzXls25SkCoOARwGuCOyWrkPKjuETy7QHafP/67x8mpR5
vJcB52I+RXRAAWkvs5pV9TcjZOkR95OdH+IaFROCF1ztM4GPSUwQJPxaY862rEZgdD50Kq9EYdLj
vJN/N5wE5RDDqI5cXV2moHYF1Ia2be1t0pTZDmZJ/brtWc22CBjXCtxEX99gGZxsEVVIh7wBQnNI
6GbFNAR1g3nzfchttWVY/Fjgnct1lHvoR6We1qJAcJ2FhXvsjZtGFKRGIK9mlZj1TJBk/Dj3ucRC
Ml5/cxCplXMgOMTOeCdlDghp9koWXPpvdIQUOFgfJ3EQSWy1ZgByp5UV+iUNM0hqJK8c06L/MsNc
0Fk8r0uLzFN5oWaV++NQG8L5rprJ3h9+MBZ/d1yEdSF05S9fCzYt/k5aR/403S/pdO04axmmMxbR
UHbN0MUgU7JCQuZ12ZN/KNUP0JjV6ta5L0Eo2F4wiXgtdeHb6h5IrGRjuMVVoketK05yhU+I77Od
tC0NRkudEsqDXZDAQa0Q61lGWtelr3//RIyLh4e64kL4xRIoiYLmR6OiSZpp4RCvw9FUjge8O+J8
KEXjOBuG4xMqLn17Fbs9iCgnYYxhJOonBnZug45mTr5G18YLApmEzP7xobTWvV5BZWLhQyeSuGRS
lT1YwK3SZuUDCfQlFanyRvuhYgzcNMmMdPJH51+GQq1gF7pI/VEtHm6o4ZoiuhVy9AEn1eCGdOFr
sK3Lo7UyhK9PqKlO7hjbglU86ApG3xwaLQfMaMYq/GMFgiOuqHb9C39plpQhB4KBcd2izvrsuu+D
Q31nly6IUTZDoUxFplp7Emq569wbElRavsMNdcBFUyHA+RsQVo3qQnQ9sjIf0AsB5EK6VNtZELUU
vd2pJPyfDu62REhfbmilne9DoalF8gyWl0DcsZAmJj6jsQ+Eh4OoOa9QaWcmmLFZicNDqHXp4Xg2
WbXiyQvrj3wgwT+eG7JOUcwSGOAMQVmJ31ovlN1SA9UbiVvinmbHAfY25SR9s5C81oeOgyJRV4p1
7EnoSYDEg4V3J0KPZqVRZ/0pmnWp/O9m7dg83FuiFnFUZTnihkKMwRGExeno3yszm7Gv1ZMQF8Bd
YMaYB4AYCjXVOsr8Ug0jLhoAm+UXIK+N0eufeXTGWrQ60wjyzYwzTGm/SOhzOEA8yrYvttgYOHS9
XvH6TsGNiA0oHryksZj+MyIaqBINY7VLaVWt1K/SarmvyyiPND9FN2R/zXT7mIgGwsjLvSf1jfDI
c+G2HsnZ01bFCKEQuFlMVkNHCJY3DSU0aVKaSagJw1H/NUQLEYLjKdeBGlJDsKC8XQbhKMfHwqNM
c1Na6MCVmlaHWiFl+VSrUt+10hMTPmyAsjuR1sLrcn2OVd6O9j59K8n8PwlnFQQ8ykn8wxweWnaZ
zc1WZdjM5N+ehf2QIiXyq67JHYxNz6qq/a/2xUXqlXo+Rp5fpg/mLFykhGHt7RRbdVVFkFHVyLVE
fJEoe57+FTqlIho87IGD4CCio649BNqMfBiC23FO1vfRwQph5fYcjHz50pPJq9QVXTObhyw9LpkY
i570rg7E6Ac5z1oA2QkR/ZhRaTYXMRLPh93Laci2EdDGqGtsXWwrthbo6HVHaEGRFxtOhDHMWh49
1icKcV8xp1ixYDJE2RUNPvQDx4xg2et1ng4aPImh6y1bv79csZAWsV9V1lphL/wmTI6T9NjXYolZ
klKUv7wd1+CpTUihHh47xvmeHLBK9IGQE+WfmHJdy+R+a8uNR+o2J/3QmrWzb1t+coryF+r+DVh+
4VFHH4yqfQ7hEJf4YhTDe8abU1Af1+t04G5N8I+lvK34MFeO28rHL96O1FwN9hBj5BeJN4YnN7Q1
aWMH56jg/VFQsSJeiRCNG4ssP1hUjRxwqPjoPeg5uZhdHRi+FTcTwRR8cp4wH3/hLN1V/jOxz0Ra
GM0YEVetCeLSPYZQgZnB5eg+35lUBURsZ18ExWjwI7XtC/ewfX32dsGmPcwjHSZYGNI1kiUui+A2
K3xVSTQODUgxl6Vvq1z8MnJhZAS3ixLBHtJq8W+YSvC+b+OygL0yhld3gjXN/1g1bNqrdLbOznj+
Wlpz5kY3GFD/DyvAPD4DJif3MNt3wBbPFGO8hVLMnuVhXdBkVL+criHW/fDeiSrjee6QVH45S5VR
e2wnCLLiI/ToKHjuRIfiNsZfC4eWmI0n6CU6UPgXQq57HFC7h+tGGEjKTBWaqDzKpeXXmMGh4spO
DcpLvsatTLUCSHBjBJhax1Ni7STcZgHqlLajD7pT2S9Cmp5ByFhDzO8cLt9w3RL2uFEegyOVmQxI
nS/pFK1jL4Mnh0/My5BpSkFC/xdVi5vrVGeMB2QFgSmchjRgEHYX8jMNFjA8criYfPfdjJLkq9Ys
Ed4Zk+/wQkonTWRmhOWvOYGjmDqVn6MH4v8wdigjtQst0KZGRn1RXvgCUAj/8MBPmznNIKYrYlo2
YEpLd2hqQT8M7GDU5jKCi6a5qkMzVHhl5MLsWmW8EKcgPUQ3w4jZ0dEqkX0JUF1UlgswSyAtCoo7
O7cmphD8oh+t9AV/C7WFnvptrpBoKJ2McJbpGGE1iY/x2Dk2/ON95ZmZAxra78nYq6PbvT67aHOi
x85Tw5d4DEzz7eXRpxCx2uT+fMwOzI+nKpCH5y/ZdsvmwOSw2fhJeaYK83kuH7nKODuma9B5C2Yt
H1xdtPM2i+ExlCzlrvufsDKoM0FGu/xdw1XES9PReDOjRsgtaY3jaG2AYJw84LKJYDT2NhBEgsml
9p+Xt6hjlvG+ETOJ4zXIkF1Pfegi+qjiTQY5W442MdqJ5lDyzrf94dtSabAjTvU7nGbHRucIoffj
iy4brZjUJPFUrjGjOuQXgiNY6FaT4P5bqgOGH4C//sktfTPq8vkHnkMBbww4mBsbbsnjKp7e0bpg
pGIuL8h3v9QWLMyJKJpGg3gvJdAR+wT13fhe+tjZcB5WH9s2LvLCmz8bIkNq8TIAuJgQ8w9hyCfQ
dkUPvcKcHYHXHlN6904mpL4WSx2u/KZyDQA/nACNA42IzOG8cdIQeM0+aNX2K6ldTMVjN/QmJ/DN
E00xPRxjL6oGV5TIRSOxtSITbZVLjGUK5fL9UkqBgygJjauz7B1iBF8LrkEZqW+1bPJetynTxw4H
Qhbv3rqlkPQR3euG7R91dn8YxpNWN/MgrXoYlShk7KRzf4JTPw9r6jp87bDVZmc+MpIOk0NRQnqP
KWicSxzhwbBg2Z4NhldkyxA77jmiOOlSSTMuijMFMI9gIWaHgYlGKlNwmhRqyVOE0VoBtU5T5aJk
akJIdXazxZbVX0yy0UfCsMR02aAlH6vahoXcbxrQKPM80lSy6NkiH9UqoYpZ4o85MbjZCdWyqeAD
mDUT0ikWGSxCqvfs3L3mkoMsKYj8Fn6vc0NfXjXLfx9NRLggKWjq0qXIgAHX7OMynzGayOzYMyDP
8M5M6xzaxb243RKlDbk8z0KyR8FrF3efJZRglYJ67XNHhlAWjXO1Pj/8V2hUHm0unjgEE3ZCowf8
Y03b4FDGD8r/+j7LdK3IIYYK+k3T+Hy/DEDWuMLdYovUEsAHHd2E3J4emUmEb/kLEae+eJXTz71Y
xYlddE8Tk98XIDzQBirkDt9YiLMXQGjCYluaT2OXKXf4sNvVq8Z6/Z7vZkoIg23BSflTUQI+d4un
dv+EPkYVj1txJFzzgZS6uj3DIsSqU7I2yxY3zUcz/dxKVbHvp4T2U3Kl/CbWbJDMhNV0qWULeSeK
YUxOyjopcjthIZbmvtNWUOns8+oOZXNnHAUeX3z60gm1XlpvcF8+o/JSHvnYFejyRsr/F5itX/FP
E1GM53QpXUlOm4ZjnDdJ7D2K/4mol84taE35elKdnGSN/8HbuUuNmXAatdmmuCbAGM/VSRCoOKIw
O+lvIFAT18jTnV+FOiTH2j0tcxzr7ZUeWETPERhp0ftC4wnJyPFq0G+I9gRtfBOljWradww5qMRG
jR0up2u8PtpdZrmtKD1jvtY0+bmMci9S30Z8y0D3wMpdqgq1M5ZJLofWKUmfvLs2H/sJTm2RlUr8
cDDxwBCOnDZK3J7vfxUS7TkKbv4a/+25D6iicoBeSzEVknaYNhNhI1bILoYXpe9q8Z7Uv4nmA9SI
QZax96dwcnv0SdFn+ZyDZdnIoh3XQO6v17lRx+XvklrxpAt2pRN2hGBMv6E7N/NRm1ZjHEpJ7y6P
onFTFks2kBFhttffjczkpC6CjB1FqKxrKd/jOGuI7fRSGvQProI+tnJF96DhWCTj/xliExnlUFdN
Gl8qKB+9NO8c7HfHjcQETGmhuJKUXqF4VB00pI23dNkhg8c8dg/ROj54L0AToOj0rZPzovk4D2uq
l660kfYa6Jinir75J7KIED/Vxsh22guzoq6dYfrtINlU7InbWi0zRRcl3K1rmKa2E+ULZLIS/Rk+
wZXFjddDUymvcFjUDJCTAaK99gKc1JRYPjRbF72ROej8F9NPLT5qDkpI+BAPgXDVayWQsfc3pyxz
E3x2wReB7+zxYqsZ2fxnJbaRCb3l3tWCSpa/EvjshKN9Gc2MvJszQlqIVGEH6R1BkKp5cpa0Ywdf
4Oas11zZCtBWH+iO/j7U3Rv32K6p7rF/w5/jqgU5JidzoqSqQwXIkKLAS/fw5sKoMy3V92XTxjWb
4Ai0CUaivxHwndU8DB50XKFJCCzzyXxwS4Iw8+CFD8WC7aJ3H2xUml7Ey62229eaANIU77p2mSVq
4mNTlAgkcccS0kxSdMiHNOpyBpcoeKSo7d32/KI+Fv8M/XH8ychY2NF9cHIiR+x9Ij8ZebGeuqeH
CwdUkKMZQNbK4S04qKYM8wPtilEMRUpuKniDCHeIDfxnJgvTNLdLI3thyDOinQBoEBUBubWUe7bw
1pTUTTiwl+zvbbuK2WYRiOl20Zk5Sx6V6BkVPgqI5C2Ovcctd2iSu19CrogSbJ9Dg5s44s/uo/kQ
NaXYcqC8+8MYn5ZUe2fXk9oRR3Q+tKq8vza+SQaaytp7zLvJ2Cww9NG3IfEe+MDz4D325J02qx54
P2unhlD6m9gFOe1nz0gORGst2v+34gZrg2gPzyZ+24dpZMePKIvVGJivsVe+z85b/TJneQpqHTHd
LgXnq9/ER/XvvOlk5y9NmVWQW4zMKIXsR1wYI6mqZOYq+IIIqa1ydndRAG394Rd4fvuVZ1khmJQg
duM097bKTaE4lOVhKRDZDm46tlBf0lQHIRCAP+NTIHpqAFyMaxkOiEAZYovpKgwpVl8pvowklcdv
sQ3gdkRgVDM/e/lyISRivid2e1VKFr230safkrB4oeeXneFPjfLt9/Pyt8oSPu2k/OpvkbxbfZVU
sM123YKoztfhs2dpRelsuMZLuFIJgMhUv85BHnYneBz7VvX8ujDYXgYjW9cvRZQeCiVJYCM5I8zn
h86O+ETAQjb20rV/ZA72j9Pug17u62zxll52C2QwIQZSkNY8wsqyjv9avP/jTyIlxF/PrJcBgWM2
tlHbn/bWGJX6eBACbneumYe5OwhoIt3zojOqJEKE55uc+tn7gGihOvMP0hMvZkeZp0bjMZ5FyHFI
6zhjmZrTQQIc7Ea/6LxK2/Z3IH/DOIRWQUj//wnMlKU0+0xBZF5F7NtDAtScX7LQWBadFPKORwnz
ihMzODe+9MJhfPEDZ5VDISWnAILiywBcOyc5xxDl2GCdJvz/47B1lPmBJMZcZEtETgfOo823DX/7
vQY6rrsYGU/74i8idGCtIbGib/CDC/NsuvlA0YIJEM9Eid4/BkVrDxommCsDexoOZP1i/iWpFmR2
DR8sVPP/5WW76lIYrAGNSM91pLEMMF7RMQiHsawqz27A1WpyJQiKH8/MddxHndzrzE1IBzG3HfbH
JiIjaPGS/sV/bJEJhUfT0vCSwD+eqUminRNoFa6/ct4BZIcKfNGagMSWub5afMemReaE2tllqj/c
zuk+NGZJ4G975kt7LxifEZHg88DB6mSzyDBu3QMb8zJQmieP7NQZEO9Z41lQqImhwL3fZvoY1R4Z
kLF3jswD4wCtfdDbKau9HSI3f6X3r3b1FCVOqADXmm4rE7HHquMPoRhWa1ztO0eKCwmwRULkfZX7
SQJyuUB1gHScemsmY23XXRx/rK0TbewyOLYiQDwQyIlmqUQO6Sh3TuCzp9900C2N/MItlM+poFfn
FfHhukB6XyD9fWbGJht4Sl5OVN7HodgVikLpWoOFbLrcoFqjcVOIgzLWiybWCReHMApCquTJGbt4
/d4blO1WFHhKGln1hE/WmeGCtc1R8LHTOGx1G7QGWEM5XLc8GmfGbnTVFBOYVzA+1ovxpOqe5Uj3
DiLMDLK99OFGpxHf4rlWti+Jq6mJ4umcuVMRVWWsYCWbcq/tKJ1GeOkB2HE+jCYbCTx0SqiOw8tx
7VNWqfSlq45fTYFwA59RWtNWieNLzhAoeG70ojJCLd9j0+Y1TsNEMMGBIeMTaK0iZab2Vu93JNPW
DBzw5l1ubAnyhOFK6vo6jWlSA9yNxUUQiMNHDxFJIzC1KTAtovKz+59/1Y5TldZYFxUbKxDbRnul
D+ynZ2ELWEReY+RCtm2SmS6SjjSggq+4jqC2lCehShkfk2Jvu2k/apUej4uAAfTnEi8to4fqsq3/
pSILN69PGtMyy4QkfvNP5pvJRL4xLRu2LP5X7FHrt2BUh2S8FpFLK8tIxxe0mfLJTLru+N3u6yi1
HNfMfK4+DhD3XJEqruhc66qjDqb12oU4cp9+HtJpWFz6QZFXXai8QtCgXlcV82yVYIaYYapcHwiW
+fiSXab5rCSf+EgD/zb4AxHHCH01a7FEmgkC37zZ6oWPXfwsSYO+0gyc+35sjaa/Oe11KmBkmag8
QoMHZz/rGQlHRDqmXQt91+74eX3qlfdeErzrd0b/W6I1OM23af1C6f5vOWkxZQmBO91br0EBTu/q
Y5Lhp5c8riJ4kUxUsom4FK/iBRfwm28CFrwItSXjS7lX6Qw7CM+OA4RrvkBj3h27ByJmXizBtBfX
gNYIlHHNON0F2W59LJcp2ROMaDkyMC0uK3JGOutIXIb4QxMl6TkB3ZlKN5lfJpk7wYSE0rZaWoVp
n94DQQ0D2yPANQKyNnFHnVg8QAm+bIe3o4Fqt4XIrggbeZKVQtiroJU4VyBz+LIAv53upM9txl5J
Vhd9XtcuwuI9xfMsNir4jFFOXaDt0L/cBldAlKCBGzl7DYK+9P1V1T+TY3r3R1BN4Pm//2kIjSRr
YmALhsXfUoOJIscI0zZOZ8vuf+scgO/qITdFb4OeNXrdD4dDg2PQTugOj45H5/RhecbBOnNhdjNK
gbWHvTw8pFELumczFpPh39RXrEpDGetvSyOsD8Y2EP51dGkDgBS5I1fHpABXeoWXTreXkV1P1Ewc
z2n0o/f+nFRxRtq6kca5OljLXJLtUT+XxmzcnCUFJYzevgIFg9FuaYTpYccjlWDHkI7l8FFTRKH0
vvyl1380jA+/MWMsYaK/genpSNRwAtLYEeIXpcBJqgbnEDKUZiOOGnGWSgT9HVctiW5n/k/nXOcY
mjWZH2X6mCLkfENdBIFsnuHg1XIHUVechxSrwRCghAINEdBvKHIvEX1CYghKu4l2LYHXuJgifkB7
IJaVzCv7nxyEcuW/m0XJoFkxiSG8a+CSYJbLo560FrMor6clV8FOPk5FCCfkxV7Esiul6UimJMQz
rJjWko/+CER0qlFuSxNXCpGmVa1R3I68lCl6GwKp+8RbeO6p/xSvKH0gRFkIw/A3+KT2ZUmxT4Pj
gHw+FA4Hjy8wrlcKuJC7MeyHQ9XaQtIFNQiBD95z21AvUAXOshIzZiV3phYToFUMz4vgR4AZCRd0
dvFIisKyCpwaevV4TBZB4thID/yYCnfB0XlTl/QyDh4bevqbuAIQEF80oeTA1LZlD33GazwS+aSM
ixhnvWqJmu6v4+mHMaufUu7ikSBJsqV34ZD2NWMHvmH/+Zj8rsQUejrXkphMkU8yQZqv2jcve8re
4dlfGoTKZSOeXiWuEwHf0P3p1Qo17+bAhTAhwTFmEC6Up4qO6HpceWDz4LKeVjRV7iqq+wwV4v3r
m4GjPETxgQcslUmTRdK2UvBo4F7y3phUP2Ji9lz1CVz0DbCwtnIx4dXddSKssMCiWuom23kgUSmC
aEjihufomRXtLsn2RyhWW9k6R2hJWMQD7UXz0z7BovE6KFt4yA5tpwEJ8vS7dIanogUviJm/MfsX
bV7Zun+9ARxMn80SIJDBkZaQrnqigwm/USlVbqrXs2K0a+cYwuQrky1QsK8A5eCLq9rqmOwElgbA
r5HBLUY6+8/TALid7KHutFdDLazMoYVSnNF1T9SGzlP9d5NkpjsB0XeMsrGt5tTG7l/XrEqZi2Jn
DhN7wy65RNv4uDLA+Ka+6bqpHQbYl2KW2BEA2FQSBX7tWNkfU9xS+zho7dmB2NnLQ70u6sv2Bgj3
0eA3XVFu0CHFmWrwXD9bm8pio4WgAm+i8jGkgpfB11le5hs3hbDQ+VyovulbPhbWCxh3+gZ0R4qp
tbYFu6vCzy21VAQM/IfTVaDw9HlLF0MSiwZdTP+lMKIjojGhJ2J/GRnQoYSpyMIC+1h93beq6r5v
ui3yFyq9RNHf4iTfGCrauaRSUc0uRTJ0uP/8xjeNmAXmL8ZacShnJ76whaOqF5zjJc9FMnMGic5w
Wy/fAd0nZwRwK7yloa25Z/m+0V33yEgKErdTR+yVHQ3pMZWH50O7WNo0Zp6iANAaBDMlpOfnCTj9
sJMVRX7R2k79frc6thGdaRPtPHSLCiAc7nfcRGKhf28aSrjCEGe5Tp0MT/N9spmuhwaw/Mhph5Hy
iKG55HLxwyiQZX6r+Ru2SF/BImsKAbmDNwXu7zCn33CMLlCfkkgQHngHi/fxB7iak1kyAcnDTNI2
T/oKEmsOja/e68vKjlEh0FpczYC8+k6AFd3i8aOm0EeRC6/G3zTxh4hY0RmRq/CWc3AZn5D31Vz0
dxdD47iYf0ptVNadYUpEkcYqeZ2QownrbE7XwykDOzISRbZoivjS7oHNkAQNFMyHcsLmJFCGWH82
tpLyi/OAoaWI5u33DP7m765M66r4jpN04DPoAX67EmzjuUbmHUGtHzQwZwoTNH8DHa57MDA8Fdg7
WDzu75jeSWsg1ogjlkdGqskLhAKllnLJI0u3NXU3BSXu9XkjZEoIZyiXs+WLZwkkdKNBdruZ2+WD
mNWLM0UhJFYcEl5h5jK6JpMIMHDSwJ2HrW8kepxw9t3RC+ontdc2Ap2dS2B9lX0Xz7ayBni+OgY/
NqqwsguZRJtlq3zSZXjhPSR3xn7nYO/pw32LNVKN7piG64XJ8oP7q1uiW16ZzlIRT1LtHlDnKpTt
8TFGmvd7g54NOkQcu4I+USBGwZFMdUsJE5FDLCXcRHGJkojCLRRk+wGT9C8e5ufVGH6KhAl3YkL5
m5oVGFeE/ot6kuPyvUcMRqAHBv+6wsx9v71cDoOW92y733+0dYEepMIjrkFR6hYi3vAcAYsi8s55
aPB+h+DYsSNwv4BbuX4YlzPke6nVO/VmrZ/FpsnYkAzl7blN4EXqR74aUNBzDelkOf9K5igTvTMV
VvKKFcpH0iOvjY8QkDITSzVUY1eh76Ds9q04FhG3JEcJNkCy6NEIzHj+GHcBihgU5T1wkgmuccBf
E8ymtBr3uMESwrFA/4HRduiLpTRG+BZvwuEyTA/wHDe40u8WNlgLdodwTo8zN+ESa/rBR0XNp3DF
qUaWETJxmLQW/QmiSBD38R1b/b4r4FIy5XpsZaONjxJk97gQGnJ2zhMnZZUo/+BoDpRWh4ZFlYLQ
hl0/qNhrhF1bC13tLB6tnjWpwTfVK8evg41TfszvSyTYJRCVqEbQONX6OOH9cFbk3DezqqPwLYRI
/cOwoK+klVWtFzm3Lphy7GTAerQgz3U7JW9eof5lm5U7FuZ8gdrRSruupP4wi6eZVVHq446YasRR
7ohqB2M+xhgBPnNRklZUUk64EEYd29+9d7M+ZwXvHh7vekJYlEFhgw0MlhIVOt3Upx346gE4ewNX
obMBjsIikZU1giBylPzJzP5JXP4bZxmSvS2ZHMs5y2oh16nuJFtQaLzY+gja64XmkcF7vlsQyVk1
EycLOwBm0R/9XCj2YOgF6KFYb6VHMNIsL1m03quqfawxnNwFb2RibAqTqU87GXypJsu5hfjBAL/h
jMu8Wo72laoZ8ZeO6xkulG+jGpslhtNlwlhBByCM5G01yUbpRqaWtrVoU0sT16fEcrevLoJNXpQh
DrUakzOfrL/CPy6cA/UkuvNXttYpjQ8cyfGIpcIZENtwMiLnJnYPgLsREu6n5MvpRgMVKqP/DTJF
7Sm+xsIsBuDnYBy/aivUAJqLjQdPtJwCip+dCw5VX9JARNqdb8SKAgNgV6QXt9Po4y1fj43+QWfc
gUE1YMI1Bk1PVubWuAERZV7DNVjeLmMmgI9RlV/Op+GjwViCOWXTIq07PP2SEc0s2bsYfdQv1tbA
BtHphKyO5mNrtwfjl3L9hIuGMqYAzl/mMQnz26GcteO7bnQyw4OgBJa4UP/Q9MHOSBqTaWxKT/Q6
tPXw7Aib8AlUMItLnLvi4Y3XkF5LMG1/EVFxJ21uYVvKGapHFtv8CK4KZsNw0pDsA6kZxS7/5iYu
B22d7yYllck6Y4kQVoM2gLvhltDHGWchwllv0C0DA+4q4MkyFL3nDChIMg795SeX4DLSAw8RIRtI
g67Ok3ioaPBk0vZc/z+430KhLylJ2gS6HMsPjW7B9nRURSHMR1ABmBPtaM6P+ZF/TY2Bul82LUNf
akWHSc05BmeusaEVdVh8boI+xONAfaGOwUNAHOyD61FLkoXUdKSQ0vQvOW0TQZYvxITbhXmN6DpD
dJi0+RM9Mv6cF4mnZjEYzaCcYkdaukNB1rYD0OVmi+nx4gkzIZ4HXRVwg100qLWI0RieCeYq6p5p
bEhG5Y4TzcAcQhK39MrfjCeOA/WY1iwJar2Qrz7IGZnlF2vGH7BS5VP4v2fehOfYeBO10YUIk0m+
WDJzxtEaiMzGUxRv31LHfl2YThHUP2dGMZ4hLN5bJhBaADSc9BMlgkSl2nFa7ac6XHni/j9ltFBF
K5uxI58sbrtTNV82mBW0c0lMa1oTFOewyq20/RrDNYAp7IBysGzs939ACOTQI0XD+VtSvz+95Y5j
Lj+7GIusaOtpP44F1f2x3aExk9WEG6O+O6KXSViPJZUSa5bkCZ3n1pXu8r0KvNRm6imVH2KJ62xs
bQaZHMI5D9jyiOfzIWQMOFFcUCcu/9aq4Jdo9HiGMzgCHscV4NDQze+qG1KwUNxERyMSHLWnhpab
lGFgyY1gok6idS6n0oCX/FMnpXCPJMXbvYKZGEkonpKDe+RRXbM8bfTX84rfsLVj7KtoWOlGtSyZ
dSkPKWpgwM6Pvx61y7wKdiltsXasrNJsPQ9LztOpTz7kqDY4OxRiwbS3bb1F3kwY1pQyZqsxTLbx
7vK8GLBb9AUfp35AkraKaOLhMJBU5NHcNJ+US8SRgwUE1lMb3Lus/5pLIN4cScQtLC9ZjFVrn6+K
crsgG9/YebQPoEkgVnDXthC5yfCb5oOSWAKOiN4v1qhRh25QCywXJbxmQgg9oklRCibGzWJS18f1
y9ST8oOXOZsm3C0y7Onr77kMAL18FcbQoJpPA41ak9Nnu1XYq380R1ivJfAQ3AaKK/BWahv5sLL5
YvAQBLyRNK6pZzIgeAAwhPGLO95JNv/vZOOi9V7Af8ZO77vYjEgEvm3yeRY8weiFM+tmz4OqAhva
DJ9GOGXdV9jNF9zTlTcCxDeWCqyF4AJwUuXYSqNzH95ewytuFa+hkedWd4DQmFO2QYOvCu3tMzSj
sNpeQTbEaCcUbdXKXpJc+odVkxWsuYTO7RamfTT/WeKKV12JRUK1nwnRSEpc3x3oOsHpNJN8a5VB
oKGpzRzqcJAasrjq4cce8rC5TI3fW7CBow9hm5TwgQaQfpOwIHyGMmjdPpnPJV+/zy12cGBqKErN
whFyFc6Vy4JvfNYjRVr6x/vAAQRui0kOBQOYCAsqV0LhkgG3S87F6/19t7Q6RrITM+DbypKbUl71
rZt0f4KlnEZYfQrosi0TIyZlbAPM7y6VLS+ZoZbpHiO8zALbC3lgKzlaqL9d2nHLwhjLbWMj0boI
uYQGjffnw1bYPf4i47P/rb2MvMcOW7idBQq7j6zGVpRzMjAkH8YUuIn++hZoazhqZ772orcb5Xz9
c+ft73PXU5SlRzMwuztpf1iXyB6dvLZQy4K6jmG1XbCDG4xe31DxCryQmVzHLt46JdNMVaDPqa8w
Abb8Z/g7GoKEg7RrYA4mdCIlIRyjrx+zAWUMTG/O5cCTvgm9bsopohlflq2/47F7Q7ZN/K1zas7b
JZ7ZWtiui43snanoO3NEO08smylj8xtTDmGbV571LO5nRWcamlmhmbVRTjOopk6H8MTLxQ3fSBOb
6Njx+cHnx5T/cLMnm2uY1kGEoIrn0HSXEzSaUoZXm35oPWT1zgeVPJT4s/1cG4b14DeIQEQ5YLRh
EzZcKFDtKlDCGRAW0+IQrOvZmpkXePNRuvO3RnPKeBOHYLKgVM7G9UAaLpL7Qz5l3OK8TOmbeBuI
vKiDPAIqw1n0Vu0ARypBilRMOAAJKbHrD8Wn01oY+3NTzohSTRHoOosTXAapH1cEzSFPyUBDsoAQ
0BamI5yWu2sNGaKPjBGm404/t3UH44VQaWo5OYGWdy+G8IH9+ymQAvvaRijeNM+WF2aNbrBuIxX3
KHdJS1jwy2NhokRdJit69lw3Cx5cWnhahvT6vc/wd9449YHdBE2nyreltEm6pkSlIuKL7i1CtJGh
YZzGjwOhlYEGMj2l/9RrtSWIiipquy89kozonzWfQ7fxGWlQlzKpWAXuj0IRQ184pee3Rsu+iuA4
/gtJ7THxdalpf0Xz71ehoqPnopLPpuSuTchOlPmktZsWvceL1zz5BRusXccb65bo4H+Y913QyxoU
TRt1WhgqgJ4dkJRts05Q74b23qYp+2HFtLf9q5ZN6SJ8IBqLckkdsmCiMwfN6/diIDA3s8ckE5Nm
pwG0+ieO5ff+2EJIClz6O35e9XbukGD8a64M4UTGSK0oUKtqY1mvpCdHobeb+xUYlub+XzSJNQ3f
YwHzxf5hOqezA/xlHTNKrE255QpWATwWGIuT00ke1yzVyEtn/LeVVLTWCfJDTYRu83dPnc1zKlgW
ra0dF0ObHH3Cr92lteXo7jTeuTCe75jLqmrkiVD1k8C8jqIdCJSLfagDz/40b1RjoxwslHnR7d8t
kTLqiYBypczDi0RObyIw/Yl4GT8ytK6yq23PJR2O2oikRHLvnDfCZcUyjJuy3RFEnvVRMo/mpnQI
M9WzgIS+HDTN+edCfoexU/iPOH4eRnNzoZWCQTCqI0Fw2fb92W5SbOysIaGjnwGXZOhHeB/yOUaF
JmVaGv8+q1HYofEfy79azMRoU8eXPtaXxVaFeOvg5ydnGxKKWd0KGgyMnK/luFp+b16P8+/f4mjx
aBA1iNhlw7XhpaBdwbJVPfMGAG9hWUjQJeY5ZE/W+M/HAEjZeYB0qf2gwPrNXrNjZjgajOfmoe12
xXOD/8opu8No50gI/j283FWrWAOrGnycuzvG8vOOZVJafXiRmy/P7rc6j/AFpvn1ngdmPDrQQVZN
2/3VCcaSfHR/7LuC7dzHduOgFEEZJ8Ne3WXCgNqzQYNCkQdzBquF4UIiHZSrV5jJEtXA8GNyf0KV
HIAtGng8afep+jZLeYhmJvur+PxoeZcsn+YcGZ07baHXpr8r/BMv5K/KLDXwoWk2Yk0zCgjRZhDW
WfiWLuF3s90fy5qtmFkd8x0/e2gEbLNq4Nd7TNtK7bWfWxLG7c3OKhw7f1zGzXAqWVc1CPbKCLLW
JrZL7eFg3P4zmjQ3R5x3lKR5iXu1Z8pf3BY0HBB3OLmVjJMU96RdL7u0QaP8BeQlCcoDO40BRXkC
MNvnkLzMGsb0xLe0pOhFbqCZvXcOklY4JWYGEiM1k1jhU2cX1qLJNULvhIZi1oezOi4uz33mgGIl
2k0NEYPVjXLZqtthWOAyvDZ5wVk5K9wnFiLnNzjv5T4segZ6Jv8+J+PqYZUb8r7Njlz2p6UWmuXy
xaoqX28HSQRu1KYNH8orwJtqPBzrVM7btHd7bv9X0JFXUDWfIsYegtjZNZ3VVtpJBt0MWY/bVSe4
OotB2ZefvkDJK2VeY04GKg9vx+baFKtrtJ8MTt8e9+wnnWvJ2ZxVWWq5BeAYBR5sv/HE1KVbince
c+JMUtWvqzBaskX+rIPX3Vy5IAwlkqA8Jixtbn6J4jPkvOfWArAluPt9A7wXo+B2lRl6pffEngsc
b0WEjshznIjhWxy2cKJc49dkqidzIK4PkrDM+HO3fOLCb2DY3mS8xMdHPgGT6n3tD24KabAlcUwt
oMkjWhPiEWwCacJX1w6aEEojivKmhXnPWLi/6qtZEKANWTPhFSQo3yMbFFBt7qHjrUApDF4JTH6m
0nLi6kbLsr7kfPgrAnzitaHZF5uqgThadwmu6u2G6V/gVTOXlFsSKcwvFf55JM7Eh3QISRZgFxgh
AydItq67tWVXW0NgukB8KOFW/MKmrJna3RtEdF/B6IPHvDoSlSLXp179UZIB9jlOHqKviOLbXfTy
VWVOQ7ZV45d8XfBw/Ap2IaIv7qZ9OmrlXLIpWl3Zx07Z6GjwwhjhFh5MoVoM2AW4hfxuZYNgKy7S
JaJDIeRD/9aq2oTeHkIiTGlmGD7RkqHjOWLrIi4BWB2mQcEekWlXyDYs+YaL3nZby1RtRlfLWpq6
mV8zoQGJYjRpvtp5EtDF3HdOpiy20Ck/5imjLAaiLfHO22WcH33vX9leNWWdVWHjd2Kvw4F8FbRE
gNnUc+Y28A109LERYP0ban6/LMRAowF2gfqqm67NKrhZ0l3CeKSDvn4c8MvzZGaGoEQuDOlFLtTn
7VDB3mJkCfuZgQSCPKV+wSuEe1YKo2BCsutXagLCIlujP1LYamLduSckhtEbanvVUz4Di3gTj1/J
RZl9xgJXpxG/VuXakrUhFVpG7iH9gB6saw6WuupjLgxBwbdP2dYu8ZmkwYtZki51/qlagEzMd6S/
C+IbkmqF0ulaNSP4IlrHqoTyDTWQnRyCwMUeqTz/gtb+DAvoUaJsJTrML9uRYfYwndRvgw7hUoiK
yetNJ3j2ITziDSAfnTsNvHAip9ogFJ3FitBhqqvXiZelq1jUFnE6xit7RigcP2HjgE3/t8lAG2Wt
74a871rhp/GP7deNgZG+veu7r2nEXiGwe8yQKX0kwcLJHIoRVFpAbI+dChKSdON0Dzb8lWwq+Jh/
VJOZBeum4H3WU9E7teu+7ZcUYqlXrFnyziDkQknbQLBXTof8l36DX/AI8Zll3geWeXyv98McDrkD
VBMunHhQ7ulGgM9iiFnMMJabC3W5R+IBXgpuyG98NZZkorRIPVPEGwN35AF6zJJCkXgbZ52jiNPm
FhToDafz8b82Gdkbd8BD9AacaOEa90Nka62N5Gahvb68pmbBGJyvp7BKPi9re6tz+6W7ZHMt9D/W
E3a8fY0hGmGVI7zd1wrDH80yUTE6eActutOQvc+IQnptv+XveuMdslZds0/I6KW1fs6mkAu7/80e
W4sbfQU6v/K8Hf1t9r8q7FAzZ3ByN0jSbNxyz7NWY4+pG51yOkTg6l4fHpP5MxovyQblDnuTY6CT
fve5MntNbK0CfeF3S+tqcDLFLkb/gKDJwDTbsMimEPIzhUlGcvPdwrBb4HMcCQvXspa8EGMlV+EL
IfoZmJCzpGn722qvSYLzy8MTOmrLAYP7j4NmcFPKb2EhSyeyXaRLU9dSo5xmcua6b/HjJHnOgNjX
1mwH2PF6pSUvn77A8HCkDVIWjveJn/lJXrHvcxiJgbEL0nYBfC28BoBJDdfVcfeooE+xsHTLuAOE
l0xu4aO5tviSKPWuVDdeYBa2GYHnUJJXd3T3SN/lXiVxtjaExS07q+mPAtP2KgRCmCjXJyWTG783
Lp/FmB88jPAkE6KRCbICTuibLTB5PBLn9ObcoyrWy5dzz+yKL4440NuX9z+Oah5JlNGsdEBn6jwh
QDs2+YNKmiiBFCLSTX1V51xU5cCXGN9hV+Fz9xcAD4UdMiH86+1yl1p4VWuT9rnlTZYWvlBS4jBl
FAWUdr4cPktRg6Tsy1/RK68uLEmPh+5577ous9k1eBnJCow7I/iTdfrF7ZGY5Ixfo/YVnGWnWrCv
0MsIC3ruqNavc4RElD/BpPBXD885PtnvAUKTiLRK1z5+rTv2zgzFtCfCGIo4pR8ND5coCb8hlkYF
njOrE6bzKnhTOoaKBDU2XQH31WS7/jG51B/NJdZ7DUMHMqTafTUJ4A+vANO7SWBHGYX5KKjNCcWS
Yyu8X7v1wBQzhohSJFHagRjiNLHfZ0EtUtbvL32EU9D9aF+UaXuHreZeB1ouamZBSPF9XGH6knRq
bL3oBZ5q+GTH5XNyZ6xloIV/UcnACvtbzcxOWQd9QNLg4qBt358croYU4sZuI/g1nRWwKDNfNdyy
gqc1xjaWuzPqU8FPlDqNruMcR5nafUKnmT1X/p8YPMUL29fDwxk9TbDbYkEJguyfxbqM3RnEC6G4
emGLwad5fVPoTpKpfsEJlT3YZBI5Uq39XMTobt6Tr8IgH5wJCYNCLm3mDYMbrQxQpz9XlQpRWryH
mqSoeh3aqQFBut491dhY05qQsEr6/iGBNyi54bXAdufv/u5qes6JnRWp5Xyo8l7QEZLTr2ie7NBt
McpVPG0CNBeba2zGzAPzubRZC6+KK2f6Hsz+71bZtk43XtQ8JX2oMuOzW8QWSDFf2AfAVD1TE5qa
KAR1ehiz45eDzRQlCMR95+npMfbND4oXMvzt6uWUgOLAeT+ai24UTE/b7jMmsAqVQUkbI/BlzQK9
R4+7vIaUu+jljNDqbtT354Z675kje3y2LvIoaULqIFELgc8gkO+j3/X+uh0caoo8stsT09psMVs/
ez1fSAjnPf7GxG9aC6KLeZAP73c0RGxjUzaCZSj4z3hUHa0giGxeXJeGDJoImJ7GXO0wQBSpPjr2
L7DTcUx7UjULikxt/82VdA6ogrTSlVSnPz9vw01oC5Ww7NF9m/FCbp0sEQiCc0ngNEeNk4HHYwFA
4D50hpZM9Aj3qiWgT2AfvVMYcaa/sBU+YL6ibE5nUDrgzSIJ4LSSOTD0HtiITs0apTY28/LRQ5xe
xZzWd1s/pIHYEm/vDWRXsl3bq8uNH9tNGAmZ+YB6zoaG1GF09JlinNyA1SHL6sFSYZhsRY1kQ1Pc
iT+Y3pwteqwPOvbxCnCLpNGhkZsi2WLJS4scfaxxuB1Bc62O35wNmVp/snpbmtb8OOagfBXa3mrj
qdcdwA9rOJrEYwoc4mrJ7xyPXOExXWzRCTXDyHh3yLWrZ04lPyBcDUoQJnKKIftarDT07S/LPqdQ
XYF73D+TXRDKqgO2qNsY1LNDIyavCjEMDK0X/6c7PdKslDfZ9k0ZMgZey8o7M1DRPqyd6Xd9Dmf+
4of4NyhBz76D0C1/Nn7eqJOJf1JUGBrWyzrT9VEmdCsAcaX70B1pSiud8Uo6vhCIH75iL81TCe9n
tU3VJvx230LZUk2Q0j8IuTzVoNOUZtcEWJmnUazvLciW65iUpW281gs2ty1/LM9tqunQpX1Tc1RY
Am0ER06tg05UejBS7tr86CVOJMy9GEhDWYeBkmOzBkSw9ZyA9WJSUk0QO4Ai2gQkb7Me9a6HIvfi
r2dfVhDYFD4+APKFPshVZ91f7JtsWCrdsagqSPzzLHK4dQ317TmVfoCjR+86V6Amv3DnWMBGi46H
biA+X5pBTvSAcSs46K0obtKiQO7ROrX8FgIKltTKmAZFw1drB1E2NWv1DZGuD7DArh7eFMY9hcIt
bru74YC16o845o8yYQSCzP0jl6wSFH9OLXUDfbySYUy9Bwt7GF15hfLTMCeh8B+/ASkDhz+i+nkR
yUhf5djc2GSubcQ0M9kDOhIN6jEXHOG4h64YN1Jk8BzQgJpk7T5T+7Pjb3ME1U/0maaYRUugVThi
8/tw2Oye2MjZMRo/exkcCRGRN4+pZqekbV4QOoYXsCtly4B93Ai+bTlNfJgjh4U7whtdPlf9lRvd
XFfD9NM7GnBHomKuZ2QG6lK2cyG1otE/+hYCYVoL45/rQEmUNeB9fFTCGeoAGrigNzpfy6YmCHUJ
uG+8wuqZeB4WUtl320dKGJrZ5Oyrj6Dc8UookxOpoFnC54CdgJKumGu5jh0jJ+Raf3NJ+9olwP1c
houPkjLoJHukWel5Mr49PORyCXeWjn8TayItJfVRwEhQ88BJHELQBkPpO6vE/jdCALInfvY2sBaD
G1yAKV0efa4kOXBleCIL/X3Ghq4H6E1C7k0LBpAGnhd6dQ3CSRxZnFLaCAbx55mK5ZSDakYR/Tkw
kxuthvj60f19IsXpVuF0Irq9g+X7qEw0BkMr4abN7SqoejRgrVd7aQnRCd14HswmRrm/VaJLk6Db
ti0foBaE9DcfQH3d2Q4LSwckqOaAOm93gnh9sgnSUtM2b+3v7f2vsKYhQR7Mg7fjmrfc9PPo+boc
6WYsNnW0mweGLs2S2jd498CtExmvMiOharuPXOZWMJkPh8HMgOq/tOb57ywjMfdWXSP3cvtmleM/
xvbgS0Ejna58Mp4pWTJatVSVzVG2VT/qEXRYZklDavJfb0Vvwm/waUxzu8zKlcfk//LTrgRDjzcs
FS8/kPYSB5L1lquzJI5B5+wu+F7IFbEIuNvwvnds40Lw4tzceV8hnOUih5IwSrNG7Mrwjs1lCNil
VQB+urCGR4V5QKwnxeK0P5ddpclUkAx8xjy7g4Q+DUelOa/SaeFa6VtWSts8C2qQSdpqH4u+JE+T
aH7DYsC6s8UFX+sOjhnkeWHPl2UYQ9fu1Zi41P007aeGNzMfuR60UhP/byuHkutC6fYigcT3WzP3
tdfNT2Ei7HE/cP/JPLyPg8A87bLqtH88qlS+3rAuyW2wlP0yHLdpD81W7Q+yiYJNWI30AC7sl7FE
C0XPAUO51eLJdShJhFHVfAQzxGofW9wz1RoxW2lWlV0MW/iu1q6z2e/bFw6OJCU/AFT6FzrByibD
3Tk5GaitlTvS+39I7rGlQVvZvqZWeRrgPWkmV3K2YrN6jkX6fjI8tCX1wGELSUvuPoI+eUFKU0xa
Y4RFeebPwPbhqSP0xP8q0VUWZi+mVW+/dB4yGAjkFH61XXY+yfYjh6M7iAo7Z6u0v4IITfr6i9PO
+i41vNeAy0eFugSiYLiB7dr5a2YBSplxMdLqchnK1SOqyQo6gBkdumg1tR33y4WtedNpEouVX6q6
TafNDrCPdpvtS04Vtadi5TTm0uy5HoA2x4y/ZdmUuUmJJcQPegWWnhjuQVZcUKR5l5H/H/fcEO9Q
CGfQwYFAysSQQXh0vQfZXJKceX08c6Xbe0SBAzPAN/tKPm9vfAoNGsx3tJnyythyuL67Q5MgtJpf
HRnENR8vV7npOhqNGKjXL48IZJkVasZ1mVW/9xgdFl8SS79CcmXkrqyrh0fWOF3Ux7GSjJXV3X12
2+nZ/wLBoTKmz4aQGO6ldqBCOczb3PHxiLjwOn/sE7cX73gQ7VBZ6eRbM7WD8ftfqYKX9wzs8LaQ
CIMpi520ZaYeklriTj24nCls+10up2DuG+8WCiUE4XdX3mldyrgqKzDF9IxsZyMkY/FR39A4QIr7
MCZNCfGjTUoR1mVgSYNJSXNckl2+fI5+qM80XQ0evqWnG/6NxT8TlTB6b6xYyTr2BXdGUyscRx+2
9yPiC8fEOn8An2kmN0eH8JzmM3SWlRR6gN1mdvTKB2PFRR46kpDSBkjS02hUEQEt941xl0SBDNYu
H5Sq7OekSbpay2We1J6LG49z1jSqeXqkUKAKosv/dk0x3Eer8m9AAx02wZsEeTxt2j0lOWqE96SQ
QclWMa2MAM8CYzqApAMnLPbR60tQk107iNS/WVMr45r7MFVKOKl3dDbwaeQVPffXnS5B6DcKJEbL
A1HyOGLgEjQFvNHvMwwPsZqfzyXzV4wAUBYFvBc8ym62vzvo0giyIHFNmTqXcYoj5EWhTWCgPjXy
Fv/Lk8t+gsbeJim1hHXfRVEDz0W7swEjLKozlN7FaW2hmfY4ndsYy5JBrz2U1LC4jVXoEY0DcKIO
Gr59oEWbN1/kM3pJXO+5n/QmEcdOxeFyU2u3uVrN9t5JxO37R1Dgd3aZbVqAEcPg459BPaj4+d1R
Ae4kHeJtXtJxCWfjJ/F9X+l3rO1mFYosqxyCuOS7YS9N47+iZlym5HRNbrMr7Gfhxo/D9DYgTCJp
iDOncgK2rBKh/XG/IRZytFypjhecPPNiY/o4MWWudIP1TezbDpa8RtgucDKcgRxbJrNDlW8UKYoL
fSl9BITt9w3MlXphNImpFmQcJ+mlNvNcsbsWiUW3UwIC61YjfD3VhHKQ+GK+xsI/OLJS7OOWLfY+
SZsPTq4Ffaf5Z/ZIl6WKWgoXp9Bf5fbsSANVYjRxX4Wqwk9y9MCT0gr8uHBE0kMZKFpJn8y03C1U
jM5N11RqJQwTPyQ1OBkBDSrzSx7eUc7Wq1fyCl96Tb9J5TYfkDRxhiYGxCkpAlI2zBkbSKGO+fhw
tjaAVAbK8IqJEZ2xcz/M+w4BdrMzQKsRYXgxRCu3y/gDWvaQ0VtZ8aJptjH+/ZTsMIg/KY2nfOU1
sXRo9KBjE3V6u/L7Z4+PPMYyNLvv0Q2ci3lfEji9qtt7gy56ec3PKGiVxCNld04uRfdfGGROKT5Q
UwWyTP0PArYvI8bhIsP0iZ3Bh+Y1qBvaOmTlpTEJgv3VLMefCNMjZtpOGlePHgURraqc6cI33mAR
PQkUvpKQSEfYSfyEIaMeSOqujzNTu/5+G2lMOudd4WZpqtW38a+HfPwjkKDz1D0Or6nItHIHlWfr
/5deYGrQr7FFA/iBGZ/4boQ/uNyYPF+kZYyD8029XJEI3PtYCM1YejEZUBUS7jdEBLNyUWLH9baD
u8vOxZAY/Qf++mOrDf96hhRJU54iXQrBHRYFF8cAhC6we8budz0DhWNzSIF18F9RvU8R+wYRlcw5
ybmJLInXaP0sRbHrZabSV9Zf+Ps8DKmwI2hWaNFJtpZuJ+CccgsrrAo8OEM3EV7IEDjSi081odUi
Ob5XV0BVGz/hxzCK+wpsEfmdqDw/yBT7VTkt59bg1X+xJk9GRRZ5UTKrbO0tU1lz5cQ/IIoQe2Zt
0808gqNB3NjX+ZkOWQOEQ8+H7fE2292RDz7Qahim3I0s+HkpH2c7xRSJrT43MimuXiHBWFogO84E
cXoHWmyy1e6EVIFNo9wEsgvZBhYEKynXYKbqCFDysshMDcJ1Y2eTtoVsKalwEMhowtTLyN9WdDt/
EgSRyFq0y8qx3zNVPIiIJ+pXdTLCum+rDW6kMKSODZzlSICg3sGnSVJIudqZT2Kj3OMvwY5h6x/b
BIDHDvazhiZQ5tN4Spl+/UB5nfvM0FBtKctEqgRCN7vL1spW0Hl/w4E48wVBdprHMGpPn6FWarui
R39jiVQO6KXMonHGanS4DHPWH7LcWkz6vdR1Fs9v/H4JOKpL3dy9FF7FXYs3VI1nH8oOC5ZPnhOQ
h3QDCX70oYXKJn0+pOS0bB+iSAgmMTh8fSRQqWkGGV7DEMuEdtTu+cqOlMejRyy/a7bGyQnrYvYH
MxhWmvsXPY3Z5NP/Yjy/M7TDF0Cf0HcjIzHd0lXyNSU6NDZPqSYqvc8FuDgL89sBPSZgkmdjvdAl
DvH5ELGocafIDVdX42XsbOrX75QKSE909On8wLozpVGhnh7Biq33zszyzTkWox9q5v797ZLx9c0w
2PMFJ0dJXAXSfq8KveoisJECm9cOlZmp5qK6p2imROGTdgM8moZ/C9idRgNKAKu/g+Zr0yi9AwnU
JrEM2p8z+rNKkEYIoNnZxjmuNp5Zyq7Ybm+n/O5LsuyMbtrgSsSD9LZiozfWXYQl8px/T+Ezhyol
4MntsG1wfJNZUS9zwiBqq5dcI7hptAwJhQIrLmGREdkG7Tl+4sGK5oZHg9eISX24zsbFupYd0Zk6
u8E6W24IaepVVXBQZ/WexsNM6qHsau+kA3iqWndmXuqkpNywWfIfbhpKFsHzZza64zrOJl4Ns//n
zwqVQRqIOcARxenlUZYBRtWasqAwh6wLOyzcywIJ0hJ08MBdWeXGyYQPrJuhA/4sgJSm4uacBF7K
eLfrylUfogs75e0tZboTntxo3TE6PEhbiziw0eNcNFn6BBmcw7Wvq6IrD0iIBAcZvcAVNQBkpzi4
ZGMQ09KoKFvdYwZ5I2yFE++hZD0hxnH078OGSrmGGh5zb4krI/qh1lxFsfkjM2v47BpxHoAQnlJX
VYKD7ildyaFFyf7mf9iqpHYoJOCj/306NUJyj7I2weKrhVpaD+xktQxCxDzGOPzi0HKW2bCg/Uup
eP5jhDP0S/aUtuN4wv1stjxyNgx0QuSSEIaDIkpF2c0uF6yy+kfX0omMuEhnp6XqGkY/r6sT0JDR
uAloozq29jDsycL9dD05o0Q7q8pGm8jG9feAaFaehNtMhTXPC5scTxsxbCLdReOpwzZ5lKGQt5Ej
fOAmRa52q6ZR/vrBa1YRehAHbFi4VatcSNb7WioYi57VdfAtWyVo7ZnMYOF29Ko+8q4+VePKw0g5
DQofEHOIslvYi6MsT0vviGNZjOWHiG6m6KP4InnRrwYtxzpikZjoZRMgKgPdfrp8zEdE/5yNv9Lq
6ofqpuwGmQjRGpX82aj6J9NlLJuIKgZqAOeuDvFiyRHYmUN6f1ho2c2vXLivX3JlnlCL1rK/VUiZ
R4TvAyAjbXh7hnST97T5wi+PzlcfrmHoAglaC/C/q7jaxDyMPEFZcBewEGm+4nUGLX48yu7uE2Z0
KYSbc6uM+HUG6ZYsG/Hvl5N2ejejpmieSW05XnrPT72n/BA/S12z+CMZkwUI1tpO/9SK5OrVqUH9
LYhXOXcxeQ3jScwO8kNONXKxDSSz8mDslhbTy/qEYKLtWww3rlrBZJ5o/xiRrKfflSyjcA0/zyzH
4SiSe7S+AOYRr+hfNN9ieCq7yWI7QDS48e95xfsDQ+Bxl2XWU2ixGCFGBPQG4cxUlEdu2NqOvHOd
IQlBUqa46EqkPNxmEOIe0ijBRLzMM5WgFjGh3Te83xO9iGQXHW3EFDOyPb5vafBaQXdGyeKPnYv6
KekAQrl5rxOxUgiVD6wPMWsAtId4M3rDHoYnN1hHk9+o2JBoDIb/NnexrUCjDCnV44ITo4CtRMGp
fMZQYd48OHZLvOTeiqFAtOTxJYcefK4lKJVC8cbgvACnr3xU2wqt1akBEwkzggfbIyCmi3bWd20x
guHGXWnOSOgpU9L+oVEDNj7RDxpF+6xf6xtQOiMlRlfuBHdrG/5KjleouMwoWQEnHD4CoMg8xknp
SCzxmG1cY+pckvmewLTOQgBgt02FkRt7GW/IRUHYvJDX8reztz7fbJ8mx8uoY67e9V4O+ghpURSF
DKQmcUNlJwJdtoHSWIX4VTnE/VrdHcl8gH+hn/DEJjD6aSDo9XOfzQaDDz+INaXR79QreDklFTr5
IU/zbR3P33Cik7k9eS0LFkrLDx62iDKPm6m/ETUgxNro8D1UFGDJOmGZCqq7yUJijhe82oIfY6rS
UxX4Fb+qsMbk2lcJEJyed5wxp669GelY7rvzBlTlGZOqGw1IC5crJQSJo/IjXEW2tRimJDW3div5
imxrT/Eo9dqBCDyxM046PQ1vPWm0eFDIDCmTSPR9AY9Uyb49VNbb04xRotMfXaO4XvY4rIbWBA4m
lRD56su9shIxgq8kwycfGFPDn+bMJSOJQ0BS6VANo+GAV40uO/yjDV4aj8EYwXIenb3xCgg/GFgO
Kx3PmwSA3Mw4GSyu3oS+FIfRNeMx7d6bqHg4IcmhoNUW99G1I7RCDeMo+tUMicY42jltziPjBfLz
2FYu5I2HXffHwP8OD/vWBDdQx9SICq1M5Ut9rZk/MYDqtiktFO2haP6BvdRpl5ZRNrFlYsqQlGxL
zzoVr4KMAKJRYSaif1fnp3u4AwcCOrJ/ZDQ0804yIo60Y4ldzusR7nwxBy0Yk80YvObNVp6JKSSw
DqZREhUvlWnzGqKpuS0tDOG6uYelUCrjmyQ/r7SZGsFqLtpoOW7LYEfzfNddJKRzzm4/2JP/lC1T
bW/9lHZMdxCHDMxWDAvcgX/T5NWvuY4iI4pOsfoLAvROP9py1p/nq4QsWukyI2/U76papbGYBGs6
fvYtcUJ0Zjj8N2EjgNas3Md88JUfy++IQZmbzET9i2EeK9tz5qJDaXKHlyP1cN3UYiScI0DfDwu7
N52VvcmlackZExxiBPZNP7yU9jN32HgaTa104Xrs7i+mz29nX8+SaFOWMmXGad9bjg4mgPoAEY15
Td8N1Gxvgskcx+DwCoqpnQQLbUdD2BUKmJs4shDl4ENIlJ/Fc3KXHlPGO7y/F0Juj1oT3svUfnSG
4CL070o6kl/Bb2py0i7j6qRG4U3OYCktDVucKUuPCTC7KbDlKWnr243oCdre2DxeHEpYB7X5m7/3
A/PvCANcKthAgIjtKGBIaLQXLY1B89qlsyk/TjZoAgr0t/Z1xIN3uvQshrXYQcDQ5YxJmpg+ixXo
OzCFCe14XEE+a+Dxy8tvH1N2UNPqkeRm6fzauWqidQPD5nAr3o9JYPnIktT9/A/z31EXH1qzUPZ0
y5xn6B6wg7feyxcjgtGgifI5KoMdFQ5C0BltK50aAAK+CKOfObOHl8gekRWrD+Z3bYXcKguJ29Mt
nLfnNu8QiWcmr54kgtagUEmpZ6WB9ao7Qo2yTPBaisf6XkgBJasR4/CgwXALQqrdYhJ46BGGdm7/
2fxSIYK4ctVbn0H9Bpdk/ESV+Qc76JpYWQ5utbEO0/b9emFhihMfEJ8YJoMZmDv+X2vqN6oE/J/2
VTGsiFOpoh9QBbApfibJn60GIyyXDdpQKglSnH4nyBajQGmAL3taxFLSIsoXVG8FY/K34UyrXSWW
83WKZR9IZAIedWjB1lok2n8eoOiZWVTTAUz3CEL1YuCfM31/sPQ11i+I4269C9lkZVkCwOVVwY+r
Lynypvfeoh5bE32Il2+kqWAoaDSE5pnn0bcRdVmuZyhGtbKjxYV4mv2UvYQyLzNyagjspfzjcvgc
a8NTCX2lqj3LeHxscrMJ5lEL97rIxNsGkrM0PMpTzeuxD0UhCfD9oTLkGXlMbUm1CnzkgTGBLUrB
B6sE584g8OdzWyuYYDzIJ+4TDY8lZb+H/oMWA9JLvHdTbA8SrLYBjaqIR2/nwWMV4LAeOIoyY4t/
hWOj4CgnZoEKUBraPkFsnXFIlNdgvOfG1ATKHCyHFU2z33MBI05YNvHqNbBI/2j9+HhUg4CrEswp
zqJrFYn/NBCaG8312jT91H2wIyguqMhz1XT7i2ftMID94pUMrp45mX8CDrCT3oWzWkBUoB3mmUs6
zhhmHH4axE6NCNzNLMgJfqX0MXCsUUwp3EC849uHh3MLNwnuksXOkEUfmHnnw4jxVqNMhJr+qlrX
qmHqyc/B/BEYfTAYBxxXLA5wyzPeYf+YeU2wuCjp+VpR0SC3zmBAFfckIToDJhL/jgyhd61Ed1+U
gFgc8q4vWLO3VV+o6RwzgMrt/wyAUVvAt37roeFOYgVO7qivWg4/rF2mEmBKGs7xZd4RUNpkatss
4vdpDDZYcuUbgwWcJ5AelQ1jyjm8ureJ0656lHnhZbfTBgEu6eIEUlzI5KMAWegD7BNGkKUW0R68
w3ctq9dus1F6zHB53lo+0M8LOvGVE+z+0yjWa9liyxEI6VNeTqqzvjbbcZo/KXNnkL5EdBpkI2lV
aUySh7llEhrvj7LKsemqEeiL46n6mNx+KwllQhN0L9JCg45Q7Fh+AuPPnloyvFHG6XW8io1AxUns
h66+TWmkxDp8AEdpz0KmX/y0rsSRrrm6C9QhGTXIebk5lCxnBREj2qoO0DphkrpUbDHIgQfV/hC+
ZD5CaYKgbbC4wpFbYheDCeSt/xwZxG/57tQZnPTjN6ykGoFidzyE1G6rj4KQC/R0GLxWuTTla6nw
mRTDvV7h5mPPQvylI8Kyvj+iLiFEHzkOIwZhy3B4zOToy0WBe6hyXEycwqCaLa9gqBUGPnTHyUod
RoLP1tQqD4leeUQx0lgwDOUMBNbXUsKU2VdyDCwWEKcH1kFcpbR1Q0Sl9+ATRcOK6A6zD8orjMrh
MU4fTYfzbrB83rrl4pWS8YpwdJV/S6/oID2jKJ6E9Mi0pzCbrWc+txOAZ5NXx7/4k6XAK8qlCnE0
oGNwuTuGsOWhXTL11yYi7ztr/EYGep6cUJe8FYH6+NoZwpubGHlUAG3xVA69gd+olQj96VbbJMdc
c5AQSFfkBe44cVNM4njrGahc06xR7oh17t1mYbcJxqyAeU13tagyXfbvUiYS/lfaGoB83mHrNFTr
KJmkUgI/AiVcyl3PBYdMe4xh7oCPUUg7mpazgb+NNNlgKClLljTVzOSZq7cbWqpKNgf0beJNWu6P
R1Uadc5+C4qCiF7Zs4BZemvt1waDjysVjgsJEDkMzM6h0UmNYWM/UEKJVhJK7McCRCaB+ycf5fIT
QghcoCdlPY/HiXjSs6r6kNPgw9Wn9J1cmogfovTvOqEhvInMzBzWkEvbpyFsd4Z5/qkS7WVIsLaF
57veYVWo6sLq36xsEtIEd72A+m1Nb56601WVg4Z3awYSmjscjJeWyb3xbd7SM7vFY1rHJGJViCJ0
4SDEZNMYAcDNVFORnpoVWCkZFe1iUcttNaXDnvh7cyPz7+VALpn6LEmkSmxHKrfHY3V7YW5NkldQ
qTrK2DbeMeQ3iQnVg/zfT79/jHVKT1nU6wKh6Xel0wDIeu02J1ETXVdnRX7xIMRNlaGzjGPgyxJD
O/vuGgVbocLcC600PHXeSvATzi1nSoKHPi9kkmF4BdRukcDJQyj98tuqbxtsCFEbYGWmXaROMAmp
BmpogdKV/HGkGtkZQ+inMe30jL0XzIDmRk3kh4G/ZqFkPDJcLhUR6O8NOoRc7CcHAPuLWDHWnxlI
zePkhUDX5i1/jJiYfk+duQ96eGWQgHJb3qW1IWG6XJF2MO4rX54ITvRFAo+F4FbaxPtG0o7wZ/NR
vj4yDHfTLcX7/W0ghMQy0r7hN+2JTuDW+pcHEA+AUr6pPPG9kAvNQPm1YUICzpJhd4fudgXZ3jnf
TAL4Fn9B8L+NqCDnbfD1NKtHY6Rfq9jdywu9o1JVlQcMJfnE+XORzgaKfRThV03RLgbc7HjiMutJ
4y3rfRxn322r3pi2rfN0K28ovM0z1ZyJOHzOymUeV2Eae0nsn/9/CQ9As/kGkbb2OoVMvqdaa8UT
M1LR4omNDYwK2+ifp/4uEF8ABATy71x1m9HYF08qdbAHUHvGmbAuum+6U+F4t0XhOENN3dYDSCx/
wFrX8r3EsNA6GBrMRQASr9PePKz1Xct1eQgkG0h0zBas5QknRUCjsHpfrKtW36/m+ZYA4IYvhbMM
abrSBdbYxToMjMbmNkyungQgMJjrgtuIx0J7Kr8mdZGcMdgALEriM6qKPwTJsVc0/AYGPVKkCk4a
kNT7qErGCR3dMhAHGfZ3FShDAxMdLsZhpyluG7CB8TtVXmw3NB3+l0HY1FdY8aQ1fNSBFLA5x6S7
Ma8YLaz8k4u3sE1spN4m4hWfKBQU6T8KOcRr9S2z3ZRjeQIKg234P5zqYl1A7fDGMgyRk98PcwyH
4kjiQPCG5CIdR/tVqKOAyVWsYrmGnS/3cdBqT7/0M0PtC/RLgOVAJiUAomweQjpAfimKkdoyTMdz
NCaNjLSGthm58jajddTMSJMDVtYHAYgc8E9UUdQeb+tr8HaOCFGiphRPMQanjfukhX2vpAao2Sms
7sSG41fF1V6/TbSgpBY8WLk4SzNNqL93W86Kf1ytMAmqJYoHSTKd/oYO6wCXi5lAChVaAxtAdwO8
EyOf2k20Yl8+IZ3dbQgzB/zvJbwwzQ5uemEf8mAOpQXNb5xgVStgI4wtF0q538+3jFD153IPylwa
5G3MH07uVCwKLYHVANSF6kYi3iM7bPqhPzXTsUwwWg1fXRp9+pML3eb/UP+5wkDDIanmpKOli8yv
1q7KN7qUAOkC2xJEPvQcXAzCiUkJEdGwXhZgNTfpTYnlY7J6pBCY5VXG0CpENn6/98b48p+QZEI4
zFaSqZE33leggH6RVDNQifboRCylhvtsN97IYN15BiB7H82jfIzk5kvnL2pR0PejmY7C1zvdT/wU
+vUHfxp6l7xOCP8GEFxMyPoTBsOEDO0zhaoNlkrxHKmLOikg+L6gBntXOQHu/AGJ3qqGPELFWJ2S
fXcO3DlkZmyw9i/PrSTdnc7xwljNxdMAdsyLmzgAQpiQ0+y5GFgvMMPCFVSwOX4nz5/r1OG/yxOi
8QRXOU6NaXKhs+Uwf88omvzkLbpS77Xm4zKx2htctnoDpeScLOaB3MxyIX83JtTVAxKMiDQ8eUqN
RVGyo+iG3CrxB5ofMSx1NyQuVu+P9dWBZG+3XUcKh1NcSHKisqjGaEFYglSgjYECKsAkhVkULomi
PNi3BhsGdep1Hk2qXIBKjikBvgouK8cL+c0F+TRWKoUSy+TxZb1t+YuqwAvp7dzFs/qKujB9VnAe
cFrkie0aCn2aM5/+3kFO4LL0f7r9NxPgpGsz1F5BAXydfLZ54JzzrXKXGRaNWUzQTsh/dH5S7kpO
rBlcJTW4/5h3qivO5MWHR3WAwGSV7RTuDpnB2Ih2uV77ap4oueMsnsFPLBQno64DedUbil1Wpaje
clDxGRdqh5hW7giTFmQg33516ygpH5Dnw/tKasNHn3xghitkxAjf2aSPY8DqXK57MMFvLPGDb799
KyjcMqSnAHXahks/iaSYW5ig4KYOKD9CkrPMEn99KsBWYTKJjcccxXQC7069MOGeL7F4qEi/AAil
3/VKTgGfAgLvAEMd0WbvHAqgPCgKJh52N2V0yYPWD4fSBdm6D+Jz5M4QuZseK5qHc/f4PK+hpFFN
Y7ODT0zeS8TR5kv+lKzTpN4EuWuEy+P+vj73c0c9XxmrkYU1EVz552x4ElNhyMWyoFPt4ndFW88y
oQ1XMxscAkf/sW9uhgcxZwW+yxR0WKA6RLgLDHbZxwqHO3DcAU/yA3bPnjN9egNEcNpgZ4fGn13d
MThK11z7TnZUx9sVP/aRfLyEA75mGeqlSQtxSl0MrNOb5SxAAHDvDYT2tErza7lfCMot1Exr4jYZ
vmTrPrjBxtFH8tQjQI+D5GVspAb/U2b7FPIJfnNC2g5CaQSTQkAZ/UAE4eg1AeVxag8Kh+iYXEaY
NPML5y2Gh89XfhIb/KlpHBIIZEhaOlD/BEeIsMVrBoDsHxn917DGBtsPiGbS+7ggS4TRcYkVmslx
SLW3r3VhH7qRojYQS04z3LgCjZzHVFZuEKNK97rYKe/stvNuClb3kHhg1vid1rhgzSqJiSuq62o5
1WJTuOg0tWJVTaJzgbD6zP9QkysNQmEmmavGXFhFZgSKiDQrhPu1pzmmfPB1FPzNANUSRZpxb3Nf
5UCY6wJnTKiNlv7QMnI3NLmDJN3uQSc6Mw3HWV8tjeN5hNsL0Y03Q6bwXERtxQexzM+gXkioo/MP
HLnLoOOiztUMMlOcWm75ZgyQtV8gpNS8BLEmXurKKVTyJijTi7Lx+TRlaRBXlC880ryPzdC3yni5
c4HDSIOk9+qeiNn1moyZhhIGVENQxzjrQudLBxm65gU7RLGlA0T8nLJ7Jrzdi9XvrCWIlIGlmI78
h8vnjgGTeVJImPPuqmyWNB9uERgQmglGNPtEdyoIJEoBvCSC9ja+VrATyXbqvjCgGBQYcy3kw0h5
CLuTLfJaoz4e+qzzixK2dr+xDWsn5vxgLMeOi5VThHEkQv+0rual+MOIWFqM39hykanS2X+70UBh
Pic8ubMlW+c5ce8k5p3NLfJsbJg1+A/WReymUteaXeSM/QxTmHrlBEWMLniX6bhfJ2t3uH1iwum4
89ZJUnmGvqKNJX8QEUe+RiGEtS/C15WoeGLsbJwNaGU8s6AGnpunpFUlUCZlAY42H2uqVxB8d+si
WpwL4QkE/De3FUT0BuIp/soEbpcgGAQG2iQLtrbLreNzkZCtBrx5TwilkSmwahm7WfcgYiCVhERb
zBX/N5YRDDx44OcmNmmfx3HAZENR8BNRN+lzwZ6Pp1z/GHoPwaR31iRyBpWgDMH1oHcaLXOWPRxc
fmU7h5yne7fgZvDueHM6GyDZTJErJWh0+566o8Sb5Mdbj2p7+Y1BZpVPgYvZtCztNr/TA3JzQhVP
jM9HUklEAOBt5b1i2U8K3217TQ799KYc1NaYhQO+oCUI6zybQisFrKtZKPy1AlJ8PdlTPk96BIpp
oHKuUxIEWzdLeBeME/QMG2J+BG7+YvWN083QMXQld/dEzZMU/KHfvqHSsVg3EeEDgprv1nf43o52
JabOWnOaEMcr5aAJq2sUOlUMRAS3Rwp9OClFEemjP0V4e1hYECM2U5nRs0NGsITutm3u7xCKNvJ7
bvXw6R2qZ0tKeL42Fk0pzhhg1h9xRUDErOTdpcjcJXQ4oniLwIRux1ph9cwYOqow4kgb1JYH8s79
29jJNM0CS36ylrHj5VtvzesBqdRj6y7ujHL+JScWn3XkdQpST5CDV/Wc9XMgwGpTcveC/Xa8Exbq
Fk+wINrDT3suQYJrpnkFTJUCyu2hV3siy2DsNV+uFuKPrUYJtxEU4+vnpRX/Od9yQNKkYlqHPb92
mInjXsH+10EZupxhQHDUQrkuYiSRU29BS243L9uV0wmGY2uoOKg650Ce703tPn9gNP1rFTVhPwka
Aos7e8fcEh/Af2pbS46kxfaq22q7wibDZmgmSUa+f4p6g7dwx0DwOvnpxVvufSo4RPb3+U8Inv53
8jLlP7hIMI9FGNxw9USpB94GWC/E9lzAB2UseBo5DoFImy2+5l6hBKfpfcOWQbFFQWaPNiG9JfTz
hXDmFDbAnQy9ID1DkdfBeOENyWQfwlRxPsR7XVDCSfOtejwJubpU6077nywmoE+gQav+Jmyfw19T
OW3Jci3vEYvkWAVax67xGy2NB7U2FXFMHQsOhvdC5KtGY6G9brkWY/2XKE/lt5MuT421gzma4tEC
GjE6ezt0T3vsr8BVMwAFWBGixKTYn/vLjuUVARwB5Fk0fW6imLM4hN+yluP7J/2RRnRuQzNkonou
QKpAXr8LKA5xS+b6zOrnDKwg9GQvSn4lU2pZclxcUYyghGhdyGp/lfjYipHtrcvYiXX0ZZF706az
i5iKbEi5ZjWkmhX2BtWOg9jkqjkLqyDyKeQfG1ubd9UzlIjoZ3grJ5p0Mu40oZ94BkcuSWEtutKD
mwg9dAPj/yUjNxC+E+4ibZhPX1ku52GglzynfQMMS7hRBxpoh/Do+H4OeYzKmoe7WjFwJCdmWLCZ
Bm+Gdr0sfCeTsqL42U91H0kqmToZxhWO/64yXpv6yHlVWlL37axRSCJ/7Rv4KmQgHHCz4lRwYU6O
2QL4JsOirU2L4vTxFR6MjHC8n0Bu00ShhFDJtZnPFmXNPrXzYQPd6ejVf+PeVU50Whxg8Hm5pNVP
vh/AlmfEdSuFJkTOURoEA7ewGlsIfRZK3ojvSR/G/beIsH1LBrdHaoRuOheC1dQb2DrlJKX3l8PW
IkDok9PZHEUQIBSp5gEwcc5SG/zNTEmP1JjoESp/76q0A/7cLq9awn5osnBR/STngv17+NwAQdH2
li4W4GAILzMCBmHhhub3rmxUWKfXj3YVrZr354Ktc1zxAASeWq1+pNJ1DWwTMDAle8qWWb92qOvF
f3LMuFHCabXio4U5jBGCPCBFgvsmidctexu2WKwxK02BpRBtOs91ppghO5B5MSib1WwwH0l7IXbP
wZi01Mtxo7jRT3GnjEDuVB6HiMIZqD2DSpCrSVrHA+QLXMcU5w3FdWlsyTwZrZd5RkoKpwkDEMfU
DlEyV0xBXzgk3+li+lK9X/oIQNRKNO1/7pzoSHKQb7HwsTkFDoVPQZDvUGtawy4XkJm3wv0bWlbe
d/tE450wzM/TYu/BVSbfpKwC2pByn623SbZZlKIFswOBeb+McmAF8HirrH4q1KsrIk+7J7yFbtEI
7OeSz4M99LQjEqNiK0ieWgDuRKWMCMrQfh4OAyQmD2xmxUndzrPuUk7vLRGJtbZ9LxTCgeXgdZWk
m1e2J13GXiOw811PLAahkhlFOR+5NYUyoJVoPxpbJmsREfVZpYWKEtyN13P4WXA88/do+QdeO5vz
7N5734vLrq2CJmkO5gmXlYDqO6pFElFslDdzxbbJdfxXPN/+ybqBGMxx/U2SgZMHM+mrhY/dCxrC
wXj8XEb4FYYo7kVXuwfLotH5ZOskcVxzCYc1VFTr9QyNJyQkFUsZTQlwaK8jCtnlKITdlnEBs548
QdBrmP490LN5t25iT4qhERGFEILOUbJGWWtZ/LEAWlK6pYUugBsL84NDczxK8lq4Tj1aYQ8+Q0WW
yEOoJLohxW3bEU+rP7+RdHihnyngu7A9kwJVazEjCa3U0D1L+1at3F5YSgru20/GvhfKA2BW1crS
vW8bbwSF7q6uX+MBNGEXZQBkjJMXLkQ561Xyt3FD1yEcNgZwZHBHm+zpd+F7j7G/hX9xqMlcFLe1
2h3UEkH7Q7VMJnSP/5xAm+Zf/h4O0G3LFyR5i2WHzhE8kGxbaoYzR3k/w8WvaZ0h2AXaia5SdU9k
TjGTF0MuB1C5ZmMfd1RJtmIKJM4/NjUCOd3TD5m1V2YBHXTZ8hpjN+DlKQkJDWIjgeCPLPHvtUh/
OX/JjBV8GzweZ5gW8/NwN79TXRCqpYTCE+/lyjCFfAsLxoxVyCJUjPSm5R7MCXngA+AzzFyzRrUk
CTekjAWvqXvMyNxn1YE8d+nmqham4//6gxQKTP1quBXZp+ZUYWlzpz0r89o5vrMsOk/3RsTYhaAl
POefu3v5MEKvxlkiPwWUny73Q+PK7P+DzjaVSsdGNZzOfzumX6nMGoktC+M/pyTyQ8WuKtnqwl7y
VunNRj5QRDAE109i98tzuIqZgjyljjJxYeMSJEzvnOg965IDJoCKjpeQqjbambeNzcCsVyPaahsr
t6i0haoBaQ3KsqB6K1aHFK9maSpnAY5zDcIx4vyCRGawCQ7l+SLYFVqNdnyvYkUJJbcfzNf9fnUi
Lj30AX4zxBuivRat5dgcBTXJy6hjRZyGMP/VfyiUD6hGd1V6BDEmdfQ5uciDu/FbMBqycFeHXOuU
Om5rpVi4QR/6TQOrIg+TsZkMB9LRuz+FW74hFGKvHzicquWvqPzG5T2eXJmJLxOfzPWAmVdskisq
7OxUfe/A2HULlJCbFtrqI/h68izYpHOQV6Iur6v4CMbW+P1e/6z553peMl1N0LixCg/xgdMWBc64
THuF777m2ybsxC0oWQciMDZk3a2fX5+zLJBArFtFZssJqNNfIquJLvZ4ScifQD9A4ohL/lfi7Usc
fXCHjtXwspkz0Gf1lVg49NML/FqsGsgiIr3Tv1RwviKNML8ZAYyhIAlYWQAOFMKna2oYHfVHXQzV
Ovn8IS5t/MvQY6K1KxNKoSl5IJQDMKfXdQ2agxLU9klBO+ibi4LfJYArg/UAd1tlF64y9QIfkrXx
cbARW3hqVez08EEC4U18qKb3gJSbnUTs6uBpdRfmsThMLlDD55VcsBPdcWIn8nFi8/28aGra47NN
kyLEMbopgIfJCIfakSdYXRrxqGDjWak/TzB/ZwtQKcJwxrefIC4BgJqaWLX/5YpJVw0NCMUQgykd
hWS4wugoQkA/5TcURt/NrselYnJhebPiyBRn2zzSfmmiHBaKarKyR/i2JyQaGj+J2pZIWX+wgqiw
CTJ7gDg5eb/LKV133zO3nTB1NznUtTopGNCrWgehVFYWmXSHrJf800o8BUMcWfKzm/eOswC9aT5i
XWQyMwx8INLhasSpucEbFpoTQ6vxVVqvq+WlplSdrM77tx3qKuD55xjoeJ3CnSRENjlcgVoHrYbY
QA4NFh1mF8j3FINxpOOnFrcHYL1gkzMPriTFoE92339qzH7GqkzEXObfPqKtsTQkViWAHmxEL0mo
oIpNETHtB87Z8pb9wIdCAW6kzJUblxhK09YqSuhYnMmEJYfVMQGO/gyLtpCLubrOPuPJ81zGhzcY
WLhWpxWU7uAAL5YOlgmYJvCbTJnTM2ZQd0v7ZngBVbRB8K5OMwid0VeJNvApCCVDfVc4a/m40AXp
2MXnt0smz1ZZbwocJ322MSe7fxtWalTA95DyZT/uwDCpd4YtXpie2fC2yI0kISw9qLg7BN5CbW/m
MgIS8gLWcJ8Xy0sJ8wwJJn60xmaL9tOdKjHWsCiyuW28j/4vXqOD4vAUPXq+PYT505PIoaiP5xUM
lm3BOsaCj+GNgk+HAnprhp+LODIaXP2QWVY/xB41bo/36SYd6A6B4IwGnMFpDOxasvCIQ+PsgQO+
y/lJtJGyRhbsaHN8u69ktSgjejLDAzWXwFlsRjroW00U3KNB8Xnfi5TgPPqc5CpT1VXSF0yWrWP3
phVgRfCm8ytjbXs3AtyviP5L5AglhvHy8tjv9jJd3p1fd5VVV/5qHDqezngQTzGM0jg5PzH1mZN/
OHmYRdS9Y8lHJC8VFLhZsAr4BWRI7YbbKouAtKmE0Gt5iLITENk2Xj0CNq2un7Rob0aYQqh8nCyb
hmMrFnj7vbUJptvkdqluvTU0oWf+8eJOrn+NtKNJcl++uDwcR72eOFM6SuGBKd+954RMRNBypRX/
SE8/UtE2+UOn5TJPbYm+dTnQX7Y2ISkA+KzP+2aPTR4ToUm6uFVntHTF3Qe7LwkVdGigPK6gxEyl
+5BhBoxolWAgortsxK6puXeycsI+YZ5+6GBTaWKfm+8qdQ+udl4KpTr1uN/SNfTDc2X/b+hGof8t
jyOM7aAk62Lqe3sQNdaOwnbpV9l0dNu8FTqjJmwSrGNMGjyyz9evZz6uql4+zc8khZRvHovsOjmK
aICJGZ7xaOYtGJsQtzHv+Y5GrUDtkv16hxi8PvO1ATqcWfQ9QQuRqnF4PWsuTYAMicLv6vQ2z7U9
DkfscyJOOiNwWhkWuLoS85mOrGfSFPRyF7V4UyB2/jwrAmGkVbi8cdjd7Giwuvj2QzMrdN9Dr1iK
HwdYdaOMUXZXy4tntBGcyHoCul+AHOdMXdEDYcK19KHQ6D0QJLyoPkTKM/Smck7zQTnsLnFCLRBR
mc0m2mfH0tPthszSL0kvDjyCST2uMqZiBAWHzcmFcUhxyM0hb7fmuIr3nuH4N97lUT7NCwihjWmZ
RvKdkQYgId3x+LkEj9/9fCVw0cBi4nk7VS5YUd/XddMpRPUft/cKmnlfbKMP3CQIKsDx1octIJSF
pRmOEuT9ONZEnMUKqOSvmKwtjcx6q9/hv/YLQWo84Oh2AHg9YinUj4nYOz5/Nl8BrZUahbK01WuR
anF44uw/V+HzRnZz88dgj+HOoaMs84NiSOX51DN0tLsaX7IFlPJoLFN3AAv5ymXlrkr8p/SM/VWf
rshVjDdyj0S3TOQgaAevL4huZaP312ugvSdqsgT24+k2XN12VJgo5HKP/5yTmXMr30R8UzC0k5pr
JIgvDSb48oTGXLRMuspvuPaNwga6pnRE7f8zZLWU1cr0U0gLv0HFl7oBum3S+jl6O9FAg7Fgtsf4
t2vyI2s6U92dO2ozjPervuPapsgL2MRAkRbb34SE/1/rDiaMsiv1YZWkwpni4wKV3Vrjb+/4tnzF
whVexgoRd++DVtZnXI315pzgYIphL7fKuHiwtJa9HbW7Yy485Q/bVptXt1Se/rqkLsSA6CdiX5Kl
tqw6RDGPDSq3boXoGXcfjw2ecEXsuA34PI+TMK0KlpQ3MFIH1KvGr3CZz/2molFTrQiHdFL1iS5U
0pWxrIDt1mt/IdV3Ld2EvQIzzj7ZFFu1Pl6dDmy70FBaCmdzB+yuuQ4nhfGBqOJLJt6XAWkO4eLK
qaH+pth83jFLQeHaL3kDAniXVmnolorJ9gMci7Bq7LFTISlBKT81VsDbjifEYfA1fdpVR29EKgju
0RyThpaFbGc9oSg9d+BnguMDF6UQlcRPww0977xs/w4TkeJbgM8UYS24TLJJBt5GY8CTFj9GrASP
jYJZW0iUnFxXE3RUA9/q2C6nfS1/d4Pq3DlMeBkeBrbDiPTnakdnVTIoz6t9OVgNi7blY0f/DFVy
ZBiWCuRcTYruEaynttzglD5oCDVwHDf9mp/YglTSorM1vcUNHtxFygkUM31Ia+6bcNtfdSYPYSLU
AhZzVIHPFTMtDKKMepiHct9GUJUxvCzuyAW+TsYIoyNQ0YOUV1Qw9vNQrOiOI+tTc5HQENkml9jn
Dnp6vHRqtRYzI11al4EUcd/MdlQ/Y1bYCo8449mtEeHdKanh0Tae6sMJP4H1ub3NCO3rSeELHYWo
BZbUR5oXDvlYYZ3laRZtB5B0Xm3GiA48ZF2PI9rmy0stUJ8Cv39avenx4n0HV78EMnLM9OySI87Q
xbf3aAHsDX8m1anAqD20R/w2UP1Rgdkz628fu1fTPlbhtjoVT69RMmrgcyHrfrwh6Y+CSe470a/X
EAY36fDFqcmCdUZDIcclkkPp2EPQT4BAr69jVjyQodtS40BCQ5AAvgIQSwfu/D1R1TcW/+nvRBzl
wk7383D1QKqhprK/nxIKfH/Usf2vd+dHnBd8k/WGK1TgizYvSj4npAUGkz9LRB8T/daEjk8prJnA
EkQKqAaNuXMS2ksbC8x4rQiJZFSj0rujV1R2YvJuhjEs1qFmr53y1cheF81bYcyyfQYpTD9ssigv
7gqYOxPeTDlOyKQ+k43epi6kZPYsG1DUkqBexSLnCH1KxRGe97qyEUEFL90WCVx5nKiu1jJqmkSc
xVDFEoqAJ+WHf/lprl7j5R//Cbt7GrzZnKzhZmV3Y42P4b012GQklRzhGCAvDy5XjngstHduf4GJ
7UpWzLeJ256FpkkW2C7m9YtCGJ11UiFjAkjl9nBVkxmJJI6fOTPOeeE0XiYEc/Iwhnspgqn+z4Jg
kKMpNRU4x7/DqnhsAWWKK05TDy+Hpp+Pn+LbHxKIP12ROGVcYkz4dEqWd7UAcW/sWswzmI0gbrnh
y/f4Loq0mgqDHUFCGO6PEM1WyDfWTpAzjcDH5cp47YazYzYxlxFi+kai9TmXkGgp0yddw8JMhkTl
h42h0L5QzM0PJDc9gpwhwIDNx+egs/RoTvwFuadsVEm4kvLzBEmX9pUfVWhwQpioItwXufQrJ3w9
PFanJ+cu6ume99r6uVBH0Sywd87WFyKUkOFRmQ6U1ZCItwGpwKKneC9Plhm5Tpmuj7W5qoTHLOpv
uV9AIJi7EtsOpDLG18msH12foEwUT0PHCSgy7dFE0yA1hXhC23eQph6INVFlxGKuaCZ93zyFs0Fa
iLTQz5wySDHRonuB+TTvsfOY1QJplgrJroeeleZreVa4JxHYXkYraWVxJtSWHyjJ4XWaa73OUihI
yhHgfSJIROvMkv/z99s+r1aD4p0LpL2583t4qchYc1uqKshMYrRGPhug9CRt9N8G2iY89Q6Vl0oW
vE4uPgUxnxtgjH1ArHfU3l6iGfGXt1yIOsZflVlHp5kJz3RJJpzAQ519UWlqBVL9+dkqoACg8FeP
JNU9GSDw7HLDppzrfNosudbSoKiCVyc0mHk51IIxAELssmCN/MJYxMYiXF9clswDyNXuXfzS1emn
7m2hYEP84xVHd57gif/ySQRdmiByeKZGu2PeapqM3l8nxRh/WWTB96WfuuZmWRkHr2PtfNH5PvRW
hOoIMyRRooxW3w1FBW2/z7FzL4uMPsG7SWhKpeuScZIkjGhSX8oSjRF925hscSHZTQmTaFXpcW6J
cZusP6HcQFYgw+EhC334SLNoIMGvj8Y2Q1YC2c/CL3kT5lJ4SO9LJqXrTLGAsDDGcgc0bk4H2du/
i3WWXaXRf5ps9/T3LeKfjZvonxCPHdSR7qINLIKNeF874bo6VDuGE9uYHSwOQ7WaX7oRWQApAHNS
J5TeVxD7XKvWaiiQVl4TV9+J+TUXqxhoF2RgIXLAU29iSoLdnOVuRgwiuoDK4cHb+9thS9+3mkjS
AmMWA99AK3/wOtI+oxe818cgDlnWHerUlcQpZV7ahP4gLEUruv0gDmtvtgifG3APnKHSRivNdQpi
R9nxNHveimrnaZCwQa8VMsCyWN+hhRHJ4BKRn0F3/4hF5CD+k0Ofb6cguqRxidJtwmxxUkHLvKME
VZil12r3OZ0lv/Hb54ayfgMCui+5pLWtzo+z0UI4m5Oj7ufyZoOGDAJoHWUELBu0mrwD6zgbWLJo
0SCrbBvef9s4SAu7awlKbm5YdFuZTShTY3Yd+OJ8psa4dURK34NkBuQVV1dhS5cx20ThqMRGL7mp
Zj0EXLsxNvw1j2b/lFiVk26Hsim493Ik6MCSnhmwR+MroTjc3z6k7ci8pxdHZmLQzwbD9bqkgMHW
DWVShG/m1QeF5pibgwr/eqmjFv7LN2cwutjPf7WJAcZcrbNr/U4E+Wa4y68/2bdEPntycW2hHvu5
cTwaHEDqvEvDIgvQ1MlDaUvty14yRUFgb+NX65cD+bFtmsXPMAJDqwMaY5dfWRLBmKuSccCvYyfb
809squnjtMjnbEHtTq68Pt9wEnl1biBGtprjm5xxidxbEiwEo81NFk35r4EnHEXxnvdta+h1UkiP
vOBUouSdZ7Q8gk3TDCbt7wD1aYBpf4T96+zMDGwtcrd2TmZw2S3aCkMmBHwEcpfTEeYNxhj/7GBR
A0jGSumzcJez+Neu+CD9B4HYWklJVjoo7MFe2qc/DdfCThEKCb6OFGokHfzHzDpyYUX7tzE0roLI
RLnnnHeb7QvgcHgKWPwwNfTKbnJwpFtiv2IKWYULGn5NQ9XCfYP8DFj6jlTAdRp5L+MIs0fM4jRI
mZcDqgLZucU4ETIGFkCQagWPQdUd2l8bhwcfBrn8QwjY3N2mrrR1a8xr4t7kcbarU5ptaLWTdX9F
9pMJuF5QDRamCPd/2d4Ik+WG0hY1Z4Apb996ebWz38V1mKRPRDqjqdTmCU8edsON+ICX5ou7mZqT
OPXmAWDsPrVRE97Lcuq26pGSbjRG5nNaUBpO4+waaE/cYwuZHF/yCvWy4gh2E6URoE8cD+9bzOV+
NLorwwX6zER3NktAzUetXFaH5/wAwb1WQCM9xnumJtkfSVU3JhCQVmLB3zu0E7H9V4hMmdtJ2b1p
vKvARpt7NRdRjQ5mIjbJxc1NH9QNw32gYQkYVaCePQ/xJhsjOEpae5zJslK7+rpqNBY9km3nypK5
xx5WWZtQlS0XIHXSvBR89n7v/pc8oQVUBmN2/KCLNAvyF0WudZidNKgLPiYLToe0Ft4JFpH7rt4r
2HWST5Rs14wjq2afOhFHMXSljDa3CYbz9yvxM0RsitU2l2C9g5Y2bGMfQSsatkUnCVmvPWNERB7F
Nv4Nabe0zusM7ZfcaMRdBQQgbz1aA7gDsWPVfpRZ0lDxPE7JPeMXC22XvzdKb85l5zKRp1S5urjo
T5l5u7WllGCH3C2P58wNzpYk74urmIT7NABSTRsv1vtaX5aJkKAvQ+sm5gpHArhQUKjhJjLXdKEA
61+m+1Ki2BhJqQf4RmQHH0fRC3pM5dqgQiQVEFqVFTV1yqNIuDxjuYQXKBYrEAxU3odoPI4Ym3Eq
UgVHGwOvAFkahbT3yAtpgtpoEgcrwNZVs9hCMDb8YqCaNvFscGJrQTlRlYpBTXT1CNl8ki8bV5Bz
4aJ02xVA9CvB8ogEv6WB2DMKE/4KV3hgt52xux0dxihXnIS04WYn6W8a4A9vbMhJwHtINCGMPdwJ
9rMSgeRW30SyV7fJyqkUJxZbUmXSz+mxal6aRY7J31SSISkyBpi4ynX/Z3NjvxVFxMm1B8oqKwGR
1Rb2O+vdrFjmLiTMNqnPZNYP79g1JCcgzD3GgrlbOQduH/WGcgk4xxAIp7rvS8xL6Wg5wcfBEfFa
IILWvsHLqu2r4iuFpx7RmobW1Vxh+G3WMYbN4tw+z1/XyvMCzLITwWYUownm2nywZCh5xqHzJ6xt
K9gDoROI//DBTZ5vqZTRR9nsIg4maFrNOmtwsmwIORvVu5yocedG84GCQbyUF3gNpG4C7PJJ4rlQ
xhXnzke8kUjQFPQX+i3lLXk36ZLedfqLRweYtABstwFprVYYyLLzPeEwVoDSwHF0gxDHJUty0bZm
Ck8QzWzs1cqBm8ojJDtDV2bxvmhYRDxDYeLxGVrb0mCo07V+xARgoE9Ve3XWNukfpiK6KUGxMbkN
c6ZX/pmwK9qRcxZfJknH5uhWi1TBB9lt/9FyfgBHoZgWLItQEC6AItI7zYp2I9BwvQNwIRgt8NPE
ubxygJSvpWP8myIQGVrY1oxKy8hqnblrTidONnsoGN8jIFgz9Bpa4Z6lw3eawqZ0Xdb38pGighFR
wujLWCBXFJNa0ukng0YYhD0den1Xn3ifYj4JE9stor1iNI1xsjvUTVhNxfNtDvH6kT/xoLtER5Zl
wP/tlpsP40SVDacL0FFKzoVNbWi+gDs+PO/p1Tue92yizznz3US9Miu60KGfsumq+z+65AGwWsoP
f6gZdTEvL6m4QseameG8txgmOXFaEPw3xEPfzXUX68fl1qOXQ+U07IsL5dXfrmhxosgyBtzYDTda
Z7Z4A2ZfoAfF0/xMeUS1DuE9K2KsBWLHP/mzReDtWRa6lDajKF+gN1CfADZYc8Xiv7Vy9cEeA9Iy
ggSV7VjpAZkc3JmmLOnKawMr2xKZX918sEzCRjUrWWtctm+/QjbVyuZuELQZnjbi4fT+OCceV5OI
UfxGnabpCAmlU3YAWzj89+v9tfsnpG6mAALfmhUqyer+YwPDsO52quo4GLc3kLuHOGbksIH/H9cT
05CMLrrMuCX9KBulxK4OKmDN7gfJDEgt5Zbisx55iN2thiLRo7P7a9OWSmRPSxo/Q8oUM+jEXIdz
QIqqkEYOnEMf7bPDx5pT/H20SW+X8lMl9Je7PuMF7I4Ht7ggnK0SCj3gKkFVWgBlBDX/S698adwc
ZQosuWzCdjQzVLGBrvDzbeavOPBylL3adcyoDCXoqGC8IwNRM252/mga1dmm+sfez/57nb/TMRCK
UTpwbfucI+/WVLTwyl0JCFH0mI5t8hvf6uVNrIcCaAZuj8+JajOoeRWb3h/z9OKkAxzJFmr+c1OX
lZWTNTVGsBcweTJZCslwiPhgTBLGVSNKfnm59+BvlFcGsFUWtN1wRQkAilzJ4jBV0scgf8zsrEV6
sJRHy1cnPsaGySAnFbU0S3t+sQKm39DP/AK9J0TMqt71kdmIywx0TyfNuYex46NbyWpZcZYVnCVe
m0mxjPzC3389fFpt63yy8JxhPhyQmaBwlIZf+r8jKT6qtCPpk8m+DA7eJ4ZXnoU8IkUloeXHI323
BR2/mYQagOCoF0E7dcWetIgkgV+ZKWMKm0taAQq/2klUDCZB3miUQdE5lN8anlN0Gi9/A9nvcYm9
wgzIOIcegBDOvLhtYY4wnJAvzAfhKxyQTEt3W6gx/l6n3yDVpHV8WIo0Upbmu/ytn9iP/Q1i34EN
WFkKo2l9LiJ8Mi59aQoTl1GgWhDWFZGITMsungn7rwgCMbQSR6MEsoHVZOzQAe4/HckjjJerPBRB
nCHO3ALZXxzST/9tpXBAYKM/gERhqklvteBfTonhGwDiQrJecpkRM75o6+dk4W+JboanaqS7c33a
KFGfoH5EyjhgTbqcCC1x7zYKMXldaBeUrU00QPOQy8o2OfvP78fmo0Fm73O2YgnaKwdYp4mh7ay/
b/xL1qFYZL9XFnOZjmnx8ZfM6dYyzmOZNJg6MGI//OIW8/dVP8WoghlHlV1XWGBKL+cNGJH2y71g
VxNLLtffhKbBa5rO9gVZgeAtjNc00+KaGqPsL87RowUKL2yVKGeRcWj2dU8BKvUMRopu5fJvlJ6S
jz2pDLNqzLymtvq/Wmc+B9bXJweKRREeU0g6+2jrS+ZQGWYBZsdHxHad4akwZ8vAubZT7uO2RRc6
y2gLduWC+w22s26pDwhcSW/nB0DXn+WSJh3sUwCF+voHy+LiU6z8QHzi0ewwGesNcZXvs1OwxAjb
C4Y3c5FOF3EeO6f25xH9Byh/IkAuEO04p3AA8F79aTcfmrH+oDVXPxhQRi+7sMl0J7tgGD+OzRw0
IPvDQogWe8HYsKRfl0qfzUhPKMbzYy8Wl+0Inbt18LTgceEv7ONPi2K5FmVnIyedrKT2JmR7ktkG
LX+0nrkBXooqovtohfrGJ5K/X3AmfbnSr0drf6RTspkeZX6YsemBsIFfz9bi+F/8vrhaxcm99qSA
WNNHoXH2YSLwBQSMhWF1LpAEPe/r5W3mPh+yt4ODAp0DiyCABgZsUwUqAHMzEz39qsB4w3C215hE
nEEm9Xo5/u8lCj5Lw+UwGRRJk5n5MIcvPUe6HaovJbzOzdhqLp0Z3Jth5R6Fh/I78mZ7fBeYUNya
fJW6tM/EE9tlqz5bzOByzkMwq4wnwIn0b95OAxIXeHEgXK4B6JdZKzzpnaGhSl6dVyPLrvnFOzta
+5bdyYta8BGSG4fMdTsAPzEoxwx/p32wPM5nq0AjusIi5cIaqN4FDkVR0hiJUuePaPajlDxZmlPK
d1c+WpKHFkRXq0Nl9VDRczNuwIwdU2PUOslCKxv424rhGqeRi5Ugloh9fNXfwR1V1h3/CLH9q/Pc
H4eNOsJ4Fk9x6i7mWIQds+HwdqCSwJFxB2kpEvwY2E3sFmXEhBiKtwyloAu2n0Z69aUEsNsSuvCS
W2GFlc39IrTlEhl1eM1C+lAKIFKeFPoMaxsQ053uEJ0GE3e28ET6ENkkp+2zAqzU0rfnAexnWnlQ
2xdzrMcF5GyuOsJwsmkuXsePIVySf0++k2O7tlr8zW48yX5BmEMaBo0SoUZgynNndqPNWBF2s/hG
IkKMT8Jm6xBvMnJh55h8PlkLfhHqJE6dYDsvmipbAlI0ZxKSYqSv4Rg1GL5pyz0OpsH8wmwl9ifX
obiR5KGR/n564tWxYmQxm6kslhFQyzr5Q+OF+uLZOlm0xJEs2cGoNPKjiOa4HL7IMLeT5oq3ULPO
NrrlDBZA6cc2nOGepOXQWMhLhh5VJw2J3VM357FgU6daTibyKCDIRy1FID/fX96WSuyyR/0EFZ+6
KoUIUJXb+cQtfkmWqds9JNvC8pUK0LNtW7UpVDEvBnv3YbL+oNwAcWWt1sL/iYp4jBu3dd9r+k73
kOU3hywk9Pf1dBVS4uU79N6/U3HwubkUvuRHHKVKGU3HNm4umTtASGB2lMjTYBwJTZTFWoMiAeSS
NFID+eff7Lr4rOEcneJxN4wLIHPyRMT18HWAtm5EhqvfPq+pQ+JKe77POaeG/7nSDkLGXQLXyBCg
WtXSVEfzBnoWuYN1VDs8xf03j7ALarrZFusm3xl6gK5T+UMssoapIIzU49v/pTs1yWhSWmbAinQL
QgakbpI7OdiIYSSQxFOuV9XkK3Dh1xMKUvnv4M0cSW/+yutrhWmwL1nVuZPZuVpyC+OT7xTOjl7a
FQjG0GlilYcDvj3QbXXU4rOm8kBqR5UyehIFhFodGV6tdq83D59hyuoRDzKzNNqHdC3gdVT29K8x
f2OIrEdzX/geZvqoldp9U3GW/5UNDa54iBknOvodTSTPU1CQ29i+aUAUWpmkmfCG/DcGrTW4jGws
wg+tdkhrtE7qhk+5T7sSzZ+85TCPI6z/UGQLRhEanazBPmvnUMCSjRVvS+fQ7MaJBdr8oV7MdXXp
wRTFVgRwO11Q8V/l9yejRmqGuMzrKLyduGKFIK1wbTTsHZBHiVEPJahkwGDzo8KeNH1L+g0VE5Tg
5mTaIJz4HC1vmfroyFdFpvXlunBddI7vIlsEvUmBgyVgDSgTJdn0Ok6iAnaAPaYsTpFkg33PWUeI
d2HxnZYuSaqrpFkInsFoJjuyU6fCs3jt6gFcnkhEsuRox1MLKxXjv/wfXfzQ/qb47Gl4lo69GOz+
ctu3pwxIfwNe+s/EIoJJPnczyhVizThnBB+Q5+YEM7wFBLE1ctIDgDoBtYCdoEhccPKmQKIzRxZc
hsklyG7Z5gYwYU9wyNl9wf0yb1Q9Iplr6XENoueGUM7cAf9z4pnAo+CPquN4d+FMLb+iAzM3af52
IKzfGcrXHj7n5xD44DddBqfoW+/7ZoAQOeR+Sth07wPKZJFYYMEqXXjk/ygb9xTnYPqR+cIzd9KC
ncQMYvDsfZzKoQHIbtsgwI9sngudMEhcHpMeGj4DFAFxh2A8aF5Xs8sRUcqzoA+pvgst4FDisamD
4QqSgNOHIBwS/jHHQobtTxhIIsvZVBp+f5RbUV2CJuNzRdrBdpIpYT3jtG8Rmfl8hxM7AQ+besSq
Nb8wHWoDLL+/TWPFt+xBTUPcUP0XhdWifN3cB8HLqc8998mHW5B2D5ZsATjvHEFQ8KBdnzv5k5Bg
RL2SkfRTITCnYZctiltrWxurQpIBghfSQTJDyW2r2ngSrEk+o/aIRq1VCngXaQA43vUcU6+mrs7w
70Idn+xHg2Jn0gLHM80ZCljq8cRxhxaNuO7XfKrR5QTKE0epgXNKvJndV+kwBGrOqw2RdFOn9yKB
/X6KJdS1hjvofhtkDtScAgtsUKYR8fJVH1VfPF/AOy1YnbcyqfatSFYp6qJHiZw0rihT1E5kJb4B
lo60d0q1/E19aHxAvvbFtfvNZdwq56K9TeW1Ap/QZQN3w2WOh6AqU16+5o6GOl6hIhqp3orztjYW
i/ubWpx2ESIP7YSt9lEyu3PYqmaI9hnEVTwAtP+12JyGY0ii5+dL1CP74BeFBgmaNFLGf3Okqo5B
CferPUqK09rSRie3OIm580vejoKDcoURju6UGIpen9gQMEd4T3tiMENgjGWUuwDYrbcao8A5mtSr
lw26ArlV1EGE4bZKdU+8yzQ/D0ndOJJA+4n3bU9oOLov6/aXWCUNC+25xjMI95hmngct/E0D0AhL
bHQzPyF62zTNiNe82jNzeVY3CKrqXkNETsodrTVS6OU5EFYvmN5EK5wXYYjCxL5tGmhSLHNVxsBl
8AQYhtiuXPCKO8Bb9reGzG9Y/Q/Y3JHnNrMo/yr0a7p82JMyYmBMw/zO96WiSuGmItpzZy5rsJqf
nz5Ej93fhSD66lC5Lp8dCrK8kq8rTX/umMa4yYplSsYSUQy7b2LQcs8fS/Pv863X8mNEWOffPzkt
KMNiK41OopgfBHBcMvcmEXeXxeBi3dLWCWBiCBUa/6xz78TZLpBBadx29RqJeJ3hNDjlbV2PMMvz
y5t0sIjOWNPNpEvm0jk5d6pkSkl6QlmDIBfmC3R2c3vqkUVAE5F1TBj8ut6bmQnrr9PulJJS2Ie3
Tvpl/lRon75DWFnXXkNeKqizCBuvMTnltwzF6xq0nCqntLIKgP501GP7fd7BWqHdQokkB0Nm2OES
FTfu9LXrc/5gd9cq0DkkxtVB4oY5hwV0cQ1PmPdMUq/x0qdt+j/l7S2Vd2tp9i/EVyygemhkvsoS
//GhH6joZICE5lrig3qzyB0kHHPTRy0yWAaBPaDvPRBS+/KtXRFJc46dGDIoP4LNTIxApB9tYi6K
a5WwVUrvw5WeGw3Q2xgCCAbBuxbFxtbUJZJZ0djN0fJ8a5kwnXKC8gCVfDOVGZUQHdXBWUPcgPfG
u3vdHvIcVD2F/z9kCZ2BrXFrHsOEbMWK20zwd+zuFUZQgSRLT24VEv1M579+nMGq/dB4I9EdRLaH
naUQs+lUhc8W2iQ23PYpF1abI+f0BtbRrIPZbvZ5I8FPKB/8Vtdwia3RNCQS0gDtrx7JZSRZ969k
GvwabrIJo99PjPdsuVrsjDsnUKAFmDBJ+AnSN+jsT6CiJmIlpdzNXipoDqIeCMCYWBBAZZdL3kYV
GbFUZCLTY0fDd0+jB/dTY+CJm67ERzeSWoAQCJV9b/4ur0tOIfyYJpwhtw4PPCfQYXWXgRexT4SG
eeVeNvf8WQX6AR5Z+Vm9bhaEFheLn9mNdmg1WtCtH7RfJcu9WUSm76tvo58FQMRJIxeq/h2qjMjc
L3N1gO5UdCQ1I6JQGQSx+vTQP455nIQF81yshDLHfmTDCNGQ/YIgqzGAJsVP1MM7a5XAbkSK+ytW
Iusl8g0h8KEq+CkFOSo7lKxQVCCzm4lPvY6UOdLhACt2UlOOtgk9C+xaez6rWmS0rAJnh0aEL7P7
Lb99uN3tOM1tnc5E9tWlc1TT6Ox/tv2neWiKDa+6etM5DVapTKtS4xSihAoQeGjgW7fVxlJ0tOIb
aptgzha5ICyr4f6ogQraA4A/r94JOx1evETsCbG7RFxppE7HUrSgfQbnVME+UJMxGtm8IAfn4i8y
wHa3LcF+5c2f+C8p7Q5i0MQBjU9C+AnZMIZHNp+Ylv/9KhqHNEomjGZUQ7lEl5G1Ho+ddvPDJmTB
SEkYdlXrERKBVP9C1TMQAdHKShn/J62jQpPRU62ojn9A/cWUf/+boxvuPrY2WBS4zNHbt2IEEffk
Vi0WQMxKSbER2g4He6J/FAHvQZn0crTF1maY45Z50M4rXe/DVxlIwqpifchUFeY3M3HAxDTgKBYG
EDkYgNkia2AOQRKAVTKVTSeAHluq3QBkxt1Csgq9KD4I7pZoJ9qIopYYbB/s1OPQvy6yV9GDaA4k
dBJFbJU0hfWPiZUpoFbbMu3PV7Vs7Gc9yMO4+/aQk3mtMCeVOUqa4GrmN4FYhGBnznRTjFFYjdKf
a9qYHkjN7ag+hTztLukB0PFeY20sjDrGqEbfGyOptBfchk2gwgkPXDmcWoW87M2pQ0Mgnd5S06ZA
6Doqtu30P4ZgGqjmolk9im3PATd1wEqK5UGJGy62JSoGrsR/XbpFc+LpNmNYijwVhaiyy19tKvOc
ljgR2hb1JEpUUL9bnnvG0joSOFlLOENYfF3Ll90HkqhRENau4LCpxQtJtxpVvAhr7JMYLe0slbux
1q6qfPC3LJsVdGF1BTA0rShigMdtTRs055/63TVKuP8yRZwEavZHTqOj79t2U1sveWi/hcBnNWj0
rAGZ4K8CSIZ9xXvMAbKxAJ5aKjPw6IQPEgIcXSCAdbSvH/LD7OQ5J3glRY80BWj55TJpaqYfykQN
7ePAEkWCPlCsFWVuhAC6dUhoQnkfFVikYMQXobTlwgYeMv29n7c18tLA9vO61wYB331gv/1+Hy2Y
hjROwbgB28GXqCEaXtERoAE2XeqtXhy1Ro5FdjduwxAJzyUoeRwAvMGoUizmiiiaj6nFmJ4cgWf7
n0jhu0E1aC38plJ2r3Xxl7FgS8SXrfCqf+DacuPaiC/5MLUI00ofAlhckvJD793RVyqpRRQnh6Wi
MmkCBQgBI+rhCiysoZ1SPTKzhEojBEim54CezWD8LNC4oFKsTkid3qsbOSq5VGBYQZbnAD8G9Otu
Fldm6I1zkgvtM7gq8st6YlDeTUlhH+41sCzo8YeLO8AGsbGZXQVCg/8AqRvFEk6Erek7bsclg3AL
97lmwQKNGdhjM7y0vATA3WXYXyLY9t7gTaOLeeo0iNd05fRH6sS3JRwb21MHYUMJuBMGij3HArWQ
fzh3nte+tBSb36gTZ/cAdOiyJKl4Gnba5kx+QBv2ovDV+jHR3u89+NLFZySFzw5zz5QpRr+9/gdD
dSu8X5Ab/eVKlpwK9LO65a82cq+HVDdmcK5NyjyWzl2agMgQk7iAtzFkR3Z8LvqlQX8GtEICa27V
2jYo8lUaFZcPUbCOfrT6Vq8jC7nXgx3eq8EH36dYG3JQYu/KOZTzeMdqgHuMzKc6mdES6z5JZQIs
ghe4aj+9DXcilURNhEwSfmG4LZbhVfCLUqg9TOCpc2O97l+IlaPiRbs9Dl/GhzZ7x2i8mZz63XlI
t1i6hy0FosATagNGx1qjDTxILux3OmlnpcJ1p/EN/ch+ts6WiAucmmr9XaAoDhNzhzkIcRMAJ6Kj
BPzDMH+pI6djoJm4cQp07EZUISR3X+TAmkdDg/Xp5rY3QZCBd/2SCA1gHtbBijqG4XVhjsoLnUWh
/YHrxErnqUKa+q9TSL6/Zaaot/1Wvunh7lo/MpPqKXNxOSLfnFRDg/Sit/K8b7F0S0kmXp8oaTy0
i0EtZbHSD4CLgI1w1v2/q4yPLPrGO9KHlxDjLwPm6CU2g0ThbN05X1ML1qicQVkec6jgpwqODZrR
545w6P/OxoUsxgSv8wlupZ23QZYo/1J9qU9DBrIqo1J4xStAdNP/pCn2CbcCOo63ctIe+ZDg9teX
NhWn+Ibg5nA2EGW8vY8KUwO1E72lBa4yNIM0BrbvsFW44OJMNDm8VSIESeU22UE5+LeYXZNRoGae
o9mAGr/xMk+CVB+pBuN9xUPrLGFtsGItS0o6bP1+JRq0W9QQbBaISw9zD4ZIHaNaV66mgubfGprE
WcbBZwCPXTs2leExKhoLyIWUW0nsDjsMu7j+Wy0pOwZuPWdaTpMP9bRDR8z1v4kG6e8fsuewv1py
M/YOXoEKtPKZXJDZJL0K86WRkwkMtE/1dOLQYCZRpEG3uHYC9kmzRWN+k9BLd6CUcawDm3U+Xa41
u5/m+ZrylOauZDCmi8ggRF7yXeUDJwORKW42apW+5uw2KjNImP2Kz+8TUFuLZuJN7zCzj+MgsyZ7
oPci3etToqAZO4qe5AwITBZe/yjlkt4ASDh5y+fKyuQETSOeKPp1F6dSlArGaWvWEFW5tKZs3aLq
lB3Cvm+cE/weEv9ypnBUFiWuliw8ZqzMPyKg+3+YQSY2JSdvbB7rI0jz9xD+B0sUOkDWtx0UEWPd
hniNYgX72T0JsZPgEFDEKoGmnyflBTsstrTM8fTofwlFG9DtzXEew8bl4M33LgndYe19kPt7mRM8
BbGYpf3EnXFqO5HWmvA/2uc3irECYvrUW+ipWQMqebVeOz6+0H9p25VaC8WHJiDUENOEo5QwsXm5
j/pZKfjjp0frnDp9ECmn3YE46qYVhlQY09HqfwRa+t6jo8qDadXmNlI8IqfkVzdOBXXrmY5H/BWe
HSlpu9ueRc6ssYskHlYD9L2ePdvl7xktIWsSZUW49wMpYO1yitAv1coE72CksB+R1dWUbT2lB7PR
60b8ijsMYo5TbWYrm4/7ayyCdEuZ3/ftQEvlMMQFaQTgq/gLVjpbKkmo8QLLaYjHRYBWVJsNYYfa
+C7EwFvoWydYkUPjjeGmdOx+2Kgs68OjdftQY0I+CGovabkvoY345OWoNWBswwiWEGsZgsFYgITD
nHA76npBgZSVMSU5ov2OSQ7kAFHko+MLH/srtPD9PzT39M00kkwaaUF6XiI+EmyTkzdK4yDSWlUM
FyxHKbsSiPPX7FjYt4UQSLXSwMaI7AYec80LMXLK7R+5m5zWl5vTh6I4Cyg5SqJjgZnL1FhfLfO5
s+7zqNOs3ohVEqh4FF0MyL5NbiewoRZlBjICL6KP7Admk3kVcDBMLwHF972W3DfyfmxzhsidfrDx
dIip8jqo5VFUBh8TPqeSbWxw8knftMXNS3ho16++171NaSyCatxPTxNBaXHUxz3WtGkx0fr9MyfD
BbDQtgsE9D8vi6UJu/dsRjanQyLLRB8XdPo+JrI6AAR5DTNzt/Usi2ArWJ20y9nkQq3hvWGNnDkd
EMfx/IZsKssx14+S7+Amq0wEzb2b7vCZ/7mx/Rs4M13qsaMlRm8ks+yLv4RH+9oMQjIdOxiWOU5n
XyIzyjtPbjnUPeSYPs79VyXaxxN8CPSfgQwMA62NcMmk0VxpLNuhMIZvPJb0p+O7bBLjcHnUurcD
C/11VTQw1aViOEVF1YVMoCIloKeMa7adZThxN/Sijl3XWuzO4ksbSivL8bIJ2d/cGbsCsA8Ry7zY
qktrqtKIuhPUSC1q9DaN+FXZ8N2QtShSOmc193ivZ33kxSp0q73ganYi3+cCPXfbqvJZkxA9hGD9
LIXAaZl+GHh3Ud//co+5khoG/JyrCiHtelmDfW6iP04Xjoc48u/tXAKgjwsAUuKzzJZE4l3vx+Mk
8zVyJPaDYnUxt3TK3PNvyecRj9ROAw5z26qtWE/JuRf5cwW8oSKo+tx8yFtDhSMpikczYhD4yPt9
Q/roHoKLciB91eoCP+fFzS2NJ8TSLRqwe3CAYGCC8EKvNrgfXjpPEps/O5u6pDIlxLL1qDQ9RtKA
+3ONbxVyfxnTclWmAAUJV5QGPdL6G+c6JXY6A3hy6FOvx7zQddidtikbUNHJjbHYZnh9Bp079TVi
FeN9XFWWjD47yxGH8sfNhLpYDNkZVGZi/v0b2u7MfGeRb8nZ4y3DrvghKSeL+0PPi0YgHBDSkTnz
J8o2F1+7u6eYmY48xEO/qpJculC5pUOGh8SeHD69N4CcoV0ZJ2r2QajYKMwPtDcIlASFSWgOXDWv
I6avYQ2f1zwiCCIWiQyIAot1I8Kwe9xj8aq1JYbXvfk1+JqRQ3osF0vuEwgToFVjGO+hXqnYdu+J
JjwxeOYfgEYsDjLunPOahahU8qbj7c3qAwJhc+0nC7TsYUVp65ch1GJ4SyPkfz59DKxUhZS1bJx+
zTZ3nhHiUM7yGTkJazaldakR88NgC4sJHPN1NW8aMcnSPmfbTy5qDbzzRTnx/3GkgYHBTR9ISVd+
vXrxHAV8lScQDySIVGOd0hkkxQ/tDBPn3eIfvGY9iN4O37VdTHyIgxghuGevWxPAl5iyqdaVfvUa
bjobEK18xdUt4uLWYR2yG0QgebAY+L21gQ36Y7kJzQdk08sWCOFfY9beMsq7comWQntcZA3rNMCG
jSrjIA0CM9mURI/zlv9Y8rwe+GmFZ6vY2Oq4brPicXpDvtHaLCxF/U+5nuZz+xE2oBPcmnTxr3FN
KhobjO81DMJ8XkU5oJna9qjYLNqXCe0uvqzFbYYUlMPr/3SDDHsOzd7vUzGRv70h/MCPTgh9Kcnk
xUTaxtae0LpyR018BiJraQOV7lSBgKQbAePaIO/jbQyxn5j1+QT46OqS8iXU5yMxL9jo25DykbAk
ab1x9KcTK/dwQ4SfrxFTUiUELJyYg8PEyu32doyjA4o4Q54yMeTYYZnwNPY9vwDc/FbwZjeESwMF
M6QAsi4vy6awoGpEnnXqMqzM5YEABC8FzFBLAx+fd316GmDaEkUpCcE+/kfzugVNOp4bcWbox25N
2Kq1rwfqnJJFKgduewkUqxi1m9yXzMC70FulR7XI29NwTuFC07OaubY+3GOAjafFFof89n5DcBQX
4cNgGNDD8rgHPi7yTIH70+3aJ4IA9m7GGzAFfr+QTTOw8Iw6pwIdDgsO5T1IKPA6IDgivQ1Qfhs8
h4RWLG5uYjsbjQgbExQ3XIz7B8a5xsg6McelRMY+F6BzLWMfQlrJqiGyXzD4BVVHCT9kudC7VQ+4
0QlVp/7CkRCubJqcEHKaUW1C8/sN5gQqzfke1N+3CETB4C5PP8e0dGU9gMFx1pMJJ+XJzfex0mNw
ucsA92tVr2tCSLPCcJvbV8FbqUVErAuw/nwSk1/qUIpsJhiZXo7NpGgUsfxiKHRHLOW6UkYevU5G
yZasU4lNWsJCitldL4zRyZi0YlIRC8ULCuiddKQveeI/zodCQe/cPKGAwBSabEDp64pDSB27367J
HMk6GuTQQCCbuuFVL+LR+sTtysf39hgxafrnOQvynNKaElVV12YnSk94958Wh0agpw2dptX0ItPx
tQ7AOxixydgpL0hXQhgpwh8d75DQoPJkxhT9tdMimvKHpX4jFG4VIdpQ7H1lA/bkR7bVUImdVAfs
Wimdyrj7AhNgVadWGoNs3JLWo/MICHmgh+ZFgbCTQGWUuuFnBupDUTzq80UqpmsvOr7rpqoDiCq9
Muhh4NaxmtaAjoG0bvVAiCwOZHnVgciUrgODG8ASvvzvQlMAQKtc3FcPdG0mUkPvwgjAeqeJ5Ber
R1/ycjA9LWWPpTgP7Sea99/7vmdy54tMWuXk1DiT0Ubt19VEyfSHIAJTVuidooht8q+dmRYDwa6+
74URvCQZfmLGrLkVCIoQWDBD+tjY70ACWgIV2ryjw5PYKTErbAkLY9aS0EIPWGxPxZ+dy/BMVvGN
e1SoSQqNF9RZ4fYifmh6sXPQLPacpEAjuLbKRNjtY8kTpV6CQmwlkIZBi9YoI2wehFi7GHlRxOmN
IpsPykCY99XRQ7FTHInHzlOFuzYjbyz7ICjlkIHF7IFMvhwFn/IQallLiXRb9EyD39IzipYEraei
ftM5f6C7NQ5yzcxPJJdbzKVObe+pzk4AZnN8jJu889CR8+ZPsiPWfr4zfHymvyijrcKVddzSNE7l
ZquycbKRzztsb94KBCAKZNfbpBQtrKAKSn62A3fsYFIxV5yYFsQl/FlZz1Zg/QT5B4dCU3qk60K6
5yug8mblqrVY+T3QSHKtLUQ7FjAIVLmm00tEm3FMFW6XVJ++5q5KynaZ6pqOBykJEwQgyoZDXF7Q
R7zlw+ZHTM4RzLdfARSLH6uvmD3VEy8TV+K9dn3p0yWgRASB3mW96EbpSJXA5+ltuSVcdklhRODK
oWnpJUrtalA6qRBOOqZ4RTPvL3A/biZgBfEIH4ZAe4dxMPsfFuE1gJqib4NJ158NAAFnTTtw83AB
OiubhfIaSeYa3fj2P7wXnWwSxRAgsa/sG7zm6aBRhL3KQSbMfBak3qvJHljdes7xT54nYJxKnhfR
bU/Nc5tHr0S+xPUatMNGX5euBvNUSQQRndCyCAhZUkAHMnrtb0sSfXzveucRxNJVw2PXmqKIShuP
BAbCGZB5TLghRiXeLX+wwk1r8b3Kch3PikE4TAI8SGcGAvljdbwxv5gSuHRHh/2D28vpA3n5G+4g
lPa1RRSMn597DsTKLYiNLuvb21fbpa0ScfmXfmj7TOgtSpsSUcJC/ziIkxDCLMQY7y3sBH5Dptdd
VOJysW/8f0oepkTmYjen48Wdo52KeAd2T0qUP4wpEnZjjZ50j1hMLv7oo9GUTHmtQM/vl/xRxrpo
gLbwEpnnvgjeYrkLcf7p59j3tBUSMK892Zdl7LUvbHbnttEOoBaF9odUP+ZTeUyLF+hl9hvI8XyD
Zlc47+GTA4B6JpeHIgetNTvGf+z0dMliYrBhvvRInCYqUblan2job8bQrZHb60pCqWKL6vhllaXN
Igt4dLIzUKXfRf1hv3pZLQHkXALH4V0jVNCothixzLio1eUGP1JW70AOqC4i2BOO7/N2BjQgjcQm
TFp77169V/lH2UmxLLXHWERzD7kz8tsFHZ611to+PtdXT29hNdKbIuG36B6hAEsOzstSMBoeklwq
HmDIVGmJmADyCcUnJCu6UNNe5GqtnlTMAexdMiPPtgeuVhSioZ0waPBhZUveNBByh5nyH4MimKb7
xwTnjYP/k5WxY5cLAYV22/yik39JgmaGkzxNggPYzSMg6dF0AB1+zYcJIfBRSJfsneEhbY8L6QDa
IytHptTV8C5P6Y6WOGwRiSIb4uI5FSReCmIH0Kot+9bEswR0q1vlyHFii5jPwrxkWUVC7FMX/BuQ
I6fLzxs4cL0keSqA73ekIscCe//87T5zTgZzciXAa+Avy7HwHudJfB/U7VgG5aWTaQ0dWhPBjlrR
Zq9gTQUJUeqwwCYZ6jh9f4W8wK1pvoxUjBfrz8p09LTVEN4W0RyjYoKGiQNuLFUpMX/0jiGl/MOJ
9ttZ5pJOBoS3IGHY3pgQmJXBIQneNT1lvJntYb4OwK8erlc8TX2QHGTlQlERNBpbqYeo9ZyMDhfH
pPzKpUYsTGsKujDSBuWOB8SaLK+3CjNoDNU6Be9qpgA99qdXnuDNEHpaCmK1cAvSWaGYrR7hFILZ
s2i7ILawMQ0oajjXKsvlH21YbXpvV0rQweoh8cq0RQOM2eMfUkIjIyX0g/VQq12FBivp4kXTevOL
UdZEuEHznABRbFXHo1ZgbInkWn/wn0Q4kMEGAIwWYiJp/cL1sciWZ2ZX9mrD+gZgcCMm+bfMdIaT
2Yzc3L+u3LONNw9H3+6d2i2bCdrLnipPT4MQ78lUUgSlzTTxQt1Zea7WKHBtcnzLqxEygBc/k8Uc
CxmLBrJlB58+p4iyhftJ42bXYGp/rmcUYbg3flhWkdPjLASlpAdbtmxjbVGjIMuJhHWzRAB3g+Z8
IT7uZZyQ4KJeuYdXgUZhqZbjYCMnZJasP24gFh8lzyOWIOk1L1RPHiW/sH9BrsmoNAKGHmggRL2o
nOfyINLus+4fY7MlRp/umBl2nqd/2wg+rVnOZ0I1ve++D8UkowFx8rgEtUpOMIxEhNRT+eLMMKEH
kl4JK9JUPgK/LHWYYLRgbxNq1J+RVdhFHJ1jF1zRrxLWp9MiZdIJRK2d5ArUxQxgE+REgPy8ZuT3
9GBH5Bvv7lG5dui0vpYh8X21Ps3h26Pxj5vRFILSU3A2XG4vA+x85x3SbvBGokoaJv6k4M4vborB
b/5fvlH0eSYM58wLjvY2ERdAm1Y5p6Js/BhF5j0leJpUKYEiyACxJeBSBpe0Du+M0TTWuznGyHOc
Fj8vIzAqZ3hFHSNT8rZX4B5BQ1E145nVNgEu8lyPJq7r021A2Rn9UHpFr7j4nFHFmSH6UGcZwVMZ
HYKhrAQIIAjl3FT+/TEfxizFHg9VWC4Q/ZyfSbOn/dvH2LSj2hfFkuXdMahHaiM5AG4Jxm5LO5bz
12I3lfxRERFmQ26bbJ57hVg7PPA3aOJcBGtOeBszsMSYDpRnF01/WqMrDtisr93SNJcEfTKc7Xmw
jbMjjyPCzTuRRdQRZ0+BVY8wIFI6NdtxbvvE1Ca8QFfG25LdnP+B5X4L+8VNSgyvXMF7VLlHSM6F
6Ap4pvC2XlasZThOq2S7YAEA4mNyd2clx5aqnO7ocWbGDSeO9sE9kzIKpf+gTldJ/4ELILIGuzNc
5MR1WIBZAg+6FJqbjQ6x2PaJb2/SmRS/w+KQ1Mq/p3aZnOihs3XM554/xv6p62JHkZJP4dQ/29Yv
JoyVyNr3ulACYzv4N4yjwWzbk09iCK40TSFXC+uWf2Qto+hiAdIQjJuF3Z2+a8W+ZxhCdaG3JcLC
WGdElCKZhA1zShaQTbrg8l+DYgCRNnyJhcSaYpIMMGuh8RCNEBSR7NQvxddWUNL/kmtd48L9vBFd
aJoxVidtUOKgMnjeRTnoAip+X1kwH4jcCX+T0f0s9zzd8y9i+xxOpFZTMdndwUNxEwHIsihJhD8k
uKlhfK3U88vJd5An4++KknxsqQUOFwPpDS7E8wA9+EUyfRD+ikUpdQQYsZyNc5QTxAOiJSzTaJIW
o4Ez0Dr+0GM/Layd8/aGNtz5CwoWdp/Pgp90GbjZgqHecEW6WGOiU04sf/RuNXioepUp3qbIqwZ1
3L+X5MkdlX5JdFyMjdkKeQFUykXKkf3+UQ1pkdgJK3Q7TYxT0uIddXgT7mQBQPJY7l4CFmqNQpKN
SsZaWXggPr+Ht3e1R3AlGEc+bbjkp8WrjEgGOdMLB/efGKp70XUkGWc21JiBpM/IGlnMM1s2e0oU
a9gY2na1tey6W5ehvCUTCs9d2ISjHHmCQfJqxlzASQqFcaEYPLHCEsQk74n2Wc8trH7Mn+i7SQaT
atbLNcR7upBfOaY4x0R07iZpwxG4fzRVVCjgzmRbB6cZXoHc5wKfO7QnRArx9BnJxcwE+VD7BOpt
uSr5WJnHyDvWdch1BqrgRlOFnD0MQoJa8Xy2Mw1ioAPKEbMPBNp2zQ3poYSHhMUBX3frIGb4l0Bf
s0diP2Omw4LyamYv81KU+kTWCSVUQIlYUKR3k1yMuBIEL1/SbGd4qDuYUn3JFy9TxZoXXkRH3buW
WfRjQW/0LWD4JC9DWFOi4eZXj1X3H20UheUG/+CkvJDystIjfSX+BhTiAwyVZxMlbaoTyZsF/rCO
IrbvO1Nv5X16d2tqBExdtjo2VYv9/Up4vHtcSfC2hQ2wk49WSdtpRLTc8DicG0vqWnt5LUHvJ+Z9
Xnzpqpr+PyV7sR/kEft7d9Wz4gGSkK7QUjdqzfshq8PrtRl+V4+B6aKMlk1Qg8wVquyvmAlXLhR6
UIs15miyznBMkRuwkPMKKN8sIaVgvbxQhAkfAv7TtIW9LPmdLknF9oDgo5rJCXzVYmuJMvl1qIWq
I3dY3KM6zZIrvFLp95h6pYzNEOPQdp7o0GROkJSHeGLNgiuHZwwcVe/qP9iWVsIZwFJfoubQLmAR
p3x5aZ1/WargdjC1B0Rkg+cDR3k2ke2uTHN0IMIF99OIX+3olW30f6kyY++T9g5BQemvF+/7brvl
tbg0iFwxa1RHFVu+a2tW0euCDjwwJvLk9ZhDbVP2EYL3ekHmNWgl1B3L1Eke9J2ZsdIdUL9rhW5e
wiCjmoZdZIptPXqMoIvzRJ1S+puDJWrlulkPGWfiu7sSig2KgeT3BcdFgu4AvjKmnuhRdkkYTPqb
2FrKtoqZxrDVUuVSSjn1pJf+sO+/cvIS9xbGJm7FoGRiK0Eixq3XEe4KaLZpwqD/zXLyIJhhFMXI
7qcDuF1ntiMlpw4KqeksW/FXufrMMwqwFgxFtZYDMZrKufTXa+XNXqMv9mCsOrPIdZRO5aNz8vbO
TAbgEiG/HQoRLcMKupsDsnpZ/cyGO2Cd+nBV5RPZm+bV9tq2H5dHOTgHOB0cHEOQYdFhR+ua5dI2
3I+cu9MhyNFYDrLVk09kdOQ2XqYFuw0BEp1tBklEIgN6obNWODKmEII0/dkUROwHqds9vv/UCOuJ
bqynV3mD5ZEgEB0hsCikNKY7xmYRJ4ULFa+jzHkk/WgCokJ+XRKe2R1uxdC4+icdyUl6i3vTLiIy
H6WvtxbQFXibVWCf8meDpxTqt2AfhIxDCSs9u8Bqkktq5bIOxM20zfLKSFoFu28wdloF9F95NYf8
P8TJTEFchpv1qN1FIYsFYxQQICjNN3k5x+9wXbYTQYDx6xpXvrj2Dr3E36HXDfNzu16WNBh90NSU
akEt3NIgIht4uF29rxv4WWR03Tt2p+moETWyiv/Gk0oPGHT83ThvOHbvA3xwQ9BJHpc5hrjF9gIw
mAwV6euatYy2p2b/lksZFtJ64p9POCz6Tc8LTrE9/QNKol1+qbINlJM+4Irp9oxvr0ru+6+GYxTl
gvd4//bXXNW83e9znmc6RYWRBDL9pOOEP+audX2Ucn23kgcZptRGBeMs6Zc3CZPIQJFoWy3h8ZP4
+MxKsNXbQmbMpKwzHX4aEEUTCE3syjs4fY2gJcX0Xo8aKI8vOnylLntS9KEz6a6e66V51RGKiwV5
lX/niYZWjQQTnoJM+swUqkBLyFaraBMTZOjjM0eZI2qC9/kqZDfFAczIaVM5MrK83/UigaPVV88Z
klytzIR5ZRCvxIuIVXPq/sDORAiwa8aNDIfqGPcTzn4BbgPDzSgPRwWe2AtM7EPTE3xWwNGfAzUY
cA1R5itwdn40PgsEOMDThNG7vX5DW1TZsbpBLy4OzvCIRdTG6f+pU+JVwiKN/lMRRKQo804poHrw
GGowjabg/j+oEoQgdXQC6UDEyxM0yvqeNrf/SMdduacLxLCRVTlvlIUr8/9Abj4I/s3blivpj2zz
rYfgLWbTV8z2kYGrjmDLG8pN9uP82KSC1JCYpbO/BN0WbpsGZ4NVo0Ei+lcnhzxqprpkZPLA6lCs
SygMOAcb5KR6Vf8MKo6asi0yPhkyFrxQS1XvZXLO6ZQYhIlHyH4ufUiXxAsMFQwU0rMUZoCOzSfW
4pawK3/eVZXMhROUInIuSMQN/vZAHw3IHgJ/F8adfj2IDJFeNKz78HVhJagTcMnccnxGa0GBpxol
6is4Oe60ZEqUBQFXLH5PKAIT9prpoY+qgMvZeVUNatj8UD6L+LNbrNU1fyZSF5NugfFAUDfYCRGj
qPXtULTGjtkR43V4tHNOiS4uust5sXRlSLpknMCz+ywZOhyCrgZnn8tgJck02mBnuTgWe4l82uRu
050WVFxALq3EOU6TvOMng4rpKrLoWYYOyx+lWpIxIq2COwdJzu5Svy5zaSRE6PTeaco9fGh2o1Tk
6y7TsJM3gepAmn3Bact3XwaKpefjLyy6O9cx5ceTRgfisLoR2pbtedFmqS+rIJF5kbSE2Aaoe8PQ
p6VA2gP+pUs9ZJGtY6IZE0q92V5XrqKYmkY0PtbseVQfqRaBF0a7F7ekxIjbi8gorEzV98oRMv5D
EezxdkU0Kq56s0YOCeW5y3iFbSC0atOryASVyJmQ08AEardMZhnXYgMHPFRLRv2w3yogBz2DWQDB
LBZ5dPGZeXX96izxCeDwTfw3SzL6mABWA57Q27OiH0hWQdu/IDd8hrRqFCKzleYGoXA59g5XqkQe
aLVIl6r3bbVcIzjuTg1tSHwLzboIV19qbDm2Q0pCk4mEHCawb1Yzkr+Ft/XNa+h1PGioY3QduX3A
2FnJilFt6TzGoMix+Hbu1prQy5OKfXJw6DT9ee5lZEHuvI2EJhDhD0WsTF/Q5GkNUmqoMgpBLiTM
N2+V63N/KN8jAZZL05kF8OPL+1RxPcuD1dugMyrG1B732qdwZBOlVve58JfgnbwboBQY0gT7R0lc
ejQRnw4GTgobgfgUG7KvpMKAEb0FT/kaAp+rvFxH1eBjDV06Z92/fl3rrOtHsmbV/B7RpAU2K+uI
TiB6JXQKYsZMCrEG83a5zxe3UxPxVlMe7e8HfXcqjgGFoP/QR8MrQc3ZJX/X9DC3cyiKbWYayYhL
SkfqC+br2Hu0mrMX2mNKt0ScfCr+Pa2MIocjYwEZc8ZLManAsi6Wedr71dAkYAWAFp5d8UToLNHz
OG7pzYY6Oeavwo97QEXcydKdUHqBj4vrSP7Y/QleGS3qQrC3eHbiSzJ42XLufLbocwc3iSeY0ADH
t4b0GBRvN39CpEC4Ya4KPEQbKrAE5MnyTqdRfTa1SoPz0Pw0H0yAA3iozEWpRBatNpZ5D77GCtM8
Pr5n0hQwk5YbCOevYsP7rfsWGLr4fbbzrx9CxDn975FLYG6pUTBl+Jx5I2pdMfp+oiW2fV0DwYiN
hLAa4WuwymO10T7jTA99Ukg2Mk77Vi6RcH+3owMM5h0m2p1zWSHCKZPMBpwN6uRmOEHLaYecnDEt
nfiGr1SUbZRJg88JeF30wwIFATmHMglL+AwjR3GtAaxl0NC9yuq7H46oxQ2gZbGqZLLZU838SlzV
St7qZW6mIYPN40FQhf8bCfVcb2Sz+rJRWLVEHs/ipv6tYQNNNikjgM+6T440c05Mw7G70ot520LK
e2bUmBYhtrGYDy5yWrVjczSeIFipKnKaa/gATXmcm41f3CQhrydTsrpzJ8b8VDGl8/Z9VvpDaFeX
b7YZSYQlhj+xCVCLz4UiBPJ9QRPRpiDg5CpKCPkn/iSNiM5A5ZjvOBAkMPbKDBGXJPUHyCJ2HipG
m5DnITeO7kLHPnOMJa2x7q5PGseg4QINfc1Ef/CSY7JGWN+qefzFAt8Fhn1eKVevM4W7xWn5zOCZ
ZUtFjq8VpnOmAuNU/wCmjnXcdmQ8JlfWerI2vvlvbU2/gGWWKU2sGPSkmlRRLLfrdOqreoRnOflt
CFWYURM0J2ce0Aop0kgyBUcXINFLs/2v5PTQ1Xhr1VO5VFL0p/CUaXrTiT+jFC3I5E6lBYPgGMHg
02hJemeU1ZjyE1XVkQaz10RJ/cvA7yGwjYDlavtb+PG5bMAtV/CPeatzMAA4ehwl05QBAh5UH1PJ
ygIvVxeb4/r+RDsHbQJpsDLtnAIK60Cy7AsR+wcky0xi6dXyxEIzUVPCjbWyJ0qYUuGFOscNGRWf
wPDmOt54u9F6hB8RUg9oC8l4vYeO/r1kXPIVnDkoBTG9/X+lkRIowGnXkqoPHq4KLADADSz8DTRs
3gQwVTa2avrjT4Ew/sBBtc/Gy8VTf7aUxypbfjsKVXvoOEuZDxI5f01+88X+vyGi9qb88M+1/Cjd
AILP50lGjCORDn3U7RATKsHUEIOqVTtgtPXEqshZee2+Oz+KBUBv5wtqKXI0KfYRr99nvNTTNYhe
pvgC4b1aoJces9YkqUIErfeP6Mhh4GGif/OGpoLfPIzqzfQa4DcfDGg+9u/Ttv+KmgfnXrFiPDuI
J6On5cdUHVBudlM7gBREjh5s6ZKmOge9tMORcF49OcNp5j9AqMn8xmmRnub33Vsje3r+6v7Xh+NL
QSr8o7CLRF8S5gvT4LuWLPfPdnUY3pVEeg5asJj1jeIaGAmMH3B03b/ccQYJlmYb28BVZWkJGaep
hURQJc17uOdfxZhJqz6meD7bQngiZB6xU+bGctGAHa7jVqoTUGZnsNRtGgJZvJLuYFXy7UOHGkPk
EIvzmucBIeB9zkdcz7l/wpykFQyNtuUFrEdy/6962AY8sTfzwdUU32yXkTkifZtGTW0s5DowyWdM
RAA56nJuRCdPEMeu9L8P4cprRumV3ygfrw/ZyHh2P61HP87mehwhnaR5NN6zDgG56LfAPsT9m5Ld
vP9q4lX5sxTmVCKBpNppFsGYt6lIN3iY74sbt0JElxldDbOY+bCpgEiXMVeyfflwOjH2MYM/Yw3N
Md+bRSL5areg0LRIN62tbWootU9xQo8JTVCwh6+Wmuv25r+/feHrlxw/oe2qCq5W0sLlY8adrU7i
CC+9pNV+Jx5iIpQYK76m/kcS0J9wchL/BqBW+yinAKTnqDNGepuKy1MW8oI78RfLMmhvHCUI2PH6
kLu/SERqns3iUShZsGXu1csDWbnLzNE0r8SwVafZKIBSKdq71SVuPbnP8zk8uP37gXn0wQKhL280
sniBW9LHQlKz9JwFdBNwM/5XK1iUZJeRNxfkuGmkhvIHk4sdUvzZsrjmutbyL/rBvFbCb4mOV+k9
MW7Gv7/E7Jbci92x7hSvysF6ISjyJKrHrq5YISJ5afkMIZ/1Xk0vsBZqFtSlBau2hL1V1lgvG203
aNSL0omPnlR+oYw5zmx8Ng/orSzfhk/T9FnlmpZ7ZAcxqfDEJihMNJlZNlUYvK1r7E5d54fiJODA
Q/GDBKHnwJ9We3X5fwNWl8MUjn1ZjKQj8STvXZAQR0hn9vRNlVx6/xAlV5a7wjeyGvevidYHBSXj
3vPoT/LE1p5AGl6kNAzcJnZPKVm9IAXv1e7rGRGCoQ/OhzX0BzxRYZ4wiYMLdQI68d7crmLWZdh8
Q/RIkBYJHWNC7tR1wxd8tRFhAZ8noV2XrSXRyr+SkCZZgQbIDMSww/Cz0Wx2vrCJnn4fOyGIok3u
2mzTf6tTI3SxxeyMRavvhyJn7qeuwQ3JyHT8GTM6WhmLzRXePUscAyrzk2T3X9CtK+eQ0busaKDZ
OdxRJlmY3PIUxjw7CDOT3wrapzyNwwLDEWi1mHm3GtjuVjeuW1f5jfsQWGk3en8M1rv2DgVxhnto
6IlVMLx2bS4E5DYy63m8cczmVfY873+CQqEVBsCUOjX1EphGLOJPg+h9bm2SCEAsnI+/UA4jWkby
oLzxUFEKdpzHFKfj7ujjfLWqN556ltfU00PRaSZ2I3MfjFis8yR4znYzdQWYK0leE4eIU+5bw+0E
4gNbce448vxFCQKsGBaiufs9COYC8ZJXvxIRiCNeqgzNiPV7QIL57JtZFp4GnYgUh1m0L2m7n70D
h4T4NA2M8bsng2OyQUxltYiAdJnCN5AWNs8dnbTrK0qyM+5fdhyz1FYHjqRxrEcvjuTG/h5uo/Qb
X3Fht2Zx/W0PumdTqT8NzUgIkbVmYeD8nGj39tI28tX3wo42DVrXUZwnnuw0BF9ByM5ev/zMj10C
3kwGULZIwb4vWKFJd/Kql7+v98Op1sNSAMZ9jTmbQGrhSDlTWv9xyy1Hfi5G1YctNw4OsH1PsvaW
BD4ppdMfsqzxjTZOjzEwpNrh4+NxeA0ZogxXo1wvxTA/vv4mjviVJFdNt+qHrCQiKxJJ3xsudjlG
xOegJdTILq9UmU2i8KONh721Rji3ZuY1bH0CKj2uAWGVWfXLtEB5184t7QIc2GJvmYhQyHMKYbQL
gxXP0sHeADNwUVQ3Pab0Nlq9DIti3h5Y51E2D8sHkzyJ/nPrA/zehYtaPgfxIUoGXd7/dhxqx8/m
k3BjMAqNx2b5zEeFn2VsXekEBS5AiUG0fBm5Gc61N3pwtIvfrz3pj55wYboCzUi3nRgR4fkGF3pN
vPL6/HTOVFeZpK5lg1je5HkmiIeGG/BnZD4io+8w9Vv5DNCwZ8Mia+tC5q5p9sTZLyoR0TcZtyMx
dIF0r4VEXW1HNQ4v7E0DQOLSBXEGQfk/RQLQqgFJuodSbWzduZjrT4ExYmLXBBe/PT0fRD7fzzsT
uKkYOk8PnIOAbIhayzOHHOrMCZfSI+IlcFNWBXZssSYCFwmk7Ic+s1brPPYh1BXECZwhhG7GdcbH
tYTiAuXBFPp45wk5SWlokr0N/UBiwUP75H65/1PECWmN5XaJWHqOPnudfcv85+nc8asMxdFeQ45V
uPSD9KybCedXrzZLux4oN7fD/3oH1oygcaXAI5mXA4MpUlvPgPP28KMEjPwN96fLfgeuW7fMEg/s
Wb9nyd49s/tbzw4v+pOpSfg3Teh0Bqv9DV4Y5e1+oHR4yfSWYJAcvM9Ao6wpYtSYU8WUMRH2lQQ7
+rhTnIVxY0rzTwQKeUIm35kjuEpM3NLfh6tEGaJH21Nnm5RTu7TXZD0NWjDskVJmvY4ECfw2ViNU
4d5BD3RxpF2Mdq8zHsvcGvmjgiEeTeXNhCrSEPyoOaW3ltdzHA9AeKLgiTJAmGNUyZcJo02VHU5+
BaemVliIdFM5XY9ca8gCXdw9HzpxkZo2rM7D+N6oXwoGQQgPgLf3QAL2KTHYWQvGGee3Hc0heOYk
uD8Njol6frRtARDBO4mzoWSGm3XIxSs5vKW9cXpI7ztsoEwKrBjhDjNRfwhw8Dh81/x5GNkfOb7E
OMqdJhqna7FKEHd/8Cmv1kNUDGvEMBX9tY5483MG+QjY8fiNa1UaiFD2z1yVtip3dfGGzPplwXYA
LIB3vfYHd2oekS2AL4qiN4suKHw6xOcrG5xBQ5u1354cvRlGfeVScWfH01/sUribVtUq02hp5O5E
CTFQ7C/DBadwNaBlToHZdI2ujpOEt7Q87jBbgPnFw3ZAd/YH/7CwV5kvIV9/T08pCN5L/QSTyCdt
K063OGUe0gBRSCyHNafuAPhvAG+m9LVZkR1gipFW+ve119p1V6hlRQzOUos4SpnAisr8DpCgNNq5
5Iac7DRMv0mRXRPg05Ea6bEbg2juaHKcgXOkv4fgrneY4R+kI/XBGCx12VQiJib0ggFMg+26XkeU
Sjg2TTDHCXmZGoC7tIRBUopRGu2dQFr83EMBeLE/89yneuZ8k2w2zeqpdIqr6W6m9RdPn1cJ7p3Y
hwReEFWAUbtTV2TBMr1ppnLX6JpmBhWN1yCTEyo3ZU+v8QKqaM/6V1Sy6xVsxSrUkaklYBypcas7
hWF8rbfg0HUwH/RMJcE6dlBamVWLIqBHcty6Pfb/elKla8f92Zon4QRSRMA5JSoS6j//7Z2yTWCz
lIOMML2VOB1T0ujxhAcev3NhX4OGoBA2riSpfaMfVEBFrA4Om6Bpeo5gi6uOsFKNSBRoo9rY4lPF
MVqDpW3wV8Pte3uLdPttdQxojpsVh9oh9Qo+LPixrP7HqF4vXeb0IYqdym1dH8iPvh8ZSpODOKbI
UngsuMfggfvKoyeuGzMvWNwV082C1szwYl1MFFEDr8eLsv/3+3Cz0Rnn4oYDHKRymL22XDRfdsto
kfFFJRR/qDAY480MIZMSg/aN6ia1Kr+/gF49w+aV7UNzahSdMkCW0KZX83c8PI7WFipyZLJo/u0c
wQiC3mCs0G5w5vagDqaakGGHM9MrJ91ymE4X8GvrVjGiwq9CVPtcAEQXZMV4Zxh4LV/BhJC/6tKE
cfndKWp8BTYeFLSdrfYQNGiov/lWTy3iR58nLqimIz3zv/Nvt4zzOxc13sNAwrinbyO2+95JB5O0
rU7NWZ09B3wee7e09GCsc3h891VI69AcPihCDRJ7VeIAn/RuK168l7Oi5luc30uzXxpjK1T3+7PJ
3KzWZ9xcRNmpZzi79D57AgAkqnuo5YM/WtLVE8SQ+V+odOlnD3llChQ+3WPu4nX+lQtOG5//L3JQ
NilDNAD1RgRJ29cHxKJbzKSe66Cq+4sGQvYBXnHhMFpBhuqkWTY8Z3xwjl/phS7OWrUKpBfFppFO
SEPVS0AcO4d/Zj6njx87lpd1tCPj+9yn0mkZfYg+2QD+F6LV8wm6PjsbFh/Z6JoYSJONUpmSJ7u8
5UDgVJKNXzaN03Pa+lLhFBijoyFT9opzfWThcInulkij17Sj6urEwGJi4oNaG6S5ECxBlXpzKfdR
fq8efjJWdKFInTQDwkTflipFsO0NyhzbhS35QAqpiDcEISb5+Udu5RsyASC4P3nmjl9G1qiuRWV0
w38gji1bsxR+Xsx9uRywGpdAY95tnE02ah2eMwfvC+iEHmBR5Y8/WFmWy3UGfPmaZJfqhcef8kv6
RnG4b8G5Lw/XNhglQsZNroZDYNkTQO3hp66svNZOzEgxTROfrk2B/YXxLikWTAVzoEFKXkry6yme
2uAo8UE/U9FSxGGd2b0L8F1mDYdmqDgJIDXK3LUDQpqguseiIyoqzln7fBbPrdq54vikzKa3cQsM
frm04zZ5RJFjjbByXpRpNYV+y7OpzOwbxaxYBevTBtgGR1TrHNmhluvuM6TXbn1QtaNL+TLMB5dk
08U8KfvQHYQoZHdUaaT3awPW7oVpCKwodci8t1oEtd5qipYjdgU5+R2LEGawIcRxbMGHvpArykr+
zApsTlBCUownH5ZuvQKcLOh/EFbn3Djwa5vJcnF2FID0rBkokQphhERue5ZZx9Cl5WedeCDeAcPC
ckpL2Ot8RxU8RBmARyhQr3e8vMevyYb00YrNQvSvmU6gsa2dDk0iiVlyeOtn25G2a+NrrJcx3mzt
EZ27qju+N1t7buJUERwwAEJe/7P8xRPGHBgNJqdkgN4O8xFMugelqZpqTkGCX0xBcW4+fTxvAzxG
HZyk7kRT7ztcIflHXm/EuuWqYt+3kQq1SFpfk5wb7bd1Fha6X2woGG2dXSAWG5qRzNfev4EBsvB9
bWolGOp5vCSxVysD3VLSuw6L5GLnbsunJVgQVT7ufJ5dDlsAci5XDa0C6QBkJW90y8RSjKdo5fPu
pXlgUlud2U1IEyzdbMwr2jlMCKhhFhFTxS8SyjVJli2Gb+T4ZPkPHy/vYpy7wcm1pbaDgsSkhf8u
wVXVyXqnyNy0nndXtXkElrGeTGT/oLgCPey0yqPj1qwltcaWDMw1cGv+83J3289evu5WtKOanJlb
6kZfy4sNZnMnThjX418+xRqDKJSFr40O8PdOOGKI6m7YQ7oFGmOJJuxKj8FXDcZjyrvaPamIgxdU
I/Regbrg0YmmI9lIJWyOnpmNmkZbtKsBzESfJAzzxBNoKYyl5yd/pDioS3xkQ4ZJe+jVL8NldAet
vzMeIRF97PtG1b38+FAWMe21F76WCX1Jre+WuT/Y5fdoVB3OPJOazJXfH/BwTDlIzRX9HwxWANWr
LJimJNvt2tjT9195myER+g0AuSg90RjaORI1yElNlb3S+lpeFld90skOdOgHRD+7sWFcu17pLJbi
O1ZSV8IB4aASPQ1F5o+Qx4e1Hpz53eTU0wHgH8xV/o0/95HO9ZSAabBZAV51B9CyedtBRP2WJD3P
o5exTkR8PmlLT07YzVxSpFd7NgpIjJzNKR/HuIFVMeTpHY/L47SnQTjVPUvqoUI/eCep38gl8R/6
ESKF5Rn9n0Q7t9KopSopk3vsRY1wzDe098foJNzN1NlTvqAK0OKzgPxNMgyMmcTPnx/EllobWjTT
4TvRsjGiEBPJ58/LsDaT7q9zyo1qeaiIsYMhu3wt4+VDv/tlqzcZMPtZjG9+kfT5vFAAXnjTs0QX
+HRf21ugKwPTXJIVbQy3WVrSaghjLSBNGOawpeBJc7LYbz6109ONzG/LyQ5OlOzcgIc7Ec4gqdGK
cAeqivAPxxHrY1vgFKYBl2NKeXNspnDfvMP3PHFFAQI3B3vR3k3ZfnI/WsBfNH6bwiRHPbK6MNdY
xrHaCtX6Z8sPtMCc9zbwh3RqN1/OWMD1Z3jHxL0OLBguDgrZoQv8bgtROqPWL5wzduvEDqSeS3T+
1/+RQZ7mrlY0+TRNN9cpPPxhZHJFkXZprbUrxF534rpYnvz2NfLE1m7499+58HxNy4c31naWm9p0
HYHipwCfOAoI21VqzeSS/NTQMMe+2n2cj04f74MyIH3NqN0xOBW2RLglUCXJrXCAIEsoD+hOhGGU
SkMNxF1OD1ZbJFWS5e27paI1pFu7dBgEV9ja7kzaWz2fPdP0ml6Y2hS0KMkD5u48ShAxfOKjPZ6/
wC+wjCXjfSVLeiMesW17vb6bCCO+f9aao37CAE39R0rVm/SZ3xzNNfmvJ7ObkTHctKA25xdqyusL
3G3wjyCxJeUpxIIPyq8ZBv/KRSX/oOzERZDoCVUj0RaWR5IwoNaUrVil4iGZh2un3XTqc+Qau5H9
3+Vya+GCGiGov0MMex1alcNOug2RZpLoE2S5JTRyXT6CgyGkDWcaKkcSbOT/F7SlTSayoWwgNj/w
Y7FW/KeS2YDzNjznkZlfcT3yRgnjLvTo2aLrUEfDHJ9eLmBE2ptXw7yraAuyfDpqaQcXuJ5DtJtv
Ky5Oi8CQX6lfdHnrSc5/E5y4LElDlEnWFJT92K/RsdOpSZ7UAJPA4A4IcC5vD85YRjRBdQk/jbwF
TM6pw0qG9ieDh9YkGkVU763w2WCjpL/kbIZl81nyI1hXb48lhm2Os3rmNYR2m1q6leIEUmV1ofZd
or2ZZs9aHhG2Oltb/0owqF3eXYJrKO/41TdkABes6aYgb/5Cb6X9QB+uO55hr3JbgFEb2+nTXfjI
6G2D4+fY4GUzQJWYw8edjyC44LdlKwVnfcmUnJaL4ZmWh/3aAI/kJMv1TkLBqchXikv/FDrMV7gZ
M1DRIiDfKUEIPxxNRKQTheozSmK1F/B8gY3vd0gOqiGqGwrcjkJ5CRT57zJyDEw0fL0aCILayXtx
2B2N/D2CByVAzO7XN4+rl6tkSCJZfldea3tCp/pSONCwIrFjVv7dTBzClhjkwsSZldcScx1nTigc
Me93ndvsPZtN0NRVMv7cUhqW8RefaCn1iZ4iyGKsaFejEdqKPrN2XJ13s7NX98zNTel3F5i8KLGW
DNXVSw9DPlGM0rlj+LVoz0czAvou7zS1osgYD/YSSKvDS45BEhm+PbaNnS+D7tHEA80XRNrNNh2B
nEWu6zH2PWUftxjbTIbEu9EE3lUom867VuRPY8hiurngXU402sAVRhEg4ebrL9NMgznpqb0FoRJ6
+IcvgtZEIU699pjAkfFgm8keoh6HaHztB6Qt6WLW06E/jDYm5J65kPgPU1FjUJAAVwYWFIjhoqAI
tJQja18Q1PzEwnX9q4MhHJDpVTgJiTaEtNWGGw7FZmgl8UC+yJs3fUrKWR4Qy6nDB3nVguGXSPqJ
mJs1B6nhUUg0MVyrRkPkqBUEamFun1UJ7DIHDBJWEpesADhIc4FUdARZfgzkd7G05jfrqR8Uxa7+
ZPQO4JToKTWYnEcXmz23YLx+UcfZ/wYeU+6D5eQ+fXTZ0UjcGGkpLcI+sWM6+OmE+4w0vILEi1TU
TGRxf94YeidmrmXuRIS4AXeB21BF1Cmc5Q502lGQ6BeTE2KBkbiSuRoyi8H5RBe8XoL4mXO/4Cnd
EnpaRfn4pJMeW/cFstR+mboXkZ8tfkQqFRSSV9YSCt56NuEpcUnSuqAWntIexQK2CxLmYjxZTxEq
Et2MO5bE6sGufZcH804yc05lPcmRcpDd1laVWrs6bMsn5u4RSIumS9AAsVykH4j/SneUsqABqlf/
w6EQMXLCs7VT7nqbNVuxLWNCJrBYoJs8AJy2tENz9Qsk8hmUMdmdae4wlhDqoaMkCtMlFhc6zr8Q
+moixR3XqW2FAsOTmjWy1U209TuzJ1e0qXlS9g5nyuuWB/A8HZsFn0unNrrR5RjLX3uTavjCYNqT
Y3Ey1QFVpRV3io0++6lCcplAmE+nmB/4ox4BzYajSiioqmSMkrkq/XaPOzQrfqF0pP5oDlNHvikS
Qk/s0ApWc0BDQ1WijwMO4LVW31ZykmosaeGO+HH6ewj3amXGLOoGsd+WnE/AhUk2a7eUscHxk/Hk
XDspyyR1KZXNkAuVHspIsK9fBPm6cTJCCUTVYvUt0KJJVvv3kW4sYfTU22CPMzm9ispjg6mU2pT7
/nJGlpLzuZ8We4DsoYUJ/Ptj2/bOuGVLDAVFEguO0yhTynIJoVbU+AIX2p5DH7/x5zHJOSKPTT5W
ma4qFy+Ubx6q5qs3wgsMklYqdEyN2JeH52PW/CoezY2wEYk2glsCy4qNnHesaT+g8Rs1j4O29VDe
tXP1i9W91NjJaBwX5N2h970Id5cASEJ6ymK+zTzJ0Jke52dZWGRFz+teo1Lc4/W0iAfvWBUg+KsH
Zo7eZmLHGXhA3NNFCDebGKskUomLBHbO1giETS7dJcOkElSTIC2SmfSHq3fMZr9bP1Ojsp7IznC4
e2SLf/iTDPHLs9nis0vNisXjIsI8zUd3rciDRCmofYYSeMTnh9G/HrzJPXxfQ4KMNbGqtjOuH9LO
iF+5/E2UC+dU532y9WJE0Ojs4PZd3LaymdnRioVdnN6QrYyNct4QQaIxH0OesGU9R6a9GROiyCs6
y796ndEThiFP1iJwDU2rEeb/Y6khv483wZURkdp+5Ecc8IEj5O3FHY5+17xvoGnSLWshsn657Cjb
GEze8gpA5yjxwek4G2PUrAq+01XQNGuW0nODnmeD8qurc/MWHwnyYigNqaRP36B568Ipu8zIB2l4
oBW+tQCOcbzvW4eMwdlbqClr4x+2IaGG5qkx8Z+mSpS4AHFUYkjJt5DH/VReQLDQ+rLiCKUht/cv
h7AbgC4v9CJoReDSkyqJ69S87QS+yKmzxoIvi+O4MNZmwP3yh0KzizLij0Zx3jj5JANAEs/JT28Q
Y6Fko2tsWUPT4KhaD5EFkwb/Y1LxW3KL/0P3/dzxs7N5RIifgErEmnfGPUBnk1Kjv08Xuf9AZxR5
gY/udCR8XxJLw7NhYvK3VYaF35DVyv3c6M6o5wRMxKuVjVjVEXOAcnd6ygbjNBGQteNUSXuwyxJm
714NetAJ6FIP1qv87mtXqRIXVIUJmPUg7U4qV9lsZYrllncZDISoQkH77Y695lY2JON2EZerQ4Ah
8J733nyh5l3RjIn0ky6aiHAK5i5P1kCYCFmcdbiBncPCecf/nG/zqRiIOTRstayNncIgA+CWR3DG
QE3aMYXsyTkuDUfcw2nVG1pJ5B9gbC2PxQ9+xd78E8/GhR46oESdIEIbwxuJupxJlmerW2XTZB4s
qeBp9V6kU/re/tJc+HrPbe44hBYtUwl6SqkOLYQBGd1WP+kxLevi0v6ef62jVW4mh3fZit0lqu7y
xbkiVD4Jg6RCOy3o1RiuuwErZcbN9hQ2MY4ZQEj4y1yxDu/c91Th4UQJYcGx0C4kEiWOB2f81WZS
+zPYMC4PaLS3SpAGgV4CVQISVekSbMDrSq1IlrBRWIUiwUVRDleMWL4Bk5MtUt5upX5WnrhHmk85
TqA/DOJnnEw9aqPwvQ2badduDKOPV/jfZh3ZgcZCqckADATgdAPA4an3eEaTHEbCMmelAqumlwil
a978aF7MCYpbzfR27Pe6DRYwnt2EFxLpXZvRpJYlYE6eYW7JP3V3t0qGcWXg2oV/lTXdy7jBigDC
L6w6gV+kSGyyuAnaXXLqtK1RZfYAsKkLxpD/2VKVGCEN1FQdosAtKfQGa/HK4PllyJlFX9x1uTQ1
8dyGUNRkNLpzZh5VO/hgG86Ct4fCHgiWxvHfo3WMOIy3QnkliHicXsO8l3R+YnY+pNMAURDvB5wJ
c7pbVycY0RPEjvbjs65iD9gX3ug/TO0HzOE0r2GR2y9SRNUdOUkguDcBrw/12ybhzyGXKBUdH+HH
dvHDIIDwu+GFd3hsMqGxXNCpNQqtRgYE8QcZFDe9M+Il1zgrcYW+gRlmDyuhoLlch8y8tIUfyeVR
Fwgd3QBqFqlt0OwzkH56I3XTS3Snpq1zWp4n/qHK8x7BHadC0UGdWDPrO0PIWAtZRhQaKB2MEGLr
/UEHkqmIfFub/NljZurWfI4xTrK2MGGoaEuWoSaDS6G3IOrzDEM4MMYLeuVyL2ircgC4be2es2jm
OLQF6K146TGO5cu3ta4G2x80jLxmmVwzajjWGTPHj5Zth2Kg8l/27pYmdJv8FGHfAWPq5bi4oZKB
y84vEniYqzV/nuC53yDYmFFibmnbwyTSKI4CplxKSjOcXkdQnKqXQVZZa+Nrk4uY9ZO6dJeNOZY8
g542W/qS3QaIOgPUq4aHBzzjjbKZjtmEpmZ25rMdcLmWfjosUdpZvy8gyw/rh6B/KvMkTwSglBS7
a1qSY96tE88LNyRtpRcBCzdPz7V43kPjGjhprrm0TQs3C8Z5Pv+VoAXdAOj0ViwpAIuRPSWdKAEE
+ckD8FxYj7QVyiGaOXez3B32XeHLz7Jd19d5XZzO77hcEVM+eNGQ2BfevF0lMru4nSKtOrivTYcr
cBKypOJtSwMVURvNc8JxICWoBo1zBwkTca0Sza/ynm/IMNfEbd2R9csUyMp0IvsEevxz3SXy6/OW
EZodZ4NOtt5Cg06ndi3BdJcQhWZ33+XyMa8RqxsKNyWibMtTc5GphNRsvbXoYBl759tjvyCA9w6F
N+lFT0zbQNJ8mz2XXfhppHCkw3WicooaCegcg86mQpF2Gyw6dka8qQFjbxN+2YDhXR760SViHbhq
Lx+W1dCT30R2dtSX3MNDjb8T+FPWApNkXNqWs7IsSsMfmRXyChsZmU41lc09DwqKX8KEd70Ee1rD
ZyKX6+QVW6sCrbW8fFd7V/ZbJ22G1rz+GQE9y/h1pfNVNJvTW829CbeSL/KZxsfcp9jtkEpUuCdn
OOv/3ujBGmsh21L9AcCG0TnLfHfKv7fseFxMZp5n+e01nLD+nMlZBkodxbD0R3j/yFHspHQSv/0t
QAhd+EyQHcejM1hcSGSIXcDMBiDW1V4b2VE0E0IZplbB5DV9Gnya66/hudcCH4XNRsWk9PKyrafb
e9HEom8dwVHjoNLkcTAvElraU6++2K/msS3BRj7YjYSqybILXqFg+2dYQBEFQu/7qb2vMczsWi6t
3MZ+Ca9KLTwAtTEjptiNBQ5z6Jo5RaBAOPdPTTq/ajt6oW3cBJo4qY1v2BydanIRiZkJoHol+qzb
haoBKBt5qRUVX3k9DQMfbsNavCrKBQfjwleTfx++TvNkMVjfDkpRx6LUaM/f4/hAhyGpCKrN0eqL
1BVZzb6uCAzRtL8M9aHgdRc6rsB+GpEjO8nyAQjhFC+gmhSrm+vAl+zHDREVGlzTywT9458I3lrO
S7ScjQb8AyuvTjUy/OUeuibOJvq3M1JGT3IDllhIibhZewoOcqo7wA56cUmaLkJtjU9655UVmc4R
sTwL3sG9zMZdehjnVJ6DXDrjfbWvjOLPTjaNKFbWfVx3TEuKhHoKsTJtL4FXCLfxvUAGtakWDbOM
dzemjg9g5/LCuDL55J0GVwgRAA2lcoL1B83t53XP9HbtZ+FQBDV4fAvmXpDrCnVJAztvBrSf5bE4
izjvKUK5w5OrQrwg3wfhBAEUxZZEMZudSIkgsFKt+7h0XPPx5Kv5NBGCpmsFBj/zyMvjX+vbccYd
o79JNc670Wk99FiWiQ1cWT9zU016MnaRIg2BOGpz5wH6Ytuh/+g2m7dht9buBtn0JULQ7EW3ZQ4Z
fmA3MoU9sovQqEZYKjl2BAa3pyT8nShBsDotpnDb4v0HoOF7NH9fq+oavxrcLTjPk8e6YW8tcHka
ujzN9W9/sLD1meIXd/l+8jhmPoWKZ8iiXi84UKcgOxZKyqAxiko1cwrvFRywpMtviCxiMi9QTNJY
QJYPjfLwu4RgKDFXvHDuUxVXn2IC6tCFS2blyq4w3kps94XR+MvWQEfIEQPSZy39XkhMyXrlTwHT
JivnF/eqAkJ4A3UsHgwiqBRqlSKLTGCLAEB1FcIN6/hyIbZ3flXGBgsKq5jfh1Jy0lGnRPsTnkjX
dJiydD7tg5SWV8JmhrglsNNfDE4ws5gsm9q86UnBv1nNRQhFJOdyDbGaOpJVwDr6+1T2DoQaEsIJ
2+Obps3l7zCT8tTqUrtmHVbJCdogJBHW+Hlj83xc1OZweIgtnewcWzg2wTArcS8HAJMm9RbRjC2p
FUeqABX3OWSDCB3lwPpyOr5XwkVacLB2OYG0nAEM8GR8XpPQAh080xcG9O5e57QkKi6CGvfwLSM7
ubOlyWHyKzHXSKbL7/uLHBCu8NRNFq9Vu+Qer9twQ/F2+BHG7QbWSTKQQjEJFpO6GHwK/tawHPZp
V8FiUdPQCox1ZltlGtsz2S+YJllsAkusicnCrjWZt0xCibOcRQQ96GLYx9iR9gF5c/aZ6zGBqsDm
tnk4ogy4HeXRIwG5/7LkOpARtzbNMjX4cwCZKDwJke89JOrQ0wIh1h8+5V0VUc9DQwi8RjT8xrXU
tMsj1aQi5ech7f5T1hdmdaaUX+gw6td3/UJEFsmuDgk4MVBhynHqpWbQ8QUUhPMQ81qAdnqCEV0q
sSb94oXBXnfKu5Gn8qDXDuvbWOFzOpSdZaNyS67cpznPZ5KOPThf+4cNeIlcONf+p1bFhP66IAU1
Rb2Tv/4u/JrFgrqOL1tbSYnbkpu40NmKZ59n4tOPj39g0rheH7CwPUKtaKSvopihRI6O5tYCX4ki
BrXJ8n9mKuNtO0l/N8mSW/pqydFOztVwHJE9V9YJxdA/ftYprJ1qhSGUYhX0NLduPOrsVElgI4Bx
MWgVE8llUucBmddZ9ah4aTqHkZLe26T6sNQ7EBj7OPQ8b9ITxaH0elF1Ne3W/Hj6PYzCVgRPOmUw
npsZIFZC3JZ0n2libtl6QCGujzgX54jAkBEW7XeQmU96mJJl6925VEB0aaR4qf2Ljndh1eDxG8zC
mMZCWANu3Lox0x5NKHpErttMz6rrtinLfF4YrP1gmsUMavsIm1CNbuNCex1N7Jcd2J+UFCkop9oW
bNgNt57JkjJsL+WFfI2mO5tsE+uxkWFR7ybC3CA108Q2RgWe3OGdh561xjHh447pfUu8bpcWO6KW
/X7P+KkANWORrhAnvYTBvjOgyAN/AY2lLiXGOVvHdQPQOgE05sABRIYQX6UJDotHV807aC/GhCgd
v+XmRLUxkUMpuWQR81ZfHz7kRjLSFIXkMFxygrJdKgV8HlOkEsfnWU8GJKrk22n7s17Ne8XRvsqf
jpP7nnUyv3ozAjwVxQz55zvXqTdvBKpgGdx82yqnWnMMuMToT1ooQm2BtsCvFhYtMY14VGPtB+Fr
I9E3Bmo14QZom5LmToMdaM9JVrUtJ7WLxGT9SpE1jnkfMSaRmaP8QNW0iz3Ee5jYT8WLxAhLCBRW
v0RU/Cer7KBg1Huowia4O/349RSXOIB2BRsxQc+wqMfn4EyWvuIzrp2C8Apoirkyjb0CB+r5fSlc
Y6nkd+8cRG0ztjGiCREIOgvecDCPuYIvpBieQFmKs+3T37burb9ik/z1xGWFbxGqZhlSDxlxsA5w
lG4ikM/4lkZVMfzmGinmDcchfeCGUZbueOaX6Fhk4TmJitMyjIeJ9qdItfw/lELwjorVzwyscIKm
GNxORFRaywwn++3prhqJJiF3DQ16OfjlvNSsey86M+JGck2Zm5+rYSIBzewb7Yxt3qD9od8tgH47
F2fLlv2fvatOwFg9ap2nnT4gItcv7cDvRhkBknIs0LX+om3eL/3C6CVUSZdihDK0lGajJxOUYxU7
TQRz2JtOiqs6lSjLTFdF7IL6138ziHCaY4dXx0glhqsxK/+a6S65qOFbh7frCZZe8F1pqbEofK1n
W9F7tWoU9gl2205WV7+vUvm9E8bkwwgzn6ExArx/yaJrmmFzklZeqZLqVBznk3DLIV0RCjumS9oS
Sh/rpWdgQnenbwBPxMtI/Y0OCwTEZW05rIM8oXHQ0ZD2dAMbHbN0zPDsbL+xsz7fOU5AM4/pl7PR
Qk8c/VJ5P97mmyzXKQEOnv7c5GIBx4azSCRsVHn1oadySugmV/1f5KJ4ZDT0ZwvoFomJhcqp9QSI
ww2h0fwT4IJZIqz1sNExGWPYWaqeD5RDPhHGAtbXXunA6E6GVZ+ut6ubt0DmADZIYRkJyAR4MWcN
+kas/ZN0gB12YfssoFfTuFD7xEhlF6QOUlWG65cmCVcm0wYA1jdwmtO6OGn1tylq1ddXXIhYid/i
QHSsVqcpiAGLZ+e0vCGBWQlD6MBpcnluBtrf31801R9PzhZAHRmgwqOnL7s0ksevnQCkNM2Cy00+
tvbjd7o1Hd/W3ybElUQ0z/RamL4dYkPCLRBST4mLJDiQ9xE/QhaiOR/b5+2Ims7ta+1il/UBz8lU
LIRPVxFxWWc+zdKPEXJc6DKoHgm9o0CBDAyDWrnq57G5JlK/T0X84aMA0G1AwGD8frjiBenEln12
xEH1ztigWEqA4/DDrwI2EsX2slMqitAik3CszrWDh+PRmmOSLf2kcPPHONJFDDUvfkF2TrAOQBcb
5KVzJ0WUwjBQiIOYczB9Rj/oicAnLevvQ1pTEEvjO4liKC5CNHF+W2ycuPtxHWtcFZn271NO8UZZ
iSYEWtIHsf6kDzCBzK6Zuk2UJP2Va03j+35EpAF95ALKP0SqW462dvTXcMMzFvSTvmWjltj//W4k
/L8gVOmS9Luf/VQnWKpDvsP7Tn4FlMOMr1+9FVodQBVRsU5nKEzL9n35Ba2Jss4yycBjxaH/aST5
MQWUEgrrVG0JLXFTtHIccDOKDN/kRtn2tUIHqdzR36BmXVwBHb73pv/dlREyQ6440Ts1KYQrmfZv
YMGLLxwm+4sQvTyqgJa99R7dwgYurfaccq+xqs6dUbKw7evF2IRX54JRZ37YACKchSYnxlwbGKKx
g6+krfzyXwX8rv4Hp7o5rCFljk+pBQzfYo7svKKyOj0xF2oCXijL3CJ7xcUvkpXyJXt4q6DwNosZ
poEU9MbfdkYBXLTatZF29OyHGBz6jY/nLr9zNndLXi/50S1XdXlyMxk11l6GB1+F6zs2tnqNLMib
gGnrXbz3Ia5knFkShMNj/k0X5a5MgQpWNwFDNjzklTpcExhb62LJfuJCQNxsFw5Lve1XVUtwFQvT
dVjudZP9qstLXoq2i45Jy0DPSY6zdNqXh745bU6tViUuEFDid4oVX7dpChBheNSeEWOpEV1t4RHK
DJYpcZNTj/IZ3C/azCHf04JvhadRTAuqzV4Njcd5LmjL1ROlBorIZdVFY1lStcAXrwnaDTq7NXZA
MZTV2fXWDAXhHpMVvPf4F+fNRODmpxVHzAPbmT4yPVNyrhjOIUJaQL4Deue0WftL51Gpe1kzR7Ms
I7eNHYfjmioLh+L6GNf8Pmr6gxPHMptwTDtL3swp/XJTIob9U7kiEqa51xg3J2U2GI5IoWNH5NMX
YG+SFNbVeDXm24yLDLQYibGJecmkuzK7LROkdIVfAuLuIe1sddu1KYFQqTHD0trTxJV6f1lJoZKG
t7gQRIrTlMTFOvTSvKqdnJcinR0r11DWITGYzRmJrYF0sGUrMR8pxTfhNddAcbuE4okB63Q1c5M5
Yc10NeJvM6T6HLHEtVXEdCqsVuUuz+hhQ8ygKoc0GJFIautPpuVZDvUT0R8Xy9BnxJ0V24u6rA8v
QbWLIySncGf9yfswPC20A9WdKdyZazAYVm3fLruWHeOTFym2QUac+LycCS+DWeb/6DIf5+IN6xix
jQ3NvnM8BPzGVtALNeN9Pz5IbCxXwUVVkoewPjRuDFCPPr0W9HobjFChz+N0nu2u/H7XcK2/O38/
+RtOkuY/FkRdQBUqXUDIa3OktFmBrStOWoDGZjNkk09fcgeQZkttHbnGjQym6c9RwL1QOOWcghDA
J0B5R0qIKcjz2756wtqieMzeuuw9Q4JX+54VRqlYt/uNZS4Zgw3JWZi6CTc3Pn5QAaYWBRaEO32v
R4lzHxkM2ke1unoSJZxlDIjgXwYjG4JSXSDfHY1DECZfl6o6yFT5N4kwEeLsbJWrIfnQW0LY77Wa
j9nLaVPYBG6n7foTpSuT976JwJBZ1d2wlqP7QTjOO0DWRcqn4fodC31FgntBkpau/qRmX1E9P0nb
oAwZsaF/3Jjb1PEIPLnC6qvKzsJurQEnX1O82nuDOPVSHzI/F+UkLcQVPbGm2FA+4Ec8L3SkSeai
XKA8m7NVKcdnjhX7IWaBpQd4sMMUfd0Ta+qAx2BYBO8EmInGImtFvYoPmqREwgARN55aHuT9Sxpi
5CpQcYQtyIuwCRdC7yf8++cyPYrzRzc3m2J8Xs1ySV9vmuJOtcjhggJEqgz+CqFEu0c/5MmM/cmu
QtP4N3OP8hJfkN8UX2XWYf47j37JQkh8sZPQCazkyuXaiz0YrqZFs54OIzb/qxNp3GDWG3VAprU9
m6gjD0oogpEX30nxA/r3qP3R3yTsOGjjp3V6NhXQyNbnpoPlQjSbbTfbni5PcDFDm2LI1pfamG9u
6Cb3L1A18yJDkHHOdvE2ERfcsjj1cSJgg9Mvf5ogkL6+xV5WIWXWBw9lYzGaI7l02oE8UMq/6Bks
Qn88xyaZCbLyfoYkpW2yQgCYRlwzFgpYOffRW0wcBH9HPAk2Hw3JouuWbWUamScD8AXOQpjG9HXX
Skn65XfLwvFAWgnIZDe/TfqNOXg+YD0oKbLAl95qn78dkzlqaO3gBxh1gD8gQIoXfRziSTNgvFfC
gX2/zmZEm1VBtvEaul2vVYtHHD70BUs2wucJVAo5FmmbtxOj6nGpy1QtkVmMfTxZ69J5JZ6mS/er
mmvDpmTCFLr+itMdgHBwShQTo9qQpFH9BRICulbK6omEFvU9vOqk+ZdEH5SN8wRtJr3XyVsRLN06
O7RogMoTgB7tETh852yZJ2TX4Bxcp2Ph+2aGP8NDLQlDCfyF9Dk8Ie0UOFh88OJWXk+/PoTmDp3f
V0NfBUigAQLrZgLKTD6Ov9AIO7qa4ArHfpBYJ07RhsqtXIi0mcRqUkIR4XaWGajK/5jymhFTKR3M
WcVSf6TcNSBNgKIizzeM2UKUZVrDXTMooPExKlUMREoAEObvyLntulEXFGtYU2oVk/LstwbzNv7Z
/WVou6GM/8C7s7xv0m/fOCKCIw9unN++eYtU1zamnm5nrwevDoBC+mzTw2iARIl1zOqZPVXaLqAb
sOBVVjQ/jPy/HHLkq9DVFui3W5/qyuSD5XaoAf1exrHUXUnew0ArVxNpmfUeuLqxuLMzSaQGm0pP
1M12CvrufDUZrDen5jk8m3IXhAQTxjzwK9MLlpZOmFHisMY9twf48uoKU0O+NRqAlYWvx9im5Drr
ie3CY4ERHLjWJZkZA9etvNy9mQT047LAgI8XCVduXGmNxTRbnL+59Dfhomr2LOhOQvDBAYf81/lT
U3SAwzBb/l9aWaUJm2SdFPEYI1vMpzdck4IWqg552gi0YXmAunjjibySh0bmQM2kX/4tJPcaYfnw
1TdidD3HIJ4WEsnC/lyuSPIcTMJ7J7gpTOZRTYlj0K+eGE/JxNewROm68ng6CfwpIWETrPAiZhx0
qz62Zfnn3nTAGDLaZ4iLvMffzEAwWW9jyoiBlJjnPm9LswXRg94nFCIyh1SUe0QXs6zPOTODlqJh
sNQpQYb7sLDmTlGDHb2H2erzsslU/tpDpMX9QdIgz/8rR9tLB7ddhxOAv9rFW8oOQq+JA0b53UXy
+scSR4MT0WtcN4NLA5mrDIf1eVoroyyLnwUuujE5PWo1LXdAVrFisBWuoYJYylgvPzJhYna6WR2H
F4MmFBSedxy6tnqb1C34dfs6hbD/8LeLThkUneyLAdu5PWvQ4VHrPUpVFUZXDm+MbfVYcu5tRyE+
I/5/TWUIkPgM7vnD/zevP7yAZzfDZHDYHweomk2zqXdoAZI8eGsnOIeQ5k0EQqxAM8R3cpTi5DqS
uMusLZiRjBc/YYkpHshUmFPpgKXA5iF7Umih0XIU62xHluwzy8Ezgis/bz7hay2EJ3biZ9OE0FSd
LEkb6Rx7zj0365VxMAc3gM7eHNItFWaZWqKnz30yX1wFpxUIfSxLSAnU3jzsxeOnKiJmQAb8OkKl
MPs5Juo6OQFKnb2ffOaLY44CLYmiUezig6aV1MnmTxPVBm4wCuqTdSmiR+p+4k3FHf84eQM9fc1Y
Mq8Ay7o8LPNdrDg9O/9vZ5CI+bzpNbQMPRrkFkSLYTFUe3R2GC2T1qoF0xa00JwbLT4KD2x73BfD
CvFC+fXagwyIbJ6IOD9QJLUBvhnUohLhNHponLePEu2QEifNzjMEpGSTvJLEG3nyyhmLx98AoqYd
TAOOfZenXio0bhtsoJYG4RfNU6XMFsn9WnTV0xK0ct9mwNNusv8ERp12k86g8eYxLcBxOW6gWyfc
HcSuCaHU9yMb9IeIjXrdGUOB51ICkfyPe1Xx5nJzvbdtuZHngelFvxf13Z0ezS7kgvkP7Lx3hrC5
ASvNeLxrpeeeotm6+x0/IqzVd8PCRQ7CKU5BCwOcb7n9s/sZxtDOUDOUW7hxnFKwmiMsPwUCptyJ
U6YFtRfp+mowGP0KBvftRDXc0zO+ePTsRYKKpcdTeCStH+nPUzGMRr+HFYef9XO0tDb/fui/I7uo
44J8WeNCQacn8M2SBbsMj11HujEErEhM6bXepYfuyaJLCic+qClv8AxnhUThVTHSLn7lXi7Pkapl
TIfaDFY+E1sQVbdWmRe6ZbKUtzoe2wIjdIuiOg1lP5LL/FYSSQ5WrBcLT3ja0/kmmPYHx+S/ppum
RVrBEzi26N0kcRxy1iT8/lp16x38dkXPs1ZmdyAY89x3dV7CKF9ZJPq/yGbVemcMMBlFsZ/SKgdj
rVBpcfvP3i2ZoOJM9vAGJ4mxQOs+6gB9z/TvYPk2uZBoZO7tR4zykKpCEmwC0FhoxHg33CexBLoz
YuuHWm2LDnaans/NfA4SaNpiuAgdwEINhjA7TRanNRxcmsDb47ySH/LSbM8wE0ncBMePzeR7P5ya
Ib29XXqc0HcGxaeBKO4VB0TBnqUCYSlvNJO1BSxqUks+O4yVk53rMbW4c3LtVz64HYQl93bUbQIt
LpQelICtyvf9zpBsEMQ4pRGYYsItvCOQWZBXnyJlwG/9dFs4j474CMa+Ggthpk3rAmaEEmvnXBgi
N7EbClC+wUHRyWNWoJpDdq6PtYlIPjuG9LapHCn2/ZBH5UAaTWvj8k8HIaP1DSkay/qIcJzO5Ljr
Tsu6gIv8Ln0NhITDGcCd/5oB2k1qwNp/Jd7kehdU0JdUPDMma3l3x1HYXRgIXA6GuLNnS+2uNN7p
Rw5wfipQiH21opu77mDkS9GM1GDX+SQJ/bs5g+/SoG8gSpYiph0pfBcR5EQJC1DQ72L07+fRwu++
YEz7BtTiyaEK+nlu3LQ47H7nmFziGuvM3GTgjJSHT9bfOKmR7txQEMdCUPXbBlZ+x+vNVvng7ptu
791cfNXjfj7vUHXZqBHkabNFXLUz1rn2193xEUcLs6p5IygNX8XznvBLq+2c5kyahTXtm2u8R6Hl
qV463LB29WjdogmRRcJc1HGGHddh+k3BcNCC0YVGy1/6zyNJP9cjQoFOE5Sxx9XQqD0xxQCm9Nwi
mWUn8NZC73bIvgoBfCJElmqrQSeJKMCPXPj1Jau3nQwy8LRd9jj7ND9IuGqcK5oUF+3zhhzGCbvL
5t8glRCmNowjYlYdz/E0bCmy4uh9Rwqd8qFPFYzf3zsGwOQbGbLYpJkRvMwvdj9qU1PpO2G3t7DU
pzPShIBwe+0HN2/jh/OYmgp7QB+M8e5GEyLpR17arXQz+83RVnig6gtA6FE4YDROlVQqUeHpodj7
uZOXqFtG784F8k0GzTJSE8U4xmOcKAIh1cnAuGBHpq9VNTENNSzVwl9/WD1MByHektJPTDFvhkYq
4ovPJuT3P3K1QC9PMDetuMw+kfGheTydMsZaDdA47joTXoBbEmM1xl9BOHlZYSGrHmIqUmS8+HCD
oI8rzvWGP6ZIqsICi0G/dZSTiFjr2E1r8Jog/OIvO6xfmT4J4iQOJ5YS3lF4z0mcvr2CUrIimY6H
QcTzCFeXz1VL+EvAknD8hUhL5wwZok8gyzIMpTyxz/Uysj6vKe2YK408iWwlL+KBpeHJ/NJFJR4X
lGasMJO2apQEBLexzh0oPXaEEIeSsoPHHsgUB23BPw74nH20/knIRNnFCh623tnhUXqe8CuSCidz
okHB1dUkXGGiudVfZkFant+LfpNoBxuLbV3owwUAHg7qL65hhEfM3uc/LVxIZZQBKfrBDnyNqgvl
2snCWWYWK6UoA3odlQd/UIH+cxDLJq32Zz2Hf3tWstSnvCeQaIitCueKq7+uHvpIkqiIWpsu3CzZ
o3tecbJzxxmL/5mhug4jDgqLKL/CTMkNpjIpaWd2eVj2+TUrotorsvdK+26a86Dstp+2RcUABUbr
iIqTF/yBc+vGE38i7sGQkEazDQV/XrqqbkapkFunJo2vUoquwu1uz4MzS7A3ZBGnCDuFEdQlqdvo
r84WAI7Nk+gHr+kxk20sLrsvrOuLosj1AKd5Zwr1gtlwMv4HsaXo6k29Is+mActey8EWysfojMl6
VimmhPYf63FItrkza7qBIWLIxS+WCv+4oT63iMytA4g18d9bk6icbBk2ULkozJ2Q73liRpjtbec4
44OEjAwiReD9YZB4JlVgH70jPtz42I0GFhCfATkNbQG5ig9Rha4JBaHbWUxLM2b/mb6wlI1jFsU3
wDEEOAI8Gc/PdBkjvSiI0RE0Ppt40VqI8usZn72priocB+AJ1WzDCobhhqWd0XCJIikt5MkCjtpi
0zz1FbgztxdwL845FMd9HEkLqLu/00qXM6lLBKuFh1bsKoWwFWPd3qwPUZ4pb7+k+xEylOz4gc7H
SwkJ9WrpdBh1+nUOQzlzpgP0BGb2AVTS6mi/WZSwraVPXEJiHtkJLDnt7MyhdM/8Kw4PDJQL/JXq
J4qKK/cDWOIMCaVF7OhvJWoiUbrW50syXIRhBsB6IEcgAP4PuZK4GNJ+XAGlRlXmWdUBs3sz4iel
4rHbS8PjanegP553GrodGmcOWZFE1wMAu2gukimcnPi4pzJW7yWP3rJiVIwMWLH2Z2VBXHC7ZP+5
u65v0GSKFjVsVjVZCFe8ofagsFisKOxHQk80Ss5SBeu3hHPp0EfM6PnHoxgU0oE8WUqY4XOf/4A/
0jzCxqJWPMIivVoycG27o6GL2U4hH9q9Ek2Kt9ptLSC5lPRZ+2hUpJ3yevlzUqMTlyKQ6oXFI4e+
CLufFzIX1Yjc+VcYKb4ho/EdAuM02co7OBkCjmnyF59x9TvLuqkFo7ioStMPczdXFZQ95mB6a5oF
SGj02lTefWoayBeIPn+Xke0iWLwHLIdY4ORS2PyhUOE9q9g8kJ3zAGl4N5/zuppPHYZSPYnpSofK
tI51zPpMcnhJMtdw/AaGGv2eiWnfLh1MYQkd3sWnfvF1kmY6xEB3AH3S4+TyHeOJZFYZem8W27eZ
2Gw38W0+xE+/D2iwyy2RZ6X2nciggirFP4ybXaiBC7dvV4GPt4xS+e9xH0m9F2Niv1Ic4b8zptSk
q+Itl1rmCvV++Ns0DqEe1xkNgFV7fx/SfknzHJ46FL5AG3LlTdNStsRct+CqhEa9WnSsGaDbcVYG
WdNagozfoG4jMBrwYfrF5ZN2nU0U0NpnRTpmL/jCVEeuTJwjUmglhhREVExSwWxgEigoBMFkoc9y
q7sL2it1sSU1vL4oPCvZdvs293Pr2QmvNPbrssUHm24g1ysKRgv7vLtdSM2Vu9cY+ZhwmDYPOEPP
j+ewRGjZZixzihPL9yJcALq30QEskCYXEATC1jhor/h2m+o45pYREemL0GM1bw1o2EfjhXIbpIcA
sf3sF7abAtT9w34P1UOmvvZPzwi+fTKDKmk4kahQ/SuJvqyvsBQJZSNLMu3TUZypDoZsHWfaQQ8P
zNxH4mxcP02j3r171dcyj9DJ5o9c5NSTKIEv7lGGV5OpAPU4q4B6AicWM+FV5DuR8V+R9CNb9Hl5
qMC6zOgtINXEmRk6TJjCR2RaYVgY58U5GXVqtKE3QiA4kvgdcYcQaiIS5qx+vQh4RZ1j8IPpjmlf
Tuh2xuLyERcdmxsQrhDXTr9VTjmONDOnEAEAfwDfDe7AHN39JnuMZSG6qBfMzBeX4KaZ7AsHoVyw
8zH/j1sr2jJdmiEbdMMZxJnD6b3OKB47Cy9m/53hXYFD1+iWvF184zKXza3wyd63BBx1pEb/AWJj
Ky9/+OpeAP/WjYUpeDQjGe4haClDsbZJFa3BfxrxSPgPegcK06yMELS6hQOM2WYETzoJFD9TVHtM
+WpwmpWLTYLGMrfkzRcvfFniDKTRZYg+2p8S5yDuqI4/xu89iSwhw3u1Oe4PKcc/7vWHQESftV9I
tUSH3H1IhxSVzILZvi5JHog+IBKBpEOgCp792HB57nRUe3m9sJmDfNYXCq0IHXYq0u4gA/iUPk8y
ek0RcLCnd/ccuWiCoOu8HKjyjbGpMi7Qf7jZTCpiroeShzOWhMVrbrJ6j8Vb8Kb9IU2w5jVciVD8
M+PazYU88X43W6RKhKcsVyQ2/WkYD4Jk1LEWfOqjgeCPzDEsHtbrx1NgWF49/tbL2SJM7YpKmGiS
F7+K3vHUJ5s8Qchgy/k7iehheHPYa8lzFsdsfEwth1aaqEd4DyUFiNbZJSL66jlhiyO2yTGMPr8i
EAILj2xe19Ttyu4oXaHZrebnhgbkzOesLDLbZj/9e5Qcv4ISxv1Cl5fKBsF7I3W7nmzRCbqj5OBk
o2d3wLypgB2E3MhAYJKeKFMNeoVbgM+WyMBhjMRb/8ufO2ksJSkZsVs7IsGKLkUyfeblqxwcaJpy
jTxLjDTAtEdOvQ9TQ6myefrpx3JQ2joF4BNKAKrcIzVPrJCCWGjAQ7uMPF9TVW23h/ujcnuCkf8J
0wjzS+NJlEGg/FnAnunBOp7JX68rshSiKSBaVViZx525ie2eUPhT0ncTf44s8vZ7W3EpsL6lvahJ
Tfj8cG0bbE1ShV/xphLFG3/q7iBbCw9DOGPNWMaNLm//BUV7HgAL/r0MXNEDwLH7mnuaY+TB4AVM
iHpgBtIW5GFsFS11nXT+vaKJCMFA2NT9eW9mENq14cQqOGOrOqmVxnNsXtAlYps82KZRXS1DMmMN
HySIefjRGrRitT80JlS134ktmc/aAl/gojACJ7dMv5AcfOGAgGdDe5E0tiJyQxUJsTOt4KVFa1+k
Db21UwdQ0BoWnXTOsZtTqaV7/r/ew77cFlyVr/zBo6rbKbHkGcyNGkz6sGDPT97FSXK/oTUkFokx
yMe7BV/g4lzaWP3rqLVG9Sk2O18zw8+K4/wQI+7LR8fzWeKkdNIJJOK6kPDIRNqKgXkuPcgGEfDW
z6TfCu/KmbqvzsDOI5WFA35XuxAL7inzOxc6dNwDlkiQoRtxLC8DVZCbnKh9XPICXRDMhlS6SnL2
OAa0ecMKMUhYpPd94ZJNbnDmBIrwUzIvTcNTa8mGAehbyt/8pmnl7Uwx5gv/qX9JRXzVqD8j6OcB
kbo5U7K/bEFOaHAhPEVO822vVkCCygzkHRADZ4oXVzbb4uV+BEsnwONyrD1tQMWW9epN7KBuE6dF
OkyheXz0IIsDe7bNQb3srifHjBE18TmF9riUZ9wf4Cukq+PePqyOpDOYmJ8Onbhkkpo++HsBINdR
7vOWPJAh3ED0m4J5ZUz6vu4JAJNmFO0NLzM2lP/f6n5Nlz/vAEsCDVOgsup/xcdT7a4N+3Vjo5b0
xFWswEAjUFBcWHeum7KDlXL2pALSl83+glodOT14Kp6syIaCHrdaI4n0O9FU9PhHeOCgYW4zu2lA
9tQja8zV68u0vCbHcnUqB661pL+CuCz1HPWauiGkzxvlc1KTUK802e966Cq++qJUM09f+IB3tGKa
U0hBNVJrPWvdbmu7GzjpvcKt3bwVT/++irxO0yKKUVhU0qN2Q2TmaEfwtF6riCadiEMkfBMQkEMT
tmtODpAytBhyVs1n8PArCP0rwLivOKJ85LiuxEZ4ccFY2rekYtX9o6nrr2HMkUKTycGvbYjVuRtm
Qp5j76JNUf/h/xbxlr+fdUJJQUViy7R6cTbfSgSNH+KqjO1ZmNDCN7yrpTkkN/vnqTXVO4NRJT3Y
WzbmpjdGTukYrVYZuAfV0Ij0slBxA2VrqJ69YmzjVadY0dnR20QznZzj0kvF5e91hB+yed+EwC7P
xnLltIwlaRqNafFIuiX2YQdOLo+yDq6Is8u4kWZMYQXyWKCKRFQ01uCJUXfsFi8z3E8UvVIfbNou
w4ftPUxlk9tOP49OMcGHg+lzhDi+GDHzfF3sHAQ+1b6thpm8upC66mHdnkyZKcpXYcvH0F8Y6lKq
dnqyivz+KxjoMQJLYLaxBh3dfQvzNTYVH2unog22N8+EuYFu1Aq/FfHT3xiuquY/pQeuD2rZJgOQ
AhpkxOs6TVB48PVzRa8/jIc6M5EvkUPgKvzUIEALVtxShVJur95IuL5TY128vWSDmkmlhe58b/Dh
4g2o6RgE/wyA2YaBJvb8QTLbZwlM1/1RfDZo0wH3hiLhcTtN8eZgZiMX3i/rRA5+tOBNxWPMN5Ts
Tr3cBM9j74VwtBtd1zQclf7+SDVdw2jKW3vg+OoNn2uG1RVrj/Q757PzeAhg3myoYYmcMXby8cMK
bvCJ/BflvQ10W2qV3yBp7Sj234R0+3WNN4pNBs84eFe33+4KGeHIQYuCMZzKNbIFx3vPojI5bDeM
7DsqgzI/lSyGTK97xgdD+qARkbSOSpXdtTABaPwXLNQQvfhk7NdCvQSZzWpj14p2T5gzCdtXSL+r
YmhQCVHdfCl2JQ1UInf4pw2t14tHynSWJQdUDIzCNNV7qj6Qw6/vTM2uvMcMD4yl1UdcK8cgfNa9
N0dg7X2Cm9taUbCyyvblT0P2ZrchAM5mNUvlj80ZLvuy7MznOu3vHkhq804w7YkkOXnX5XMib7cU
QCnr4THOYnFNWvhPzzbQxdUqWLD9mS+xCnhwKlLn2YaQchggm/1MdHht3Dyp/dUtqdpqvDgTjeBh
WKg3IIelpufjXbatytbWZ9luWldLAauojc/OOrRqgZcnWVPovguc06nHmn+UAF6T9MrC9xYnrnuC
ZIM2rFbhjm0ahLvvj1Udmgs4zsE1C4uwW3j6XdLRsfNy83zp4okngCOIe5ong9AnAklyTxEbvOj5
PrIFK+cjIpZMw+Zaj7Sr45D7An27qhnzCBbR6MUJHFdgHTr8dNoUo/fS1yXZMHkVutaGxxzmlQX8
qXaRpSq0ZjzXwDHVIg6EFX6dxURJPa7yiDcLPEexbRwIu3QaQiWO1ETwMXExQHmsL5p2kL0TExai
x1YxvUPXJvCoKPaem6SR1hgtPXhJECv5dxh8PCz1XyRKAbKsBCCEm2ovJRdQnCMcFMjqw1ysnPO2
51cg9+MdLXwlxEmF7WKg8Sch16WXB/TJCB1DA9IFMOAPo9N5AKqyzDYjoENZw9JLS+EejCdo1pY9
Wvx8Cj5sLsDGm7IfSkCTgnbiRujlqugDXm8RPNFznzl/wCCQ2h3MwlWCRkxk3GqQWRzrZcWm+OOQ
RFE30IZln9YBkmtAS2kxpKaCcEuL5azrXHzpYz9WNBPNErldIVcUToRKdGdsiuWyai+hwPiadYzd
2IU9NKnmxvvAiOzzONnC0ZlaTMIbubNBDPZ5NitIvlbcYh0W/n7Br3FPl5RybinR7SoqoOV3nEvT
9y1Vv864DDqYnXRtGBRCaXMp1z7NSS3wyeOh6PhzSXmubA9Xj26rSkkllY2nIP3cTCmeAk43sTpS
jTn+R3288S2LngjZv/CXDFK7SYtmeL5zbPyVT0wZxL2WuRyh6U5LcFovMZengG5g/HdXWxu0sfao
Q0PSRdTVzjWjKsBH2kZCPQD/uO5oXNn6uIpP0vIUOpZf29RCPJkEurGI6Gb22X6Gx9aN8PB54s6i
R17fXnkWJWihowwPcH7xpdAL+C4e5foZ3i/hJHmtrKnJ9+xP1gpyUifZatEKv7J0aHv44ZvZSzGK
ZsMkCUtXEl+v6rjWEIbntWpwO1bNIZUqjVst50fjIkSdBzzq1OiqdA1zHjm5QuyDEqlBd5zbY5h4
+908q9IpgRq15dm08trUfdDGXTDgJN8/SOyzQ4blLUOl8qo726pn1Zl6TTwZuOSuhNuAp516xRng
Ex4V0fzp3E0yiIVt1wl+uJEwOkADXwLI82Rxh7C9Nx1J0cEglMnk95am4oGidcc0yjnIj+TeVMmp
YnuqtIiq/iIoQGQP3jEEV7u2mellAvNmIcGsWTqZNl/fANTsK/iLtoHW2G+NVWYs2hYlFVwp8tb2
9e6V9rvbg79YOAELCZURKNzlg103KrQd3TbMh78LUZD3pSj/hZFhLETB8amtOMPORY97YXcCe1wt
cr61xmPm+eHDl16WTqVbxjpWQ2jArnKPBCVTw/ynvL5odrMCz0j3U3XFBoY76IK4YlIHJ6BBcaeC
wc3xJufLwNxg/bH7UZBRdMOSbPa/QXx8yIcAjwugLD/eM8GW6HNdXp9EfKkFjT0tjJ000Vr4re6j
S5e3ZAmy4azx2mtYVZ5nd7f/IPLyxUMYCzwk/nMUjwJhgUx7+cdjmUbK6Tu0vQ3M9Z9ZbZs/9WjG
CCOr7loqYDHue5TDQSENocaQ958vc+WwekXoteqB1yxhlWbv0EoYV/cKevvGKADC/I4z2OM8Lu6w
CqVZz5N7dLCJiMkIuCDyjuhxlOCxCWagmTiF++sYi5kQYOX7lOTiSq5SVwihEBcUwZP+HEraY6X9
oNxp7xRpFN9gBgVMKixJbAum8qf7WvmsFEmb2F9ZDhAtDOacK4Pqe8TXhUvNWAqcXKkL3RAKBtEa
SCkKBz0uLDjOgaQwa8G4Nltbk4xHzwF4w9DK/DojYC6g4eJ3dn1AQd1YZSQPVrYQXlFa3roItEbC
B5I76EWXlf8Ow/dBHpgKLi6Tja0rWEUpKPIG9djf/+ZdbcVP07/5H2CXhky9rs3IyJ0Cw322tpO+
+SIOrC/Fw1Grc6ujcEUQeCo6bhe5rvEw8Vm43A8RLYA87uZYlPquWoO2UjG7T5Aw3xWFZ2xN6EIc
75aNh9u2bPk/qcmq6399/AFIepZ/fbuoKHzmt5DnP0ZYE2uda+swnSn+AvljGNuCmAVMc25jX86G
3nEHOQ0y8P+nYufEvQCRNAl+rdbgGv0GhR1RE6Ki3sErrEyMsnksXCrUCft0Lp6jm8Kc6/gZnUVB
gkhbWitM3PYLujiQpC6jATp9ZIdIwlHqHYYBsr3H4gxGT+/qmJwmArcBIhCtTJiQXpH61LjZLh+T
aMwl3ogE8peWXWpvHUDMtF6PhCgvv0k/QQPeQa+gqUaAk8R6C2e+/6FM7+iK
`protect end_protected
